// ================================================================
// NVDLA Open Source Project
//
// Copyright(c) 2016 - 2017 NVIDIA Corporation. Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with
// this distribution for more information.
// ================================================================
// File Name: NV_NVDLA_SDP_CORE_Y_inp.v
`timescale 10ps/1ps
module SDP_Y_INP_mgc_in_wire_wait_v1 (ld, vd, d, lz, vz, z);
  parameter integer rscid = 1;
  parameter integer width = 8;
  input ld;
  output vd;
  output [width-1:0] d;
  output lz;
  input vz;
  input [width-1:0] z;
  wire vd;
  wire [width-1:0] d;
  wire lz;
  assign d = z;
  assign lz = ld;
  assign vd = vz;
endmodule
//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/SDP_Y_INP_mgc_out_stdreg_wait_v1.v
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
// All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------
module SDP_Y_INP_mgc_out_stdreg_wait_v1 (ld, vd, d, lz, vz, z);
  parameter integer rscid = 1;
  parameter integer width = 8;
  input ld;
  output vd;
  input [width-1:0] d;
  output lz;
  input vz;
  output [width-1:0] z;
  wire vd;
  wire lz;
  wire [width-1:0] z;
  assign z = d;
  assign lz = ld;
  assign vd = vz;
endmodule
//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/SDP_Y_INP_mgc_in_wire_v1.v
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
// All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------
module SDP_Y_INP_mgc_in_wire_v1 (d, z);
  parameter integer rscid = 1;
  parameter integer width = 8;
  output [width-1:0] d;
  input [width-1:0] z;
  wire [width-1:0] d;
  assign d = z;
endmodule
//------> ../td_ccore_solutions/leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_0/rtl.v
// ----------------------------------------------------------------------
// HLS HDL: Verilog Netlister
// HLS Version: 10.0/264918 Production Release
// HLS Date: Mon Aug 8 13:35:54 PDT 2016
//
// Generated by: ezhang@hk-sim-11-221
// Generated date: Wed May 31 23:39:52 2017
// ----------------------------------------------------------------------
//
// ------------------------------------------------------------------
// Design Unit: SDP_Y_INP_leading_sign_35_0
// ------------------------------------------------------------------
module SDP_Y_INP_leading_sign_35_0 (
  mantissa, rtn
);
  input [34:0] mantissa;
  output [5:0] rtn;
// Interconnect Declarations
  wire IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_6_2_sdt_2;
  wire IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_18_3_sdt_3;
  wire IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_26_2_sdt_2;
  wire IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_42_4_sdt_4;
  wire IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_50_2_sdt_2;
  wire IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_62_3_sdt_3;
  wire IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_70_2_sdt_2;
  wire IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_90_5_sdt_5;
  wire IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_6_2_sdt_1;
  wire IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_14_2_sdt_1;
  wire IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_26_2_sdt_1;
  wire IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_34_2_sdt_1;
  wire IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_50_2_sdt_1;
  wire IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_58_2_sdt_1;
  wire IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_70_2_sdt_1;
  wire IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_78_2_sdt_1;
  wire IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_96_2_sdt_1;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_9;
  wire c_h_1_12;
  wire c_h_1_13;
  wire c_h_1_14;
  wire c_h_1_16;
  wire[0:0] IntLeadZero_35U_leading_sign_35_0_rtn_and_133_nl;
  wire[0:0] IntLeadZero_35U_leading_sign_35_0_rtn_and_131_nl;
  wire[0:0] IntLeadZero_35U_leading_sign_35_0_rtn_and_138_nl;
  wire[0:0] IntLeadZero_35U_leading_sign_35_0_rtn_and_139_nl;
  wire[0:0] IntLeadZero_35U_leading_sign_35_0_rtn_IntLeadZero_35U_leading_sign_35_0_rtn_or_1_nl;
// Interconnect Declarations for Component Instantiations
  assign IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_6_2_sdt_2 = ~((mantissa[32:31]!=2'b00));
  assign IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_6_2_sdt_1 = ~((mantissa[34:33]!=2'b00));
  assign IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_14_2_sdt_1 = ~((mantissa[30:29]!=2'b00));
  assign c_h_1_2 = IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_6_2_sdt_1 & IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_6_2_sdt_2;
  assign IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_18_3_sdt_3 = (mantissa[28:27]==2'b00)
      & IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_14_2_sdt_1;
  assign IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_26_2_sdt_2 = ~((mantissa[24:23]!=2'b00));
  assign IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_26_2_sdt_1 = ~((mantissa[26:25]!=2'b00));
  assign IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_34_2_sdt_1 = ~((mantissa[22:21]!=2'b00));
  assign c_h_1_5 = IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_26_2_sdt_1 & IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_18_3_sdt_3;
  assign IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_42_4_sdt_4 = (mantissa[20:19]==2'b00)
      & IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_34_2_sdt_1 & c_h_1_5;
  assign IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_50_2_sdt_2 = ~((mantissa[16:15]!=2'b00));
  assign IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_50_2_sdt_1 = ~((mantissa[18:17]!=2'b00));
  assign IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_58_2_sdt_1 = ~((mantissa[14:13]!=2'b00));
  assign c_h_1_9 = IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_50_2_sdt_1 & IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_50_2_sdt_2;
  assign IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_62_3_sdt_3 = (mantissa[12:11]==2'b00)
      & IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_58_2_sdt_1;
  assign IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_70_2_sdt_2 = ~((mantissa[8:7]!=2'b00));
  assign IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_70_2_sdt_1 = ~((mantissa[10:9]!=2'b00));
  assign IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_78_2_sdt_1 = ~((mantissa[6:5]!=2'b00));
  assign c_h_1_12 = IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_70_2_sdt_1 & IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_70_2_sdt_2;
  assign c_h_1_13 = c_h_1_9 & IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_62_3_sdt_3;
  assign c_h_1_14 = c_h_1_6 & IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_42_4_sdt_4;
  assign IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_90_5_sdt_5 = (mantissa[4:3]==2'b00)
      & IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_78_2_sdt_1 & c_h_1_12 & c_h_1_13;
  assign IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_96_2_sdt_1 = ~((mantissa[2:1]!=2'b00));
  assign c_h_1_16 = c_h_1_14 & IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_90_5_sdt_5;
  assign IntLeadZero_35U_leading_sign_35_0_rtn_and_133_nl = c_h_1_14 & (~ IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_90_5_sdt_5);
  assign IntLeadZero_35U_leading_sign_35_0_rtn_and_131_nl = c_h_1_6 & (c_h_1_13 |
      (~ IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_42_4_sdt_4)) & (~ c_h_1_16);
  assign IntLeadZero_35U_leading_sign_35_0_rtn_and_138_nl = c_h_1_2 & (c_h_1_5 |
      (~ IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_18_3_sdt_3)) & (~((~(c_h_1_9
      & (c_h_1_12 | (~ IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_62_3_sdt_3))))
      & c_h_1_14)) & (~ c_h_1_16);
  assign IntLeadZero_35U_leading_sign_35_0_rtn_and_139_nl = IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_6_2_sdt_1
      & (IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_14_2_sdt_1 | (~ IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_6_2_sdt_2))
      & (~((~(IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_26_2_sdt_1 & (IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_34_2_sdt_1
      | (~ IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_26_2_sdt_2)))) & c_h_1_6))
      & (~((~(IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_50_2_sdt_1 & (IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_58_2_sdt_1
      | (~ IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_50_2_sdt_2)) & (~((~(IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_70_2_sdt_1
      & (IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_78_2_sdt_1 | (~ IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_70_2_sdt_2))))
      & c_h_1_13)))) & c_h_1_14)) & (IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_96_2_sdt_1
      | (~ c_h_1_16));
  assign IntLeadZero_35U_leading_sign_35_0_rtn_IntLeadZero_35U_leading_sign_35_0_rtn_or_1_nl
      = ((~((mantissa[34]) | (~((mantissa[33:32]!=2'b01))))) & (~(((mantissa[30])
      | (~((mantissa[29:28]!=2'b01)))) & c_h_1_2)) & (~((~((~((mantissa[26]) | (~((mantissa[25:24]!=2'b01)))))
      & (~(((mantissa[22]) | (~((mantissa[21:20]!=2'b01)))) & c_h_1_5)))) & c_h_1_6))
      & (~((~((~((mantissa[18]) | (~((mantissa[17:16]!=2'b01))))) & (~(((mantissa[14])
      | (~((mantissa[13:12]!=2'b01)))) & c_h_1_9)) & (~((~((~((mantissa[10]) | (~((mantissa[9:8]!=2'b01)))))
      & (~(((mantissa[6]) | (~((mantissa[5:4]!=2'b01)))) & c_h_1_12)))) & c_h_1_13))))
      & c_h_1_14)) & (~((~((mantissa[2:1]==2'b01))) & c_h_1_16))) | ((~ (mantissa[0]))
      & IntLeadZero_35U_leading_sign_35_0_rtn_wrs_c_96_2_sdt_1 & c_h_1_16);
  assign rtn = {c_h_1_16 , (IntLeadZero_35U_leading_sign_35_0_rtn_and_133_nl) , (IntLeadZero_35U_leading_sign_35_0_rtn_and_131_nl)
      , (IntLeadZero_35U_leading_sign_35_0_rtn_and_138_nl) , (IntLeadZero_35U_leading_sign_35_0_rtn_and_139_nl)
      , (IntLeadZero_35U_leading_sign_35_0_rtn_IntLeadZero_35U_leading_sign_35_0_rtn_or_1_nl)};
endmodule
//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v4.v
module SDP_Y_INP_mgc_shift_l_v4(a,s,z);
   parameter width_a = 4;
   parameter signd_a = 1;
   parameter width_s = 2;
   parameter width_z = 8;
   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;
   generate
   if (signd_a)
   begin: SIGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSIGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate
//Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      int olen = width_z;
      int ilen = width_a+1;
      int len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 = result[olen-1:0];
      end
   endfunction // fshl_u
//Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u
endmodule
//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/mgc_shift_bl_beh_v4.v
module SDP_Y_INP_mgc_shift_bl_v4(a,s,z);
   parameter width_a = 4;
   parameter signd_a = 1;
   parameter width_s = 2;
   parameter width_z = 8;
   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;
   generate if ( signd_a )
   begin: SIGNED
     assign z = fshl_s(a,s,a[width_a-1]);
   end
   else
   begin: UNSIGNED
     assign z = fshl_s(a,s,1'b0);
   end
   endgenerate
//Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      int olen = width_z;
      int ilen = width_a+1;
      int len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 = result[olen-1:0];
      end
   endfunction // fshl_u
//Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u
//Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      int olen = width_z;
      int ilen = signd_a ? width_a : width_a+1;
      int len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u = result[olen-1:0];
      end
   endfunction // fshl_u
//Shift left - signed shift argument
   function [width_z-1:0] fshl_s;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      reg [width_a:0] sbit_arg1;
      begin
// Ignoring the possibility that arg2[width_s-1] could be X
// because of customer complaints regarding X'es in simulation results
        if ( arg2[width_s-1] == 1'b0 )
        begin
          sbit_arg1[width_a:0] = {(width_a+1){1'b0}};
          fshl_s = fshl_u(arg1, arg2, sbit);
        end
        else
        begin
          sbit_arg1[width_a] = sbit;
          sbit_arg1[width_a-1:0] = arg1;
          fshl_s = fshr_u(sbit_arg1[width_a:1], ~arg2, sbit);
        end
      end
   endfunction
endmodule
//------> ../td_ccore_solutions/leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_0/rtl.v
// ----------------------------------------------------------------------
// HLS HDL: Verilog Netlister
// HLS Version: 10.0/264918 Production Release
// HLS Date: Mon Aug 8 13:35:54 PDT 2016
//
// Generated by: ezhang@hk-sim-11-136
// Generated date: Fri Jun 16 21:48:25 2017
// ----------------------------------------------------------------------
//
// ------------------------------------------------------------------
// Design Unit: SDP_Y_INP_leading_sign_49_0
// ------------------------------------------------------------------
module SDP_Y_INP_leading_sign_49_0 (
  mantissa, rtn
);
  input [48:0] mantissa;
  output [5:0] rtn;
// Interconnect Declarations
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_2;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_2;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_2;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_2;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_2;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_2;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1;
  wire IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_9;
  wire c_h_1_12;
  wire c_h_1_13;
  wire c_h_1_14;
  wire c_h_1_17;
  wire c_h_1_20;
  wire c_h_1_21;
  wire c_h_1_22;
  wire c_h_1_23;
  wire[0:0] IntLeadZero_49U_leading_sign_49_0_rtn_and_189_nl;
  wire[0:0] IntLeadZero_49U_leading_sign_49_0_rtn_and_187_nl;
  wire[0:0] IntLeadZero_49U_leading_sign_49_0_rtn_and_194_nl;
  wire[0:0] IntLeadZero_49U_leading_sign_49_0_rtn_and_195_nl;
  wire[0:0] IntLeadZero_49U_leading_sign_49_0_rtn_IntLeadZero_49U_leading_sign_49_0_rtn_or_1_nl;
// Interconnect Declarations for Component Instantiations
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_2 = ~((mantissa[46:45]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1 = ~((mantissa[48:47]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1 = ~((mantissa[44:43]!=2'b00));
  assign c_h_1_2 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_2;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3 = (mantissa[42:41]==2'b00)
      & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_2 = ~((mantissa[38:37]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1 = ~((mantissa[40:39]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1 = ~((mantissa[36:35]!=2'b00));
  assign c_h_1_5 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4 = (mantissa[34:33]==2'b00)
      & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1 & c_h_1_5;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_2 = ~((mantissa[30:29]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1 = ~((mantissa[32:31]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1 = ~((mantissa[28:27]!=2'b00));
  assign c_h_1_9 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_2;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3 = (mantissa[26:25]==2'b00)
      & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_2 = ~((mantissa[22:21]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1 = ~((mantissa[24:23]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1 = ~((mantissa[20:19]!=2'b00));
  assign c_h_1_12 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_2;
  assign c_h_1_13 = c_h_1_9 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3;
  assign c_h_1_14 = c_h_1_6 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5 = (mantissa[18:17]==2'b00)
      & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1 & c_h_1_12 & c_h_1_13;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_2 = ~((mantissa[14:13]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1 = ~((mantissa[16:15]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1 = ~((mantissa[12:11]!=2'b00));
  assign c_h_1_17 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_2;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3 = (mantissa[10:9]==2'b00)
      & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_2 = ~((mantissa[6:5]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1 = ~((mantissa[8:7]!=2'b00));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1 = ~((mantissa[4:3]!=2'b00));
  assign c_h_1_20 = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_2;
  assign c_h_1_21 = c_h_1_17 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4 = (mantissa[2:1]==2'b00)
      & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1 & c_h_1_20;
  assign c_h_1_22 = c_h_1_21 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4;
  assign c_h_1_23 = c_h_1_14 & IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5;
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_189_nl = c_h_1_14 & (c_h_1_22
      | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_90_5_sdt_5));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_187_nl = c_h_1_6 & (c_h_1_13 |
      (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_42_4_sdt_4)) & (~((~(c_h_1_21
      & (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_134_4_sdt_4))) & c_h_1_23));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_194_nl = c_h_1_2 & (c_h_1_5 |
      (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_18_3_sdt_3)) & (~((~(c_h_1_9
      & (c_h_1_12 | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_62_3_sdt_3))))
      & c_h_1_14)) & (~(((~(c_h_1_17 & (c_h_1_20 | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_110_3_sdt_3))))
      | c_h_1_22) & c_h_1_23));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_and_195_nl = IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_1
      & (IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_14_2_sdt_1 | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_6_2_sdt_2))
      & (~((~(IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_1 & (IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_34_2_sdt_1
      | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_26_2_sdt_2)))) & c_h_1_6))
      & (~((~(IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_1 & (IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_58_2_sdt_1
      | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_50_2_sdt_2)) & (~((~(IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_1
      & (IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_78_2_sdt_1 | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_70_2_sdt_2))))
      & c_h_1_13)))) & c_h_1_14)) & (~(((~(IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_1
      & (IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_106_2_sdt_1 | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_98_2_sdt_2))
      & (~((~(IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_1 & (IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_126_2_sdt_1
      | (~ IntLeadZero_49U_leading_sign_49_0_rtn_wrs_c_118_2_sdt_2)))) & c_h_1_21))))
      | c_h_1_22) & c_h_1_23));
  assign IntLeadZero_49U_leading_sign_49_0_rtn_IntLeadZero_49U_leading_sign_49_0_rtn_or_1_nl
      = ((~((mantissa[48]) | (~((mantissa[47:46]!=2'b01))))) & (~(((mantissa[44])
      | (~((mantissa[43:42]!=2'b01)))) & c_h_1_2)) & (~((~((~((mantissa[40]) | (~((mantissa[39:38]!=2'b01)))))
      & (~(((mantissa[36]) | (~((mantissa[35:34]!=2'b01)))) & c_h_1_5)))) & c_h_1_6))
      & (~((~((~((mantissa[32]) | (~((mantissa[31:30]!=2'b01))))) & (~(((mantissa[28])
      | (~((mantissa[27:26]!=2'b01)))) & c_h_1_9)) & (~((~((~((mantissa[24]) | (~((mantissa[23:22]!=2'b01)))))
      & (~(((mantissa[20]) | (~((mantissa[19:18]!=2'b01)))) & c_h_1_12)))) & c_h_1_13))))
      & c_h_1_14)) & (~(((~((~((mantissa[16]) | (~((mantissa[15:14]!=2'b01))))) &
      (~(((mantissa[12]) | (~((mantissa[11:10]!=2'b01)))) & c_h_1_17)) & (~((~((~((mantissa[8])
      | (~((mantissa[7:6]!=2'b01))))) & (~(((mantissa[4]) | (~((mantissa[3:2]!=2'b01))))
      & c_h_1_20)))) & c_h_1_21)))) | c_h_1_22) & c_h_1_23))) | ((~ (mantissa[0]))
      & c_h_1_22 & c_h_1_23);
  assign rtn = {c_h_1_23 , (IntLeadZero_49U_leading_sign_49_0_rtn_and_189_nl) , (IntLeadZero_49U_leading_sign_49_0_rtn_and_187_nl)
      , (IntLeadZero_49U_leading_sign_49_0_rtn_and_194_nl) , (IntLeadZero_49U_leading_sign_49_0_rtn_and_195_nl)
      , (IntLeadZero_49U_leading_sign_49_0_rtn_IntLeadZero_49U_leading_sign_49_0_rtn_or_1_nl)};
endmodule
//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/mgc_shift_r_beh_v4.v
module SDP_Y_INP_mgc_shift_r_v4(a,s,z);
   parameter width_a = 4;
   parameter signd_a = 1;
   parameter width_s = 2;
   parameter width_z = 8;
   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;
   generate
     if (signd_a)
     begin: SIGNED
       assign z = fshr_u(a,s,a[width_a-1]);
     end
     else
     begin: UNSIGNED
       assign z = fshr_u(a,s,1'b0);
     end
   endgenerate
//Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      int olen = width_z;
      int ilen = signd_a ? width_a : width_a+1;
      int len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u = result[olen-1:0];
      end
   endfunction // fshl_u
endmodule
//------> ../td_ccore_solutions/leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_0/rtl.v
// ----------------------------------------------------------------------
// HLS HDL: Verilog Netlister
// HLS Version: 10.0/264918 Production Release
// HLS Date: Mon Aug 8 13:35:54 PDT 2016
//
// Generated by: ezhang@hk-sim-10-192
// Generated date: Thu Dec 8 22:25:07 2016
// ----------------------------------------------------------------------
//
// ------------------------------------------------------------------
// Design Unit: SDP_Y_INP_leading_sign_23_0
// ------------------------------------------------------------------
module SDP_Y_INP_leading_sign_23_0 (
  mantissa, rtn
);
  input [22:0] mantissa;
  output [4:0] rtn;
// Interconnect Declarations
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_2;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_2;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_2;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_9;
  wire c_h_1_10;
  wire[0:0] IntLeadZero_23U_leading_sign_23_0_rtn_and_85_nl;
  wire[0:0] IntLeadZero_23U_leading_sign_23_0_rtn_and_83_nl;
  wire[0:0] IntLeadZero_23U_leading_sign_23_0_rtn_and_90_nl;
  wire[0:0] IntLeadZero_23U_leading_sign_23_0_rtn_IntLeadZero_23U_leading_sign_23_0_rtn_or_2_nl;
// Interconnect Declarations for Component Instantiations
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_2 = ~((mantissa[20:19]!=2'b00));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1 = ~((mantissa[22:21]!=2'b00));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1 = ~((mantissa[18:17]!=2'b00));
  assign c_h_1_2 = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1 & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_2;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3 = (mantissa[16:15]==2'b00)
      & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_2 = ~((mantissa[12:11]!=2'b00));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1 = ~((mantissa[14:13]!=2'b00));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1 = ~((mantissa[10:9]!=2'b00));
  assign c_h_1_5 = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1 & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4 = (mantissa[8:7]==2'b00)
      & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1 & c_h_1_5;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_2 = ~((mantissa[4:3]!=2'b00));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1 = ~((mantissa[6:5]!=2'b00));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1 = ~((mantissa[2:1]!=2'b00));
  assign c_h_1_9 = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1 & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_2;
  assign c_h_1_10 = c_h_1_6 & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_and_85_nl = c_h_1_6 & (~ IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4);
  assign IntLeadZero_23U_leading_sign_23_0_rtn_and_83_nl = c_h_1_2 & (c_h_1_5 | (~
      IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3)) & (c_h_1_9 | (~ c_h_1_10));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_and_90_nl = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1
      & (IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1 | (~ IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_2))
      & (~((~(IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1 & (IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1
      | (~ IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_2)))) & c_h_1_6))
      & (~((~(IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1 & (IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1
      | (~ IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_2)))) & c_h_1_10));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_IntLeadZero_23U_leading_sign_23_0_rtn_or_2_nl
      = ((~((mantissa[22]) | (~((mantissa[21:20]!=2'b01))))) & (~(((mantissa[18])
      | (~((mantissa[17:16]!=2'b01)))) & c_h_1_2)) & (~((~((~((mantissa[14]) | (~((mantissa[13:12]!=2'b01)))))
      & (~(((mantissa[10]) | (~((mantissa[9:8]!=2'b01)))) & c_h_1_5)))) & c_h_1_6))
      & (~((~((~((mantissa[6]) | (~((mantissa[5:4]!=2'b01))))) & (~((~((mantissa[2:1]==2'b01)))
      & c_h_1_9)))) & c_h_1_10))) | ((~ (mantissa[0])) & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1
      & c_h_1_9 & c_h_1_10);
  assign rtn = {c_h_1_10 , (IntLeadZero_23U_leading_sign_23_0_rtn_and_85_nl) , (IntLeadZero_23U_leading_sign_23_0_rtn_and_83_nl)
      , (IntLeadZero_23U_leading_sign_23_0_rtn_and_90_nl) , (IntLeadZero_23U_leading_sign_23_0_rtn_IntLeadZero_23U_leading_sign_23_0_rtn_or_2_nl)};
endmodule
//------> ../td_ccore_solutions/leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_0/rtl.v
// ----------------------------------------------------------------------
// HLS HDL: Verilog Netlister
// HLS Version: 10.0/264918 Production Release
// HLS Date: Mon Aug 8 13:35:54 PDT 2016
//
// Generated by: ezhang@hk-sim-11-123
// Generated date: Thu May 11 16:20:10 2017
// ----------------------------------------------------------------------
//
// ------------------------------------------------------------------
// Design Unit: SDP_Y_INP_leading_sign_10_0
// ------------------------------------------------------------------
module SDP_Y_INP_leading_sign_10_0 (
  mantissa, rtn
);
  input [9:0] mantissa;
  output [3:0] rtn;
// Interconnect Declarations
  wire IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_6_2_sdt_2;
  wire IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_18_3_sdt_3;
  wire IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_6_2_sdt_1;
  wire IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_14_2_sdt_1;
  wire c_h_1_2;
  wire c_h_1_3;
  wire IntLeadZero_10U_leading_sign_10_0_rtn_and_35_ssc;
  wire[0:0] IntLeadZero_10U_leading_sign_10_0_rtn_and_31_nl;
  wire[0:0] IntLeadZero_10U_leading_sign_10_0_rtn_IntLeadZero_10U_leading_sign_10_0_rtn_or_nl;
  wire[0:0] IntLeadZero_10U_leading_sign_10_0_rtn_IntLeadZero_10U_leading_sign_10_0_rtn_nor_6_nl;
// Interconnect Declarations for Component Instantiations
  assign IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_6_2_sdt_2 = ~((mantissa[7:6]!=2'b00));
  assign IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_6_2_sdt_1 = ~((mantissa[9:8]!=2'b00));
  assign IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_14_2_sdt_1 = ~((mantissa[5:4]!=2'b00));
  assign c_h_1_2 = IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_6_2_sdt_1 & IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_6_2_sdt_2;
  assign IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_18_3_sdt_3 = (mantissa[3:2]==2'b00)
      & IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_14_2_sdt_1;
  assign c_h_1_3 = c_h_1_2 & IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_18_3_sdt_3;
  assign IntLeadZero_10U_leading_sign_10_0_rtn_and_35_ssc = (mantissa[1:0]==2'b00)
      & c_h_1_3;
  assign IntLeadZero_10U_leading_sign_10_0_rtn_and_31_nl = c_h_1_2 & (~ IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_18_3_sdt_3);
  assign IntLeadZero_10U_leading_sign_10_0_rtn_IntLeadZero_10U_leading_sign_10_0_rtn_or_nl
      = (IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_6_2_sdt_1 & (IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_14_2_sdt_1
      | (~ IntLeadZero_10U_leading_sign_10_0_rtn_wrs_c_6_2_sdt_2)) & (~ c_h_1_3))
      | IntLeadZero_10U_leading_sign_10_0_rtn_and_35_ssc;
  assign IntLeadZero_10U_leading_sign_10_0_rtn_IntLeadZero_10U_leading_sign_10_0_rtn_nor_6_nl
      = ~((mantissa[9]) | (~((mantissa[8:7]!=2'b01))) | (((mantissa[5]) | (~((mantissa[4:3]!=2'b01))))
      & c_h_1_2) | ((mantissa[1]) & c_h_1_3) | IntLeadZero_10U_leading_sign_10_0_rtn_and_35_ssc);
  assign rtn = {c_h_1_3 , (IntLeadZero_10U_leading_sign_10_0_rtn_and_31_nl) , (IntLeadZero_10U_leading_sign_10_0_rtn_IntLeadZero_10U_leading_sign_10_0_rtn_or_nl)
      , (IntLeadZero_10U_leading_sign_10_0_rtn_IntLeadZero_10U_leading_sign_10_0_rtn_nor_6_nl)};
endmodule
//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/mgc_shift_br_beh_v4.v
module SDP_Y_INP_mgc_shift_br_v4(a,s,z);
   parameter width_a = 4;
   parameter signd_a = 1;
   parameter width_s = 2;
   parameter width_z = 8;
   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;
   generate
     if (signd_a)
     begin: SIGNED
       assign z = fshr_s(a,s,a[width_a-1]);
     end
     else
     begin: UNSIGNED
       assign z = fshr_s(a,s,1'b0);
     end
   endgenerate
//Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      int olen = width_z;
      int ilen = width_a+1;
      int len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 = result[olen-1:0];
      end
   endfunction // fshl_u
//Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      int olen = width_z;
      int ilen = signd_a ? width_a : width_a+1;
      int len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u = result[olen-1:0];
      end
   endfunction // fshr_u
//Shift right - signed shift argument
   function [width_z-1:0] fshr_s;
     input [width_a-1:0] arg1;
     input [width_s-1:0] arg2;
     input sbit;
     begin
       if ( arg2[width_s-1] == 1'b0 )
       begin
         fshr_s = fshr_u(arg1, arg2, sbit);
       end
       else
       begin
         fshr_s = fshl_u_1({arg1, 1'b0},~arg2, sbit);
       end
     end
   endfunction
endmodule
//------> ./rtl.v
// ----------------------------------------------------------------------
// HLS HDL: Verilog Netlister
// HLS Version: 10.0/264918 Production Release
// HLS Date: Mon Aug 8 13:35:54 PDT 2016
//
// Generated by: ezhang@hk-sim-10-159
// Generated date: Mon Jul 3 16:24:03 2017
// ----------------------------------------------------------------------
//
// ------------------------------------------------------------------
// Design Unit: SDP_Y_INP_chn_inp_out_rsci_unreg
// ------------------------------------------------------------------
module SDP_Y_INP_chn_inp_out_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_Y_INP_chn_inp_in_rsci_unreg
// ------------------------------------------------------------------
module SDP_Y_INP_chn_inp_in_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: NV_NVDLA_SDP_CORE_Y_inp_core_core_fsm
// FSM Module
// ------------------------------------------------------------------
module NV_NVDLA_SDP_CORE_Y_inp_core_core_fsm (
  nvdla_core_clk, nvdla_core_rstn, core_wen, fsm_output
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;
// FSM State Type Declaration for NV_NVDLA_SDP_CORE_Y_inp_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;
  reg [0:0] state_var;
  reg [0:0] state_var_NS;
// Interconnect Declarations for Component Instantiations
  always @(*)
  begin : NV_NVDLA_SDP_CORE_Y_inp_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
// core_rlp_C_0
      default : begin
        fsm_output = 2'b1;
        state_var_NS = main_C_0;
      end
    endcase
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: NV_NVDLA_SDP_CORE_Y_inp_core_staller
// ------------------------------------------------------------------
module NV_NVDLA_SDP_CORE_Y_inp_core_staller (
  nvdla_core_clk, nvdla_core_rstn, core_wen, chn_inp_in_rsci_wen_comp, core_wten,
      chn_inp_out_rsci_wen_comp
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output core_wen;
  input chn_inp_in_rsci_wen_comp;
  output core_wten;
  reg core_wten;
  input chn_inp_out_rsci_wen_comp;
// Interconnect Declarations for Component Instantiations
  assign core_wen = chn_inp_in_rsci_wen_comp & chn_inp_out_rsci_wen_comp;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      core_wten <= 1'b0;
    end
    else begin
      core_wten <= ~ core_wen;
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_out_rsci_chn_inp_out_wait_dp
// ------------------------------------------------------------------
module NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_out_rsci_chn_inp_out_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_inp_out_rsci_oswt, chn_inp_out_rsci_bawt,
      chn_inp_out_rsci_wen_comp, chn_inp_out_rsci_biwt, chn_inp_out_rsci_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_inp_out_rsci_oswt;
  output chn_inp_out_rsci_bawt;
  output chn_inp_out_rsci_wen_comp;
  input chn_inp_out_rsci_biwt;
  input chn_inp_out_rsci_bdwt;
// Interconnect Declarations
  reg chn_inp_out_rsci_bcwt;
// Interconnect Declarations for Component Instantiations
  assign chn_inp_out_rsci_bawt = chn_inp_out_rsci_biwt | chn_inp_out_rsci_bcwt;
  assign chn_inp_out_rsci_wen_comp = (~ chn_inp_out_rsci_oswt) | chn_inp_out_rsci_bawt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_out_rsci_bcwt <= 1'b0;
    end
    else begin
      chn_inp_out_rsci_bcwt <= ~((~(chn_inp_out_rsci_bcwt | chn_inp_out_rsci_biwt))
          | chn_inp_out_rsci_bdwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_out_rsci_chn_inp_out_wait_ctrl
// ------------------------------------------------------------------
module NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_out_rsci_chn_inp_out_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_inp_out_rsci_oswt, core_wen, core_wten, chn_inp_out_rsci_iswt0,
      chn_inp_out_rsci_ld_core_psct, chn_inp_out_rsci_biwt, chn_inp_out_rsci_bdwt,
      chn_inp_out_rsci_ld_core_sct, chn_inp_out_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_inp_out_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_inp_out_rsci_iswt0;
  input chn_inp_out_rsci_ld_core_psct;
  output chn_inp_out_rsci_biwt;
  output chn_inp_out_rsci_bdwt;
  output chn_inp_out_rsci_ld_core_sct;
  input chn_inp_out_rsci_vd;
// Interconnect Declarations
  wire chn_inp_out_rsci_ogwt;
  wire chn_inp_out_rsci_pdswt0;
  reg chn_inp_out_rsci_icwt;
// Interconnect Declarations for Component Instantiations
  assign chn_inp_out_rsci_pdswt0 = (~ core_wten) & chn_inp_out_rsci_iswt0;
  assign chn_inp_out_rsci_biwt = chn_inp_out_rsci_ogwt & chn_inp_out_rsci_vd;
  assign chn_inp_out_rsci_ogwt = chn_inp_out_rsci_pdswt0 | chn_inp_out_rsci_icwt;
  assign chn_inp_out_rsci_bdwt = chn_inp_out_rsci_oswt & core_wen;
  assign chn_inp_out_rsci_ld_core_sct = chn_inp_out_rsci_ld_core_psct & chn_inp_out_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_out_rsci_icwt <= 1'b0;
    end
    else begin
      chn_inp_out_rsci_icwt <= ~((~(chn_inp_out_rsci_icwt | chn_inp_out_rsci_pdswt0))
          | chn_inp_out_rsci_biwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_in_rsci_chn_inp_in_wait_dp
// ------------------------------------------------------------------
module NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_in_rsci_chn_inp_in_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_inp_in_rsci_oswt, chn_inp_in_rsci_bawt, chn_inp_in_rsci_wen_comp,
      chn_inp_in_rsci_d_mxwt, chn_inp_in_rsci_biwt, chn_inp_in_rsci_bdwt, chn_inp_in_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_inp_in_rsci_oswt;
  output chn_inp_in_rsci_bawt;
  output chn_inp_in_rsci_wen_comp;
  output [739:0] chn_inp_in_rsci_d_mxwt;
  input chn_inp_in_rsci_biwt;
  input chn_inp_in_rsci_bdwt;
  input [739:0] chn_inp_in_rsci_d;
// Interconnect Declarations
  reg chn_inp_in_rsci_bcwt;
  reg [739:0] chn_inp_in_rsci_d_bfwt;
// Interconnect Declarations for Component Instantiations
  assign chn_inp_in_rsci_bawt = chn_inp_in_rsci_biwt | chn_inp_in_rsci_bcwt;
  assign chn_inp_in_rsci_wen_comp = (~ chn_inp_in_rsci_oswt) | chn_inp_in_rsci_bawt;
  assign chn_inp_in_rsci_d_mxwt = MUX_v_740_2_2(chn_inp_in_rsci_d, chn_inp_in_rsci_d_bfwt,
      chn_inp_in_rsci_bcwt);
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_rsci_bcwt <= 1'b0;
      chn_inp_in_rsci_d_bfwt <= 740'b0;
    end
    else begin
      chn_inp_in_rsci_bcwt <= ~((~(chn_inp_in_rsci_bcwt | chn_inp_in_rsci_biwt))
          | chn_inp_in_rsci_bdwt);
      chn_inp_in_rsci_d_bfwt <= chn_inp_in_rsci_d_mxwt;
    end
  end
  function [739:0] MUX_v_740_2_2;
    input [739:0] input_0;
    input [739:0] input_1;
    input [0:0] sel;
    reg [739:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_740_2_2 = result;
  end
  endfunction
endmodule
// ------------------------------------------------------------------
// Design Unit: NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_in_rsci_chn_inp_in_wait_ctrl
// ------------------------------------------------------------------
module NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_in_rsci_chn_inp_in_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_inp_in_rsci_oswt, core_wen, chn_inp_in_rsci_iswt0,
      chn_inp_in_rsci_ld_core_psct, core_wten, chn_inp_in_rsci_biwt, chn_inp_in_rsci_bdwt,
      chn_inp_in_rsci_ld_core_sct, chn_inp_in_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_inp_in_rsci_oswt;
  input core_wen;
  input chn_inp_in_rsci_iswt0;
  input chn_inp_in_rsci_ld_core_psct;
  input core_wten;
  output chn_inp_in_rsci_biwt;
  output chn_inp_in_rsci_bdwt;
  output chn_inp_in_rsci_ld_core_sct;
  input chn_inp_in_rsci_vd;
// Interconnect Declarations
  wire chn_inp_in_rsci_ogwt;
  wire chn_inp_in_rsci_pdswt0;
  reg chn_inp_in_rsci_icwt;
// Interconnect Declarations for Component Instantiations
  assign chn_inp_in_rsci_pdswt0 = (~ core_wten) & chn_inp_in_rsci_iswt0;
  assign chn_inp_in_rsci_biwt = chn_inp_in_rsci_ogwt & chn_inp_in_rsci_vd;
  assign chn_inp_in_rsci_ogwt = chn_inp_in_rsci_pdswt0 | chn_inp_in_rsci_icwt;
  assign chn_inp_in_rsci_bdwt = chn_inp_in_rsci_oswt & core_wen;
  assign chn_inp_in_rsci_ld_core_sct = chn_inp_in_rsci_ld_core_psct & chn_inp_in_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_rsci_icwt <= 1'b0;
    end
    else begin
      chn_inp_in_rsci_icwt <= ~((~(chn_inp_in_rsci_icwt | chn_inp_in_rsci_pdswt0))
          | chn_inp_in_rsci_biwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_out_rsci
// ------------------------------------------------------------------
module NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_out_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_inp_out_rsc_z, chn_inp_out_rsc_vz, chn_inp_out_rsc_lz,
      chn_inp_out_rsci_oswt, core_wen, core_wten, chn_inp_out_rsci_iswt0, chn_inp_out_rsci_bawt,
      chn_inp_out_rsci_wen_comp, chn_inp_out_rsci_ld_core_psct, chn_inp_out_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output [127:0] chn_inp_out_rsc_z;
  input chn_inp_out_rsc_vz;
  output chn_inp_out_rsc_lz;
  input chn_inp_out_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_inp_out_rsci_iswt0;
  output chn_inp_out_rsci_bawt;
  output chn_inp_out_rsci_wen_comp;
  input chn_inp_out_rsci_ld_core_psct;
  input [127:0] chn_inp_out_rsci_d;
// Interconnect Declarations
  wire chn_inp_out_rsci_biwt;
  wire chn_inp_out_rsci_bdwt;
  wire chn_inp_out_rsci_ld_core_sct;
  wire chn_inp_out_rsci_vd;
// Interconnect Declarations for Component Instantiations
  SDP_Y_INP_mgc_out_stdreg_wait_v1 #(.rscid(32'sd3),
  .width(32'sd128)) chn_inp_out_rsci (
      .ld(chn_inp_out_rsci_ld_core_sct),
      .vd(chn_inp_out_rsci_vd),
      .d(chn_inp_out_rsci_d),
      .lz(chn_inp_out_rsc_lz),
      .vz(chn_inp_out_rsc_vz),
      .z(chn_inp_out_rsc_z)
    );
  NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_out_rsci_chn_inp_out_wait_ctrl NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_out_rsci_chn_inp_out_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_inp_out_rsci_oswt(chn_inp_out_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_inp_out_rsci_iswt0(chn_inp_out_rsci_iswt0),
      .chn_inp_out_rsci_ld_core_psct(chn_inp_out_rsci_ld_core_psct),
      .chn_inp_out_rsci_biwt(chn_inp_out_rsci_biwt),
      .chn_inp_out_rsci_bdwt(chn_inp_out_rsci_bdwt),
      .chn_inp_out_rsci_ld_core_sct(chn_inp_out_rsci_ld_core_sct),
      .chn_inp_out_rsci_vd(chn_inp_out_rsci_vd)
    );
  NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_out_rsci_chn_inp_out_wait_dp NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_out_rsci_chn_inp_out_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_inp_out_rsci_oswt(chn_inp_out_rsci_oswt),
      .chn_inp_out_rsci_bawt(chn_inp_out_rsci_bawt),
      .chn_inp_out_rsci_wen_comp(chn_inp_out_rsci_wen_comp),
      .chn_inp_out_rsci_biwt(chn_inp_out_rsci_biwt),
      .chn_inp_out_rsci_bdwt(chn_inp_out_rsci_bdwt)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_in_rsci
// ------------------------------------------------------------------
module NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_in_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_inp_in_rsc_z, chn_inp_in_rsc_vz, chn_inp_in_rsc_lz,
      chn_inp_in_rsci_oswt, core_wen, chn_inp_in_rsci_iswt0, chn_inp_in_rsci_bawt,
      chn_inp_in_rsci_wen_comp, chn_inp_in_rsci_ld_core_psct, chn_inp_in_rsci_d_mxwt,
      core_wten
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [739:0] chn_inp_in_rsc_z;
  input chn_inp_in_rsc_vz;
  output chn_inp_in_rsc_lz;
  input chn_inp_in_rsci_oswt;
  input core_wen;
  input chn_inp_in_rsci_iswt0;
  output chn_inp_in_rsci_bawt;
  output chn_inp_in_rsci_wen_comp;
  input chn_inp_in_rsci_ld_core_psct;
  output [739:0] chn_inp_in_rsci_d_mxwt;
  input core_wten;
// Interconnect Declarations
  wire chn_inp_in_rsci_biwt;
  wire chn_inp_in_rsci_bdwt;
  wire chn_inp_in_rsci_ld_core_sct;
  wire chn_inp_in_rsci_vd;
  wire [739:0] chn_inp_in_rsci_d;
// Interconnect Declarations for Component Instantiations
  SDP_Y_INP_mgc_in_wire_wait_v1 #(.rscid(32'sd1),
  .width(32'sd740)) chn_inp_in_rsci (
      .ld(chn_inp_in_rsci_ld_core_sct),
      .vd(chn_inp_in_rsci_vd),
      .d(chn_inp_in_rsci_d),
      .lz(chn_inp_in_rsc_lz),
      .vz(chn_inp_in_rsc_vz),
      .z(chn_inp_in_rsc_z)
    );
  NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_in_rsci_chn_inp_in_wait_ctrl NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_in_rsci_chn_inp_in_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_inp_in_rsci_oswt(chn_inp_in_rsci_oswt),
      .core_wen(core_wen),
      .chn_inp_in_rsci_iswt0(chn_inp_in_rsci_iswt0),
      .chn_inp_in_rsci_ld_core_psct(chn_inp_in_rsci_ld_core_psct),
      .core_wten(core_wten),
      .chn_inp_in_rsci_biwt(chn_inp_in_rsci_biwt),
      .chn_inp_in_rsci_bdwt(chn_inp_in_rsci_bdwt),
      .chn_inp_in_rsci_ld_core_sct(chn_inp_in_rsci_ld_core_sct),
      .chn_inp_in_rsci_vd(chn_inp_in_rsci_vd)
    );
  NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_in_rsci_chn_inp_in_wait_dp NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_in_rsci_chn_inp_in_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_inp_in_rsci_oswt(chn_inp_in_rsci_oswt),
      .chn_inp_in_rsci_bawt(chn_inp_in_rsci_bawt),
      .chn_inp_in_rsci_wen_comp(chn_inp_in_rsci_wen_comp),
      .chn_inp_in_rsci_d_mxwt(chn_inp_in_rsci_d_mxwt),
      .chn_inp_in_rsci_biwt(chn_inp_in_rsci_biwt),
      .chn_inp_in_rsci_bdwt(chn_inp_in_rsci_bdwt),
      .chn_inp_in_rsci_d(chn_inp_in_rsci_d)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: NV_NVDLA_SDP_CORE_Y_inp_core
// ------------------------------------------------------------------
module NV_NVDLA_SDP_CORE_Y_inp_core (
  nvdla_core_clk, nvdla_core_rstn, chn_inp_in_rsc_z, chn_inp_in_rsc_vz, chn_inp_in_rsc_lz,
      cfg_precision_rsc_z, chn_inp_out_rsc_z, chn_inp_out_rsc_vz, chn_inp_out_rsc_lz,
      chn_inp_in_rsci_oswt, chn_inp_in_rsci_oswt_unreg, chn_inp_out_rsci_oswt, chn_inp_out_rsci_oswt_unreg
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [739:0] chn_inp_in_rsc_z;
  input chn_inp_in_rsc_vz;
  output chn_inp_in_rsc_lz;
  input [1:0] cfg_precision_rsc_z;
  output [127:0] chn_inp_out_rsc_z;
  input chn_inp_out_rsc_vz;
  output chn_inp_out_rsc_lz;
  input chn_inp_in_rsci_oswt;
  output chn_inp_in_rsci_oswt_unreg;
  input chn_inp_out_rsci_oswt;
  output chn_inp_out_rsci_oswt_unreg;
// Interconnect Declarations
  wire core_wen;
  reg chn_inp_in_rsci_iswt0;
  wire chn_inp_in_rsci_bawt;
  wire chn_inp_in_rsci_wen_comp;
  reg chn_inp_in_rsci_ld_core_psct;
  wire [739:0] chn_inp_in_rsci_d_mxwt;
  wire core_wten;
  wire [1:0] cfg_precision_rsci_d;
  reg chn_inp_out_rsci_iswt0;
  wire chn_inp_out_rsci_bawt;
  wire chn_inp_out_rsci_wen_comp;
  reg chn_inp_out_rsci_d_127;
  reg [2:0] chn_inp_out_rsci_d_126_124;
  reg [9:0] chn_inp_out_rsci_d_118_109;
  reg [2:0] chn_inp_out_rsci_d_108_106;
  reg [8:0] chn_inp_out_rsci_d_105_97;
  reg chn_inp_out_rsci_d_96;
  reg chn_inp_out_rsci_d_95;
  reg [2:0] chn_inp_out_rsci_d_94_92;
  reg [9:0] chn_inp_out_rsci_d_86_77;
  reg [2:0] chn_inp_out_rsci_d_76_74;
  reg [8:0] chn_inp_out_rsci_d_73_65;
  reg chn_inp_out_rsci_d_64;
  reg chn_inp_out_rsci_d_63;
  reg [2:0] chn_inp_out_rsci_d_62_60;
  reg [9:0] chn_inp_out_rsci_d_54_45;
  reg [2:0] chn_inp_out_rsci_d_44_42;
  reg [8:0] chn_inp_out_rsci_d_41_33;
  reg chn_inp_out_rsci_d_32;
  reg chn_inp_out_rsci_d_31;
  reg [2:0] chn_inp_out_rsci_d_30_28;
  reg [9:0] chn_inp_out_rsci_d_22_13;
  reg [2:0] chn_inp_out_rsci_d_12_10;
  reg [8:0] chn_inp_out_rsci_d_9_1;
  reg chn_inp_out_rsci_d_0;
  reg chn_inp_out_rsci_d_123;
  reg [3:0] chn_inp_out_rsci_d_122_119;
  reg chn_inp_out_rsci_d_91;
  reg [3:0] chn_inp_out_rsci_d_90_87;
  reg chn_inp_out_rsci_d_59;
  reg [3:0] chn_inp_out_rsci_d_58_55;
  reg chn_inp_out_rsci_d_27;
  reg [3:0] chn_inp_out_rsci_d_26_23;
  wire [1:0] fsm_output;
  wire IsDenorm_5U_10U_or_3_tmp;
  wire IsDenorm_5U_10U_3_or_3_tmp;
  wire IsDenorm_5U_10U_2_or_3_tmp;
  wire inp_lookup_4_FpMantRNE_36U_11U_1_else_and_tmp;
  wire IsDenorm_5U_10U_or_2_tmp;
  wire IsDenorm_5U_10U_3_or_2_tmp;
  wire IsDenorm_5U_10U_2_or_2_tmp;
  wire inp_lookup_3_FpMantRNE_36U_11U_1_else_and_tmp;
  wire IsDenorm_5U_10U_or_1_tmp;
  wire IsDenorm_5U_10U_3_or_1_tmp;
  wire IsDenorm_5U_10U_2_or_1_tmp;
  wire inp_lookup_2_FpMantRNE_36U_11U_1_else_and_tmp;
  wire IsDenorm_5U_10U_or_tmp;
  wire IsNaN_8U_23U_nor_tmp;
  wire IsDenorm_5U_10U_3_or_tmp;
  wire IsDenorm_5U_10U_2_or_tmp;
  wire inp_lookup_1_FpMantRNE_36U_11U_1_else_and_tmp;
  wire IsNaN_6U_10U_6_nor_3_tmp;
  wire FpMul_6U_10U_2_if_2_FpMul_6U_10U_2_if_2_or_7_tmp;
  wire [4:0] FpFractionToFloat_35U_6U_10U_1_mux_42_tmp;
  wire inp_lookup_4_FpMantRNE_36U_11U_else_and_tmp;
  wire IsNaN_6U_10U_6_nor_2_tmp;
  wire FpMul_6U_10U_2_if_2_FpMul_6U_10U_2_if_2_or_5_tmp;
  wire [4:0] FpFractionToFloat_35U_6U_10U_1_mux_41_tmp;
  wire inp_lookup_3_FpMantRNE_36U_11U_else_and_tmp;
  wire IsNaN_6U_10U_6_nor_1_tmp;
  wire [4:0] FpFractionToFloat_35U_6U_10U_1_mux_40_tmp;
  wire inp_lookup_2_FpMantRNE_36U_11U_else_and_tmp;
  wire IsNaN_6U_10U_6_nor_tmp;
  wire [4:0] FpFractionToFloat_35U_6U_10U_1_mux_tmp;
  wire inp_lookup_1_FpMantRNE_36U_11U_else_and_tmp;
  wire FpNormalize_8U_49U_if_FpNormalize_8U_49U_if_nand_3_tmp;
  wire [21:0] inp_lookup_4_FpMul_6U_10U_2_p_mant_p1_mul_tmp;
  wire IsNaN_6U_10U_4_nor_3_tmp;
  wire FpMul_6U_10U_1_if_2_FpMul_6U_10U_1_if_2_or_6_tmp;
  wire FpNormalize_8U_49U_if_FpNormalize_8U_49U_if_nand_2_tmp;
  wire [21:0] inp_lookup_3_FpMul_6U_10U_2_p_mant_p1_mul_tmp;
  wire IsNaN_6U_10U_4_nor_2_tmp;
  wire FpMul_6U_10U_1_if_2_FpMul_6U_10U_1_if_2_or_4_tmp;
  wire FpNormalize_8U_49U_if_FpNormalize_8U_49U_if_nand_1_tmp;
  wire [21:0] inp_lookup_2_FpMul_6U_10U_2_p_mant_p1_mul_tmp;
  wire IsNaN_6U_10U_4_nor_1_tmp;
  wire FpMul_6U_10U_1_if_2_FpMul_6U_10U_1_if_2_or_2_tmp;
  wire FpNormalize_8U_49U_if_FpNormalize_8U_49U_if_nand_tmp;
  wire [21:0] inp_lookup_1_FpMul_6U_10U_2_p_mant_p1_mul_tmp;
  wire IsNaN_6U_10U_4_nor_tmp;
  wire FpMul_6U_10U_1_if_2_FpMul_6U_10U_1_if_2_or_tmp;
  wire inp_lookup_4_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp;
  wire inp_lookup_4_FpMantRNE_49U_24U_else_and_tmp;
  wire [21:0] inp_lookup_4_FpMul_6U_10U_1_p_mant_p1_mul_tmp;
  wire inp_lookup_3_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp;
  wire inp_lookup_3_FpMantRNE_49U_24U_else_and_tmp;
  wire [21:0] inp_lookup_3_FpMul_6U_10U_1_p_mant_p1_mul_tmp;
  wire inp_lookup_2_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp;
  wire inp_lookup_2_FpMantRNE_49U_24U_else_and_tmp;
  wire [21:0] inp_lookup_2_FpMul_6U_10U_1_p_mant_p1_mul_tmp;
  wire inp_lookup_1_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp;
  wire inp_lookup_1_FpMantRNE_49U_24U_else_and_tmp;
  wire [21:0] inp_lookup_1_FpMul_6U_10U_1_p_mant_p1_mul_tmp;
  wire IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_3_tmp;
  wire IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_2_tmp;
  wire IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_1_tmp;
  wire IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_tmp;
  wire inp_lookup_4_FpMantRNE_49U_24U_1_else_and_tmp;
  wire inp_lookup_3_FpMantRNE_49U_24U_1_else_and_tmp;
  wire inp_lookup_2_FpMantRNE_49U_24U_1_else_and_tmp;
  wire inp_lookup_1_FpMantRNE_49U_24U_1_else_and_tmp;
  wire IsNaN_6U_10U_IsNaN_6U_10U_nor_3_tmp;
  wire FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_6_tmp;
  wire inp_lookup_4_FpMantRNE_23U_11U_1_else_and_tmp;
  wire IsNaN_6U_10U_IsNaN_6U_10U_nor_2_tmp;
  wire FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_4_tmp;
  wire inp_lookup_3_FpMantRNE_23U_11U_1_else_and_tmp;
  wire IsNaN_6U_10U_IsNaN_6U_10U_nor_1_tmp;
  wire FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_2_tmp;
  wire inp_lookup_2_FpMantRNE_23U_11U_1_else_and_tmp;
  wire IsNaN_6U_10U_IsNaN_6U_10U_nor_tmp;
  wire FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_tmp;
  wire inp_lookup_1_FpMantRNE_23U_11U_1_else_and_tmp;
  wire inp_lookup_4_FpAdd_6U_10U_is_a_greater_oif_equal_tmp;
  wire inp_lookup_3_FpAdd_6U_10U_is_a_greater_oif_equal_tmp;
  wire inp_lookup_2_FpAdd_6U_10U_is_a_greater_oif_equal_tmp;
  wire inp_lookup_1_FpAdd_6U_10U_is_a_greater_oif_equal_tmp;
  wire IsNaN_6U_23U_IsNaN_6U_23U_nor_3_tmp;
  wire inp_lookup_4_FpMantRNE_23U_11U_else_and_tmp;
  wire IsNaN_6U_23U_IsNaN_6U_23U_nor_2_tmp;
  wire inp_lookup_3_FpMantRNE_23U_11U_else_and_tmp;
  wire IsNaN_6U_23U_IsNaN_6U_23U_nor_1_tmp;
  wire inp_lookup_2_FpMantRNE_23U_11U_else_and_tmp;
  wire IsNaN_6U_23U_IsNaN_6U_23U_nor_tmp;
  wire inp_lookup_1_FpMantRNE_23U_11U_else_and_tmp;
  wire inp_lookup_4_FpMantRNE_22U_11U_2_else_and_tmp;
  wire inp_lookup_3_FpMantRNE_22U_11U_2_else_and_tmp;
  wire inp_lookup_2_FpMantRNE_22U_11U_2_else_and_tmp;
  wire inp_lookup_1_FpMantRNE_22U_11U_2_else_and_tmp;
  wire inp_lookup_4_FpMantRNE_22U_11U_1_else_and_tmp;
  wire inp_lookup_3_FpMantRNE_22U_11U_1_else_and_tmp;
  wire inp_lookup_2_FpMantRNE_22U_11U_1_else_and_tmp;
  wire inp_lookup_1_FpMantRNE_22U_11U_1_else_and_tmp;
  wire inp_lookup_4_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp;
  wire inp_lookup_3_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp;
  wire inp_lookup_2_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp;
  wire inp_lookup_1_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp;
  wire IsNaN_8U_23U_4_IsNaN_8U_23U_4_nor_3_tmp;
  wire IsNaN_8U_23U_4_IsNaN_8U_23U_4_nor_2_tmp;
  wire IsNaN_8U_23U_4_IsNaN_8U_23U_4_nor_1_tmp;
  wire IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_tmp;
  wire IsNaN_8U_23U_4_nor_tmp;
  wire [21:0] inp_lookup_4_FpMul_6U_10U_p_mant_p1_mul_tmp;
  wire [21:0] inp_lookup_3_FpMul_6U_10U_p_mant_p1_mul_tmp;
  wire [21:0] inp_lookup_2_FpMul_6U_10U_p_mant_p1_mul_tmp;
  wire [21:0] inp_lookup_1_FpMul_6U_10U_p_mant_p1_mul_tmp;
  wire FpNormalize_6U_23U_if_FpNormalize_6U_23U_if_nand_3_tmp;
  wire FpNormalize_6U_23U_if_FpNormalize_6U_23U_if_nand_2_tmp;
  wire FpNormalize_6U_23U_if_FpNormalize_6U_23U_if_nand_1_tmp;
  wire FpNormalize_6U_23U_if_FpNormalize_6U_23U_if_nand_tmp;
  wire inp_lookup_4_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_tmp;
  wire inp_lookup_3_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_tmp;
  wire inp_lookup_2_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_tmp;
  wire inp_lookup_1_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_tmp;
  wire inp_lookup_3_IsNaN_6U_10U_7_aif_IsNaN_6U_10U_7_aelse_IsNaN_6U_10U_7_aelse_or_tmp;
  wire IsNaN_8U_23U_3_IsNaN_8U_23U_3_nand_3_tmp;
  wire IsNaN_8U_23U_3_nor_3_tmp;
  wire IsNaN_8U_23U_3_IsNaN_8U_23U_3_nor_2_tmp;
  wire IsNaN_8U_23U_3_IsNaN_8U_23U_3_nor_1_tmp;
  wire IsNaN_8U_23U_3_IsNaN_8U_23U_3_nor_tmp;
  wire inp_lookup_4_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp;
  wire inp_lookup_3_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp;
  wire inp_lookup_2_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp;
  wire inp_lookup_1_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp;
  wire IsNaN_6U_10U_3_IsNaN_6U_10U_3_nor_3_tmp;
  wire IsNaN_6U_10U_3_IsNaN_6U_10U_3_nor_2_tmp;
  wire IsNaN_6U_10U_3_IsNaN_6U_10U_3_nor_1_tmp;
  wire IsNaN_6U_10U_3_IsNaN_6U_10U_3_nor_tmp;
  wire IsNaN_6U_10U_9_nor_3_tmp;
  wire IsNaN_6U_10U_9_nor_2_tmp;
  wire IsNaN_6U_10U_9_nor_1_tmp;
  wire IsNaN_6U_10U_9_nor_tmp;
  wire and_dcpl_21;
  wire and_dcpl_38;
  wire and_dcpl_40;
  wire and_dcpl_42;
  wire and_dcpl_49;
  wire and_dcpl_57;
  wire and_dcpl_65;
  wire or_tmp_6;
  wire or_tmp_8;
  wire not_tmp_34;
  wire or_tmp_21;
  wire mux_tmp_6;
  wire not_tmp_45;
  wire or_tmp_52;
  wire or_tmp_85;
  wire not_tmp_69;
  wire or_tmp_114;
  wire nand_tmp_3;
  wire not_tmp_101;
  wire mux_tmp_50;
  wire nand_tmp_5;
  wire or_tmp_213;
  wire or_tmp_234;
  wire or_tmp_238;
  wire or_tmp_241;
  wire not_tmp_126;
  wire nand_tmp_8;
  wire or_tmp_277;
  wire or_tmp_306;
  wire not_tmp_152;
  wire nand_tmp_12;
  wire or_tmp_347;
  wire or_tmp_374;
  wire or_tmp_439;
  wire and_tmp_29;
  wire or_tmp_440;
  wire not_tmp_182;
  wire and_tmp_33;
  wire mux_tmp_127;
  wire mux_tmp_133;
  wire or_tmp_461;
  wire nand_tmp_14;
  wire and_tmp_34;
  wire or_tmp_463;
  wire and_tmp_35;
  wire mux_tmp_163;
  wire and_tmp_38;
  wire mux_tmp_165;
  wire mux_tmp_171;
  wire or_tmp_523;
  wire nand_tmp_16;
  wire and_tmp_39;
  wire or_tmp_525;
  wire and_tmp_42;
  wire mux_tmp_201;
  wire and_tmp_45;
  wire mux_tmp_203;
  wire mux_tmp_209;
  wire or_tmp_584;
  wire and_tmp_48;
  wire nand_tmp_18;
  wire or_tmp_597;
  wire nand_tmp_20;
  wire and_tmp_49;
  wire or_tmp_599;
  wire or_tmp_621;
  wire and_tmp_50;
  wire or_tmp_630;
  wire or_tmp_631;
  wire mux_tmp_247;
  wire mux_tmp_250;
  wire mux_tmp_251;
  wire nand_tmp_24;
  wire mux_tmp_260;
  wire mux_tmp_262;
  wire mux_tmp_278;
  wire or_tmp_679;
  wire not_tmp_282;
  wire or_tmp_701;
  wire nand_tmp_29;
  wire and_tmp_54;
  wire or_tmp_704;
  wire or_tmp_736;
  wire or_tmp_753;
  wire nand_tmp_37;
  wire and_tmp_56;
  wire or_tmp_756;
  wire not_tmp_345;
  wire or_tmp_792;
  wire not_tmp_346;
  wire or_tmp_798;
  wire or_tmp_808;
  wire nand_tmp_45;
  wire and_tmp_59;
  wire or_tmp_811;
  wire nand_tmp_47;
  wire nand_tmp_50;
  wire not_tmp_374;
  wire or_tmp_850;
  wire or_tmp_880;
  wire nand_tmp_53;
  wire or_tmp_899;
  wire or_tmp_945;
  wire or_tmp_957;
  wire or_tmp_959;
  wire not_tmp_424;
  wire or_tmp_962;
  wire mux_tmp_441;
  wire mux_tmp_444;
  wire not_tmp_428;
  wire or_tmp_990;
  wire or_tmp_992;
  wire mux_tmp_454;
  wire mux_tmp_457;
  wire or_tmp_1009;
  wire not_tmp_442;
  wire mux_tmp_465;
  wire mux_tmp_467;
  wire or_tmp_1038;
  wire mux_tmp_475;
  wire mux_tmp_478;
  wire or_tmp_1058;
  wire or_tmp_1060;
  wire nor_tmp_139;
  wire or_tmp_1098;
  wire or_tmp_1106;
  wire nor_tmp_146;
  wire or_tmp_1143;
  wire or_tmp_1147;
  wire or_tmp_1151;
  wire or_tmp_1182;
  wire or_tmp_1185;
  wire or_tmp_1198;
  wire or_tmp_1232;
  wire or_tmp_1239;
  wire or_tmp_1253;
  wire or_tmp_1255;
  wire nor_tmp_161;
  wire nor_tmp_166;
  wire not_tmp_537;
  wire or_tmp_1302;
  wire or_tmp_1310;
  wire or_tmp_1312;
  wire nor_tmp_172;
  wire not_tmp_546;
  wire or_tmp_1338;
  wire or_tmp_1340;
  wire nor_tmp_176;
  wire or_tmp_1363;
  wire or_tmp_1369;
  wire or_tmp_1389;
  wire or_tmp_1393;
  wire or_tmp_1399;
  wire or_tmp_1418;
  wire or_tmp_1422;
  wire or_tmp_1428;
  wire or_tmp_1444;
  wire or_tmp_1448;
  wire or_tmp_1454;
  wire or_tmp_1467;
  wire or_tmp_1502;
  wire nor_tmp_199;
  wire or_tmp_1537;
  wire nor_tmp_208;
  wire nor_tmp_216;
  wire nor_tmp_224;
  wire not_tmp_698;
  wire nor_tmp_227;
  wire not_tmp_703;
  wire nor_tmp_230;
  wire not_tmp_708;
  wire nor_tmp_232;
  wire not_tmp_711;
  wire nor_tmp_234;
  wire mux_tmp_698;
  wire or_tmp_1661;
  wire or_tmp_1665;
  wire or_tmp_1671;
  wire or_tmp_1687;
  wire mux_tmp_708;
  wire or_tmp_1690;
  wire or_tmp_1697;
  wire or_tmp_1699;
  wire or_tmp_1701;
  wire mux_tmp_715;
  wire or_tmp_1724;
  wire or_tmp_1728;
  wire or_tmp_1734;
  wire not_tmp_733;
  wire or_tmp_1736;
  wire or_tmp_1741;
  wire or_tmp_1770;
  wire or_tmp_1774;
  wire or_tmp_1784;
  wire or_tmp_1786;
  wire or_tmp_1806;
  wire mux_tmp_754;
  wire or_tmp_1818;
  wire nor_tmp_250;
  wire or_tmp_1826;
  wire nor_tmp_252;
  wire or_tmp_1840;
  wire nor_tmp_253;
  wire or_tmp_1845;
  wire or_tmp_1849;
  wire nor_tmp_256;
  wire or_tmp_1856;
  wire not_tmp_772;
  wire not_tmp_773;
  wire nand_tmp_90;
  wire not_tmp_776;
  wire or_tmp_1891;
  wire and_tmp_111;
  wire nand_tmp_91;
  wire not_tmp_789;
  wire not_tmp_790;
  wire nand_tmp_94;
  wire not_tmp_793;
  wire or_tmp_1929;
  wire and_tmp_116;
  wire nand_tmp_95;
  wire not_tmp_806;
  wire not_tmp_807;
  wire nand_tmp_98;
  wire not_tmp_810;
  wire or_tmp_1967;
  wire and_tmp_121;
  wire nand_tmp_99;
  wire or_tmp_2199;
  wire or_tmp_2234;
  wire not_tmp_940;
  wire mux_tmp_950;
  wire mux_tmp_966;
  wire mux_tmp_967;
  wire nand_tmp_126;
  wire or_tmp_2441;
  wire or_tmp_2486;
  wire or_tmp_2490;
  wire or_tmp_2494;
  wire or_tmp_2498;
  wire mux_tmp_1008;
  wire not_tmp_1029;
  wire and_tmp_158;
  wire mux_tmp_1015;
  wire or_tmp_2531;
  wire nand_tmp_138;
  wire mux_tmp_1025;
  wire not_tmp_1046;
  wire and_tmp_162;
  wire mux_tmp_1032;
  wire nand_tmp_142;
  wire mux_tmp_1042;
  wire not_tmp_1063;
  wire and_tmp_166;
  wire mux_tmp_1049;
  wire nand_tmp_146;
  wire mux_tmp_1059;
  wire not_tmp_1080;
  wire mux_tmp_1067;
  wire or_tmp_2643;
  wire nand_tmp_148;
  wire or_tmp_2695;
  wire not_tmp_1108;
  wire mux_tmp_1092;
  wire or_tmp_2703;
  wire or_tmp_2710;
  wire or_tmp_2717;
  wire or_tmp_2723;
  wire or_tmp_2738;
  wire or_tmp_2768;
  wire or_tmp_2804;
  wire nand_tmp_162;
  wire nand_tmp_163;
  wire nand_tmp_164;
  wire nand_tmp_165;
  wire or_tmp_2924;
  wire or_tmp_2935;
  wire not_tmp_1202;
  wire or_tmp_2953;
  wire not_tmp_1208;
  wire or_tmp_2974;
  wire not_tmp_1212;
  wire and_tmp_181;
  wire mux_tmp_1183;
  wire and_tmp_182;
  wire or_tmp_2986;
  wire mux_tmp_1187;
  wire and_tmp_184;
  wire or_tmp_2990;
  wire and_tmp_187;
  wire or_tmp_2993;
  wire mux_tmp_1195;
  wire and_tmp_188;
  wire or_tmp_2997;
  wire or_tmp_2999;
  wire or_tmp_3002;
  wire or_tmp_3007;
  wire or_tmp_3011;
  wire mux_tmp_1209;
  wire or_tmp_3017;
  wire or_tmp_3020;
  wire or_tmp_3025;
  wire or_tmp_3029;
  wire mux_tmp_1221;
  wire or_tmp_3035;
  wire or_tmp_3038;
  wire or_tmp_3043;
  wire or_tmp_3047;
  wire mux_tmp_1233;
  wire or_tmp_3053;
  wire or_tmp_3056;
  wire or_tmp_3061;
  wire or_tmp_3065;
  wire mux_tmp_1245;
  wire or_tmp_3087;
  wire or_tmp_3123;
  wire or_tmp_3132;
  wire or_tmp_3152;
  wire or_tmp_3153;
  wire or_tmp_3156;
  wire or_tmp_3160;
  wire or_tmp_3180;
  wire or_tmp_3200;
  wire or_tmp_3224;
  wire or_tmp_3227;
  wire or_tmp_3230;
  wire or_tmp_3233;
  wire or_tmp_3235;
  wire or_tmp_3246;
  wire or_tmp_3257;
  wire or_tmp_3268;
  wire not_tmp_1369;
  wire nor_tmp_464;
  wire not_tmp_1373;
  wire not_tmp_1377;
  wire not_tmp_1381;
  wire mux_tmp_1367;
  wire not_tmp_1388;
  wire not_tmp_1391;
  wire not_tmp_1425;
  wire mux_tmp_1450;
  wire mux_tmp_1452;
  wire mux_tmp_1454;
  wire mux_tmp_1458;
  wire or_tmp_3510;
  wire or_tmp_3512;
  wire or_tmp_3514;
  wire or_tmp_3516;
  wire mux_tmp_1485;
  wire mux_tmp_1488;
  wire mux_tmp_1494;
  wire nor_tmp_522;
  wire or_tmp_3530;
  wire or_tmp_3534;
  wire or_tmp_3538;
  wire or_tmp_3542;
  wire nor_tmp_532;
  wire nor_tmp_533;
  wire nor_tmp_535;
  wire mux_tmp_1509;
  wire mux_tmp_1511;
  wire mux_tmp_1513;
  wire mux_tmp_1518;
  wire nor_tmp_545;
  wire or_tmp_3562;
  wire or_tmp_3564;
  wire or_tmp_3566;
  wire or_tmp_3568;
  wire nor_tmp_551;
  wire nor_tmp_552;
  wire nor_tmp_553;
  wire nor_tmp_555;
  wire or_tmp_3612;
  wire or_tmp_3614;
  wire or_tmp_3616;
  wire or_tmp_3618;
  wire nor_tmp_560;
  wire mux_tmp_1543;
  wire mux_tmp_1545;
  wire mux_tmp_1548;
  wire mux_tmp_1553;
  wire nor_tmp_569;
  wire or_tmp_3627;
  wire or_tmp_3629;
  wire or_tmp_3631;
  wire or_tmp_3633;
  wire and_tmp_225;
  wire and_tmp_226;
  wire and_tmp_227;
  wire and_tmp_228;
  wire not_tmp_1550;
  wire mux_tmp_1573;
  wire mux_tmp_1575;
  wire mux_tmp_1577;
  wire mux_tmp_1579;
  wire mux_tmp_1581;
  wire mux_tmp_1583;
  wire mux_tmp_1585;
  wire mux_tmp_1587;
  wire nand_tmp_218;
  wire nand_tmp_219;
  wire nand_tmp_220;
  wire nand_tmp_221;
  wire nand_tmp_222;
  wire or_tmp_3798;
  wire or_tmp_3802;
  wire or_tmp_3819;
  wire or_tmp_3836;
  wire and_tmp_240;
  wire and_tmp_242;
  wire and_tmp_244;
  wire and_tmp_246;
  wire or_tmp_3973;
  wire nand_tmp_230;
  wire nand_tmp_231;
  wire nand_tmp_232;
  wire nand_tmp_233;
  wire nand_tmp_234;
  wire nand_tmp_235;
  wire nor_tmp_653;
  wire nor_tmp_656;
  wire nor_tmp_657;
  wire nor_tmp_660;
  wire nor_tmp_661;
  wire nor_tmp_664;
  wire nor_tmp_665;
  wire nor_tmp_668;
  wire and_dcpl_78;
  wire or_dcpl_4;
  wire and_dcpl_96;
  wire and_dcpl_98;
  wire or_dcpl_8;
  wire and_dcpl_105;
  wire and_dcpl_106;
  wire and_dcpl_107;
  wire and_dcpl_109;
  wire and_dcpl_132;
  wire and_dcpl_138;
  wire and_dcpl_141;
  wire and_dcpl_142;
  wire and_dcpl_144;
  wire or_dcpl_44;
  wire and_dcpl_145;
  wire and_dcpl_173;
  wire and_dcpl_176;
  wire and_dcpl_177;
  wire and_dcpl_178;
  wire and_dcpl_180;
  wire and_dcpl_203;
  wire and_dcpl_209;
  wire and_dcpl_212;
  wire and_dcpl_214;
  wire or_dcpl_80;
  wire and_dcpl_215;
  wire and_dcpl_243;
  wire and_dcpl_246;
  wire and_dcpl_247;
  wire and_dcpl_248;
  wire and_dcpl_250;
  wire and_dcpl_273;
  wire and_dcpl_279;
  wire and_dcpl_282;
  wire and_dcpl_284;
  wire or_dcpl_116;
  wire and_dcpl_285;
  wire and_dcpl_313;
  wire and_dcpl_316;
  wire and_dcpl_317;
  wire and_dcpl_318;
  wire and_dcpl_320;
  wire and_dcpl_343;
  wire and_dcpl_349;
  wire and_dcpl_352;
  wire and_dcpl_354;
  wire or_dcpl_152;
  wire and_dcpl_355;
  wire and_dcpl_383;
  wire and_dcpl_390;
  wire and_dcpl_393;
  wire and_dcpl_394;
  wire and_dcpl_398;
  wire and_dcpl_401;
  wire and_dcpl_402;
  wire and_dcpl_406;
  wire and_dcpl_409;
  wire and_dcpl_410;
  wire and_dcpl_412;
  wire and_dcpl_415;
  wire and_dcpl_416;
  wire and_dcpl_419;
  wire and_dcpl_423;
  wire and_dcpl_427;
  wire and_dcpl_428;
  wire and_dcpl_433;
  wire and_dcpl_437;
  wire and_dcpl_453;
  wire and_dcpl_454;
  wire or_dcpl_159;
  wire and_dcpl_458;
  wire and_dcpl_459;
  wire and_dcpl_464;
  wire and_dcpl_465;
  wire and_dcpl_468;
  wire and_dcpl_471;
  wire and_dcpl_488;
  wire or_dcpl_163;
  wire and_dcpl_495;
  wire and_dcpl_496;
  wire and_dcpl_498;
  wire and_dcpl_504;
  wire and_dcpl_524;
  wire and_dcpl_526;
  wire or_dcpl_167;
  wire and_dcpl_530;
  wire and_dcpl_535;
  wire and_dcpl_539;
  wire and_dcpl_559;
  wire and_dcpl_560;
  wire and_dcpl_564;
  wire and_dcpl_565;
  wire and_dcpl_567;
  wire and_dcpl_573;
  wire and_dcpl_575;
  wire and_dcpl_582;
  wire and_dcpl_583;
  wire and_dcpl_584;
  wire and_dcpl_585;
  wire and_dcpl_591;
  wire and_dcpl_593;
  wire and_dcpl_597;
  wire and_dcpl_600;
  wire and_dcpl_601;
  wire and_dcpl_603;
  wire and_dcpl_609;
  wire and_dcpl_611;
  wire and_dcpl_613;
  wire and_dcpl_615;
  wire and_dcpl_627;
  wire and_dcpl_630;
  wire and_dcpl_631;
  wire and_dcpl_633;
  wire or_dcpl_186;
  wire and_dcpl_639;
  wire or_tmp_4220;
  wire and_dcpl_641;
  wire and_dcpl_642;
  wire and_dcpl_645;
  wire and_dcpl_654;
  wire and_dcpl_655;
  wire and_dcpl_662;
  wire and_dcpl_663;
  wire and_dcpl_670;
  wire and_dcpl_671;
  wire mux_tmp_1821;
  wire and_dcpl_678;
  wire and_dcpl_679;
  wire and_dcpl_688;
  wire and_dcpl_690;
  wire and_dcpl_691;
  wire and_dcpl_699;
  wire and_dcpl_701;
  wire and_dcpl_702;
  wire and_dcpl_712;
  wire and_dcpl_713;
  wire nor_tmp_686;
  wire and_dcpl_717;
  wire and_dcpl_719;
  wire and_dcpl_720;
  wire and_dcpl_740;
  wire and_dcpl_741;
  wire and_dcpl_752;
  wire and_dcpl_753;
  wire and_dcpl_764;
  wire and_dcpl_765;
  wire and_dcpl_776;
  wire and_dcpl_777;
  wire and_dcpl_784;
  wire and_dcpl_785;
  wire and_dcpl_787;
  wire and_dcpl_798;
  wire and_dcpl_801;
  wire and_dcpl_807;
  wire and_dcpl_808;
  wire and_dcpl_810;
  wire and_dcpl_821;
  wire and_dcpl_825;
  wire and_dcpl_831;
  wire and_dcpl_832;
  wire and_dcpl_834;
  wire and_dcpl_845;
  wire and_dcpl_847;
  wire and_dcpl_856;
  wire and_dcpl_857;
  wire and_dcpl_859;
  wire and_dcpl_870;
  wire and_dcpl_872;
  wire and_dcpl_874;
  wire or_dcpl_257;
  wire or_dcpl_264;
  wire or_dcpl_267;
  wire or_dcpl_269;
  wire or_dcpl_276;
  wire or_dcpl_278;
  wire and_dcpl_927;
  wire mux_tmp_1835;
  wire or_dcpl_280;
  wire and_dcpl_930;
  wire and_dcpl_935;
  wire and_dcpl_936;
  wire and_dcpl_937;
  wire mux_tmp_1836;
  wire or_dcpl_283;
  wire and_dcpl_940;
  wire and_dcpl_941;
  wire and_dcpl_943;
  wire and_dcpl_944;
  wire and_dcpl_945;
  wire and_dcpl_947;
  wire mux_tmp_1837;
  wire or_dcpl_286;
  wire and_dcpl_949;
  wire and_dcpl_954;
  wire and_dcpl_955;
  wire and_dcpl_958;
  wire mux_tmp_1838;
  wire or_dcpl_289;
  wire and_dcpl_959;
  wire and_dcpl_961;
  wire and_dcpl_962;
  wire or_dcpl_294;
  wire or_dcpl_295;
  wire or_dcpl_336;
  wire or_dcpl_342;
  wire or_dcpl_357;
  wire or_dcpl_409;
  wire and_dcpl_1007;
  wire and_dcpl_1009;
  wire mux_tmp_1845;
  wire and_dcpl_1060;
  wire or_dcpl_499;
  wire or_dcpl_542;
  wire or_dcpl_585;
  wire or_dcpl_628;
  wire or_dcpl_630;
  wire or_dcpl_631;
  wire or_dcpl_634;
  wire or_dcpl_637;
  wire or_dcpl_640;
  wire and_dcpl_1217;
  wire and_dcpl_1219;
  wire and_dcpl_1224;
  wire and_dcpl_1226;
  wire and_dcpl_1230;
  wire and_dcpl_1232;
  wire or_dcpl_660;
  wire and_dcpl_1243;
  wire and_dcpl_1247;
  wire and_dcpl_1252;
  wire and_dcpl_1256;
  wire and_dcpl_1261;
  wire and_dcpl_1265;
  wire and_dcpl_1270;
  wire and_dcpl_1274;
  wire or_dcpl_699;
  wire and_dcpl_1335;
  wire or_dcpl_727;
  wire and_dcpl_1338;
  wire and_dcpl_1348;
  wire or_dcpl_732;
  wire and_dcpl_1351;
  wire and_dcpl_1361;
  wire or_dcpl_737;
  wire and_dcpl_1364;
  wire mux_tmp_1861;
  wire and_dcpl_1373;
  wire and_dcpl_1374;
  wire or_dcpl_742;
  wire and_dcpl_1377;
  wire mux_tmp_1862;
  wire and_dcpl_1404;
  wire and_dcpl_1415;
  wire and_dcpl_1426;
  wire and_dcpl_1437;
  wire and_dcpl_1448;
  wire and_dcpl_1450;
  wire and_dcpl_1452;
  wire and_dcpl_1454;
  wire and_dcpl_1473;
  wire and_dcpl_1481;
  wire and_dcpl_1484;
  wire and_dcpl_1488;
  wire and_dcpl_1497;
  wire and_dcpl_1504;
  wire and_dcpl_1534;
  wire or_dcpl_818;
  wire and_dcpl_1541;
  wire and_dcpl_1545;
  wire and_dcpl_1556;
  wire and_dcpl_1566;
  wire and_dcpl_1577;
  wire or_tmp_4282;
  wire and_dcpl_1588;
  wire and_dcpl_1596;
  wire and_dcpl_1617;
  wire and_dcpl_1619;
  wire and_dcpl_1624;
  wire and_dcpl_1626;
  wire and_dcpl_1632;
  wire and_dcpl_1634;
  wire and_dcpl_1639;
  wire and_dcpl_1641;
  wire or_dcpl_897;
  wire or_dcpl_903;
  wire or_dcpl_906;
  wire or_dcpl_913;
  wire and_dcpl_1722;
  wire and_dcpl_1731;
  wire and_dcpl_1758;
  wire and_dcpl_1759;
  wire and_dcpl_1760;
  wire and_dcpl_1764;
  wire and_dcpl_1772;
  wire and_dcpl_1773;
  wire and_dcpl_1777;
  wire and_dcpl_1785;
  wire and_dcpl_1786;
  wire and_dcpl_1790;
  wire and_dcpl_1798;
  wire and_dcpl_1799;
  wire and_dcpl_1803;
  wire and_dcpl_1852;
  wire and_dcpl_1853;
  wire and_dcpl_1854;
  wire and_dcpl_1856;
  wire and_dcpl_1857;
  wire and_dcpl_1858;
  wire and_dcpl_1859;
  wire and_dcpl_1860;
  wire and_dcpl_1862;
  wire and_dcpl_1863;
  wire or_dcpl_985;
  wire or_dcpl_990;
  wire or_dcpl_995;
  wire or_dcpl_1000;
  wire or_dcpl_1005;
  wire or_dcpl_1010;
  wire and_dcpl_1927;
  wire or_dcpl_1015;
  wire and_dcpl_1947;
  wire and_dcpl_1953;
  wire and_dcpl_1957;
  wire and_dcpl_1961;
  wire and_dcpl_1979;
  wire and_dcpl_1980;
  wire and_dcpl_1984;
  wire and_dcpl_1989;
  wire and_dcpl_1993;
  wire and_dcpl_2005;
  wire and_dcpl_2011;
  wire and_dcpl_2015;
  wire or_tmp_4339;
  wire or_tmp_4457;
  reg inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs;
  reg inp_lookup_1_FpMantRNE_24U_11U_else_and_svs;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_3;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3;
  reg inp_lookup_1_FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs;
  reg [21:0] FpMul_6U_10U_p_mant_p1_1_sva;
  reg IsNaN_6U_10U_1_land_1_lpi_1_dfm;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_3;
  reg inp_lookup_1_FpAdd_6U_10U_is_a_greater_oif_equal_svs;
  reg IsNaN_6U_23U_land_1_lpi_1_dfm;
  reg IsInf_6U_23U_land_1_lpi_1_dfm;
  reg [5:0] IntLeadZero_35U_1_leading_sign_35_0_rtn_1_sva;
  reg inp_lookup_1_FpMantRNE_36U_11U_1_else_and_svs;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_3;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_3;
  reg inp_lookup_1_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs;
  reg [21:0] FpMul_6U_10U_1_p_mant_p1_1_sva;
  reg FpMantRNE_22U_11U_1_else_carry_1_sva_1;
  reg IsNaN_6U_10U_5_land_1_lpi_1_dfm;
  reg inp_lookup_1_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs;
  reg [21:0] FpMul_6U_10U_2_p_mant_p1_1_sva;
  reg IsNaN_6U_10U_7_land_1_lpi_1_dfm;
  reg inp_lookup_1_FpAdd_6U_10U_1_is_a_greater_oif_equal_svs;
  reg IsInf_6U_23U_1_land_1_lpi_1_dfm;
  reg inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs;
  reg inp_lookup_2_FpMantRNE_24U_11U_else_and_svs;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_3;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3;
  reg inp_lookup_2_FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs;
  reg [21:0] FpMul_6U_10U_p_mant_p1_2_sva;
  reg IsNaN_6U_10U_1_land_2_lpi_1_dfm;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_3;
  reg inp_lookup_2_FpAdd_6U_10U_is_a_greater_oif_equal_svs;
  reg IsNaN_6U_23U_land_2_lpi_1_dfm;
  reg IsInf_6U_23U_land_2_lpi_1_dfm;
  reg [5:0] IntLeadZero_35U_1_leading_sign_35_0_rtn_2_sva;
  reg inp_lookup_2_FpMantRNE_36U_11U_1_else_and_svs;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_3;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_3;
  reg inp_lookup_2_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs;
  reg [21:0] FpMul_6U_10U_1_p_mant_p1_2_sva;
  reg FpMantRNE_22U_11U_1_else_carry_2_sva_1;
  reg IsNaN_6U_10U_5_land_2_lpi_1_dfm;
  reg inp_lookup_2_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs;
  reg [21:0] FpMul_6U_10U_2_p_mant_p1_2_sva;
  reg IsNaN_6U_10U_7_land_2_lpi_1_dfm;
  reg inp_lookup_2_FpAdd_6U_10U_1_is_a_greater_oif_equal_svs;
  reg IsInf_6U_23U_1_land_2_lpi_1_dfm;
  reg [22:0] FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2;
  reg inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs;
  reg inp_lookup_3_FpMantRNE_24U_11U_else_and_svs;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_3;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3;
  reg inp_lookup_3_FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs;
  reg [21:0] FpMul_6U_10U_p_mant_p1_3_sva;
  reg IsNaN_6U_10U_1_land_3_lpi_1_dfm;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_3;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_3;
  reg inp_lookup_3_FpAdd_6U_10U_is_a_greater_oif_equal_svs;
  reg IsNaN_6U_23U_land_3_lpi_1_dfm;
  reg IsInf_6U_23U_land_3_lpi_1_dfm;
  reg [5:0] IntLeadZero_35U_1_leading_sign_35_0_rtn_3_sva;
  reg inp_lookup_3_FpMantRNE_36U_11U_1_else_and_svs;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_3_lpi_1_dfm_3;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_3_lpi_1_dfm_3;
  reg inp_lookup_3_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs;
  reg [21:0] FpMul_6U_10U_1_p_mant_p1_3_sva;
  reg FpMantRNE_22U_11U_1_else_carry_3_sva_1;
  reg IsNaN_6U_10U_5_land_3_lpi_1_dfm;
  reg inp_lookup_3_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs;
  reg [21:0] FpMul_6U_10U_2_p_mant_p1_3_sva;
  reg IsNaN_6U_10U_7_land_3_lpi_1_dfm;
  reg inp_lookup_3_FpAdd_6U_10U_1_is_a_greater_oif_equal_svs;
  reg IsInf_6U_23U_1_land_3_lpi_1_dfm;
  reg FpAdd_8U_23U_o_sign_lpi_1_dfm_1;
  reg inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs;
  reg inp_lookup_4_FpMantRNE_24U_11U_else_and_svs;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_3;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_3;
  reg inp_lookup_4_FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs;
  reg [21:0] FpMul_6U_10U_p_mant_p1_sva;
  reg IsNaN_6U_10U_1_land_lpi_1_dfm;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_3;
  reg inp_lookup_4_FpAdd_6U_10U_is_a_greater_oif_equal_svs;
  reg IsNaN_6U_23U_land_lpi_1_dfm;
  reg IsInf_6U_23U_land_lpi_1_dfm;
  reg [5:0] IntLeadZero_35U_1_leading_sign_35_0_rtn_sva;
  reg inp_lookup_4_FpMantRNE_36U_11U_1_else_and_svs;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_3;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_3;
  reg inp_lookup_4_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs;
  reg [21:0] FpMul_6U_10U_1_p_mant_p1_sva;
  reg FpMantRNE_22U_11U_1_else_carry_sva;
  reg IsNaN_6U_10U_5_land_lpi_1_dfm;
  reg inp_lookup_4_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs;
  reg [21:0] FpMul_6U_10U_2_p_mant_p1_sva;
  reg IsNaN_6U_10U_7_land_lpi_1_dfm;
  reg inp_lookup_4_FpAdd_6U_10U_1_is_a_greater_oif_equal_svs;
  reg IsInf_6U_23U_1_land_lpi_1_dfm;
  reg main_stage_v_1;
  reg main_stage_v_2;
  reg main_stage_v_3;
  reg main_stage_v_4;
  reg main_stage_v_5;
  reg main_stage_v_6;
  reg main_stage_v_7;
  reg main_stage_v_8;
  reg main_stage_v_9;
  reg main_stage_v_10;
  reg main_stage_v_11;
  reg main_stage_v_12;
  reg FpAdd_6U_10U_1_is_a_greater_lor_lpi_1_dfm_5;
  reg FpMul_6U_10U_2_o_sign_lpi_1_dfm_6;
  reg FpMul_6U_10U_2_o_sign_lpi_1_dfm_7;
  reg FpMul_6U_10U_2_o_sign_lpi_1_dfm_8;
  reg FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_5;
  reg FpMul_6U_10U_o_sign_lpi_1_dfm_5;
  reg FpAdd_6U_10U_1_is_a_greater_lor_3_lpi_1_dfm_5;
  reg FpMul_6U_10U_2_o_sign_3_lpi_1_dfm_6;
  reg FpMul_6U_10U_2_o_sign_3_lpi_1_dfm_7;
  reg FpMul_6U_10U_2_o_sign_3_lpi_1_dfm_8;
  reg FpAdd_6U_10U_is_a_greater_lor_3_lpi_1_dfm_5;
  reg FpMul_6U_10U_o_sign_3_lpi_1_dfm_5;
  reg FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_5;
  reg FpMul_6U_10U_2_o_sign_2_lpi_1_dfm_6;
  reg FpMul_6U_10U_2_o_sign_2_lpi_1_dfm_7;
  reg FpMul_6U_10U_2_o_sign_2_lpi_1_dfm_8;
  reg FpAdd_6U_10U_is_a_greater_lor_2_lpi_1_dfm_5;
  reg FpMul_6U_10U_o_sign_2_lpi_1_dfm_5;
  reg FpAdd_6U_10U_1_is_a_greater_lor_1_lpi_1_dfm_5;
  reg FpMul_6U_10U_2_o_sign_1_lpi_1_dfm_6;
  reg FpMul_6U_10U_2_o_sign_1_lpi_1_dfm_7;
  reg FpMul_6U_10U_2_o_sign_1_lpi_1_dfm_8;
  reg FpAdd_6U_10U_is_a_greater_lor_1_lpi_1_dfm_5;
  reg FpMul_6U_10U_o_sign_1_lpi_1_dfm_5;
  reg IsNaN_6U_23U_3_land_lpi_1_dfm_7;
  reg IsNaN_6U_23U_3_land_lpi_1_dfm_8;
  reg IsNaN_6U_23U_3_land_lpi_1_dfm_9;
  reg IsNaN_6U_23U_3_land_lpi_1_dfm_10;
  reg [9:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_lpi_1_dfm_9;
  reg [9:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_lpi_1_dfm_10;
  reg [9:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_lpi_1_dfm_11;
  reg [9:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_lpi_1_dfm_12;
  reg IsNaN_6U_10U_8_land_lpi_1_dfm_4;
  reg FpMul_6U_10U_1_o_sign_lpi_1_dfm_6;
  reg FpMul_6U_10U_1_o_sign_lpi_1_dfm_7;
  reg FpMul_6U_10U_1_o_sign_lpi_1_dfm_8;
  reg IsNaN_6U_10U_2_land_lpi_1_dfm_15;
  reg IsNaN_6U_10U_2_land_lpi_1_dfm_16;
  reg IsNaN_6U_10U_2_land_lpi_1_dfm_17;
  reg IsNaN_6U_10U_2_land_lpi_1_dfm_18;
  reg IsNaN_6U_10U_2_land_lpi_1_dfm_19;
  reg IsNaN_6U_10U_2_land_lpi_1_dfm_20;
  reg IsNaN_6U_10U_2_land_lpi_1_dfm_21;
  reg IsNaN_6U_10U_2_land_lpi_1_dfm_22;
  reg IsNaN_6U_10U_2_land_lpi_1_dfm_23;
  reg IsNaN_6U_10U_2_land_lpi_1_dfm_24;
  reg IsNaN_6U_10U_2_land_lpi_1_dfm_25;
  reg IsNaN_6U_10U_2_land_lpi_1_dfm_26;
  reg IsNaN_6U_10U_9_land_lpi_1_dfm_6;
  reg IsNaN_6U_10U_9_land_lpi_1_dfm_7;
  reg IsNaN_6U_10U_9_land_lpi_1_dfm_8;
  reg IsNaN_6U_10U_3_land_lpi_1_dfm_6;
  reg IsNaN_6U_10U_3_land_lpi_1_dfm_7;
  reg IsNaN_6U_10U_3_land_lpi_1_dfm_8;
  reg IsNaN_8U_23U_3_land_lpi_1_dfm_5;
  reg IsNaN_8U_23U_3_land_lpi_1_dfm_6;
  reg IsNaN_8U_23U_1_land_lpi_1_dfm_4;
  reg IsNaN_6U_23U_3_land_3_lpi_1_dfm_7;
  reg IsNaN_6U_23U_3_land_3_lpi_1_dfm_8;
  reg IsNaN_6U_23U_3_land_3_lpi_1_dfm_9;
  reg IsNaN_6U_23U_3_land_3_lpi_1_dfm_10;
  reg [9:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_3_lpi_1_dfm_9;
  reg [9:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_3_lpi_1_dfm_10;
  reg [9:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_3_lpi_1_dfm_11;
  reg [9:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_3_lpi_1_dfm_12;
  reg IsNaN_6U_10U_8_land_3_lpi_1_dfm_4;
  reg FpMul_6U_10U_1_o_sign_3_lpi_1_dfm_6;
  reg FpMul_6U_10U_1_o_sign_3_lpi_1_dfm_7;
  reg FpMul_6U_10U_1_o_sign_3_lpi_1_dfm_8;
  reg IsNaN_6U_10U_2_land_3_lpi_1_dfm_15;
  reg IsNaN_6U_10U_2_land_3_lpi_1_dfm_16;
  reg IsNaN_6U_10U_2_land_3_lpi_1_dfm_17;
  reg IsNaN_6U_10U_2_land_3_lpi_1_dfm_18;
  reg IsNaN_6U_10U_2_land_3_lpi_1_dfm_19;
  reg IsNaN_6U_10U_2_land_3_lpi_1_dfm_20;
  reg IsNaN_6U_10U_2_land_3_lpi_1_dfm_21;
  reg IsNaN_6U_10U_2_land_3_lpi_1_dfm_22;
  reg IsNaN_6U_10U_2_land_3_lpi_1_dfm_23;
  reg IsNaN_6U_10U_2_land_3_lpi_1_dfm_24;
  reg IsNaN_6U_10U_2_land_3_lpi_1_dfm_25;
  reg IsNaN_6U_10U_2_land_3_lpi_1_dfm_26;
  reg IsNaN_6U_10U_9_land_3_lpi_1_dfm_6;
  reg IsNaN_6U_10U_9_land_3_lpi_1_dfm_7;
  reg IsNaN_6U_10U_9_land_3_lpi_1_dfm_8;
  reg IsNaN_6U_10U_3_land_3_lpi_1_dfm_6;
  reg IsNaN_6U_10U_3_land_3_lpi_1_dfm_7;
  reg IsNaN_6U_10U_3_land_3_lpi_1_dfm_8;
  reg IsNaN_8U_23U_3_land_3_lpi_1_dfm_6;
  reg IsNaN_8U_23U_3_land_3_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_3_lpi_1_dfm_4;
  reg IsNaN_6U_23U_3_land_2_lpi_1_dfm_7;
  reg IsNaN_6U_23U_3_land_2_lpi_1_dfm_8;
  reg IsNaN_6U_23U_3_land_2_lpi_1_dfm_9;
  reg IsNaN_6U_23U_3_land_2_lpi_1_dfm_10;
  reg [9:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_2_lpi_1_dfm_9;
  reg [9:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_2_lpi_1_dfm_10;
  reg [9:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_2_lpi_1_dfm_11;
  reg [9:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_2_lpi_1_dfm_12;
  reg IsNaN_6U_10U_8_land_2_lpi_1_dfm_4;
  reg FpMul_6U_10U_1_o_sign_2_lpi_1_dfm_6;
  reg FpMul_6U_10U_1_o_sign_2_lpi_1_dfm_7;
  reg FpMul_6U_10U_1_o_sign_2_lpi_1_dfm_8;
  reg IsNaN_6U_10U_2_land_2_lpi_1_dfm_15;
  reg IsNaN_6U_10U_2_land_2_lpi_1_dfm_16;
  reg IsNaN_6U_10U_2_land_2_lpi_1_dfm_17;
  reg IsNaN_6U_10U_2_land_2_lpi_1_dfm_18;
  reg IsNaN_6U_10U_2_land_2_lpi_1_dfm_19;
  reg IsNaN_6U_10U_2_land_2_lpi_1_dfm_20;
  reg IsNaN_6U_10U_2_land_2_lpi_1_dfm_21;
  reg IsNaN_6U_10U_2_land_2_lpi_1_dfm_22;
  reg IsNaN_6U_10U_2_land_2_lpi_1_dfm_23;
  reg IsNaN_6U_10U_2_land_2_lpi_1_dfm_24;
  reg IsNaN_6U_10U_2_land_2_lpi_1_dfm_25;
  reg IsNaN_6U_10U_2_land_2_lpi_1_dfm_26;
  reg IsNaN_6U_10U_9_land_2_lpi_1_dfm_6;
  reg IsNaN_6U_10U_9_land_2_lpi_1_dfm_7;
  reg IsNaN_6U_10U_9_land_2_lpi_1_dfm_8;
  reg IsNaN_6U_10U_3_land_2_lpi_1_dfm_6;
  reg IsNaN_6U_10U_3_land_2_lpi_1_dfm_7;
  reg IsNaN_6U_10U_3_land_2_lpi_1_dfm_8;
  reg IsNaN_8U_23U_3_land_2_lpi_1_dfm_6;
  reg IsNaN_8U_23U_3_land_2_lpi_1_dfm_7;
  reg IsNaN_8U_23U_1_land_2_lpi_1_dfm_4;
  reg IsNaN_6U_23U_3_land_1_lpi_1_dfm_7;
  reg IsNaN_6U_23U_3_land_1_lpi_1_dfm_8;
  reg IsNaN_6U_23U_3_land_1_lpi_1_dfm_9;
  reg IsNaN_6U_23U_3_land_1_lpi_1_dfm_10;
  reg [9:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_1_lpi_1_dfm_9;
  reg [9:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_1_lpi_1_dfm_10;
  reg [9:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_1_lpi_1_dfm_11;
  reg [9:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_1_lpi_1_dfm_12;
  reg IsNaN_6U_10U_8_land_1_lpi_1_dfm_6;
  reg IsNaN_6U_10U_8_land_1_lpi_1_dfm_7;
  reg FpMul_6U_10U_1_o_sign_1_lpi_1_dfm_6;
  reg FpMul_6U_10U_1_o_sign_1_lpi_1_dfm_7;
  reg FpMul_6U_10U_1_o_sign_1_lpi_1_dfm_8;
  reg IsNaN_6U_10U_2_land_1_lpi_1_dfm_15;
  reg IsNaN_6U_10U_2_land_1_lpi_1_dfm_16;
  reg IsNaN_6U_10U_2_land_1_lpi_1_dfm_17;
  reg IsNaN_6U_10U_2_land_1_lpi_1_dfm_18;
  reg IsNaN_6U_10U_2_land_1_lpi_1_dfm_19;
  reg IsNaN_6U_10U_2_land_1_lpi_1_dfm_20;
  reg IsNaN_6U_10U_2_land_1_lpi_1_dfm_21;
  reg IsNaN_6U_10U_2_land_1_lpi_1_dfm_22;
  reg IsNaN_6U_10U_2_land_1_lpi_1_dfm_23;
  reg IsNaN_6U_10U_2_land_1_lpi_1_dfm_24;
  reg IsNaN_6U_10U_2_land_1_lpi_1_dfm_25;
  reg IsNaN_6U_10U_2_land_1_lpi_1_dfm_26;
  reg IsNaN_6U_10U_9_land_1_lpi_1_dfm_6;
  reg IsNaN_6U_10U_9_land_1_lpi_1_dfm_7;
  reg IsNaN_6U_10U_9_land_1_lpi_1_dfm_8;
  reg IsNaN_6U_10U_3_land_1_lpi_1_dfm_6;
  reg IsNaN_6U_10U_3_land_1_lpi_1_dfm_7;
  reg IsNaN_6U_10U_3_land_1_lpi_1_dfm_8;
  reg IsNaN_8U_23U_3_land_1_lpi_1_dfm_6;
  reg IsNaN_8U_23U_3_land_1_lpi_1_dfm_7;
  reg inp_lookup_if_unequal_tmp_12;
  reg inp_lookup_else_unequal_tmp_32;
  reg inp_lookup_else_unequal_tmp_33;
  reg inp_lookup_else_unequal_tmp_35;
  reg inp_lookup_else_unequal_tmp_36;
  reg inp_lookup_else_unequal_tmp_37;
  reg inp_lookup_else_unequal_tmp_38;
  reg inp_lookup_if_unequal_tmp_19;
  reg inp_lookup_else_unequal_tmp_55;
  reg [17:0] IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_7;
  wire [18:0] nl_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_7;
  reg [17:0] IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_8;
  reg [17:0] IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_9;
  reg [17:0] IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_10;
  reg [17:0] IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_11;
  reg [17:0] IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_12;
  reg [2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_lpi_1_dfm_9;
  reg [2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_lpi_1_dfm_10;
  reg [2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_lpi_1_dfm_11;
  reg [2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_lpi_1_dfm_12;
  reg [9:0] FpFractionToFloat_35U_6U_10U_1_o_mant_lpi_1_dfm_6;
  reg FpFractionToFloat_35U_6U_10U_1_if_else_else_if_slc_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_5_mdf_sva_2;
  reg [31:0] IntSaturation_51U_32U_o_lpi_1_dfm_11;
  reg [31:0] IntSaturation_51U_32U_o_lpi_1_dfm_12;
  reg [31:0] IntSaturation_51U_32U_o_lpi_1_dfm_13;
  reg [31:0] IntSaturation_51U_32U_o_lpi_1_dfm_14;
  reg [31:0] IntSaturation_51U_32U_o_lpi_1_dfm_15;
  reg [31:0] IntSaturation_51U_32U_o_lpi_1_dfm_16;
  reg [31:0] IntSaturation_51U_32U_o_lpi_1_dfm_17;
  reg FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_sva_2;
  reg [49:0] FpAdd_8U_23U_1_int_mant_p1_sva_3;
  reg [7:0] FpAdd_8U_23U_o_expo_lpi_1_dfm_10;
  reg [48:0] FpAdd_8U_23U_int_mant_1_sva_5;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_sva_2;
  reg [17:0] IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_7;
  wire [18:0] nl_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_7;
  reg [17:0] IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_8;
  reg [17:0] IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_9;
  reg [17:0] IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_10;
  reg [17:0] IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_11;
  reg [17:0] IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_12;
  reg [2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_3_lpi_1_dfm_9;
  reg [2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_3_lpi_1_dfm_10;
  reg [2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_3_lpi_1_dfm_11;
  reg [2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_3_lpi_1_dfm_12;
  reg [9:0] FpFractionToFloat_35U_6U_10U_1_o_mant_3_lpi_1_dfm_6;
  reg FpFractionToFloat_35U_6U_10U_1_if_else_else_if_slc_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_5_mdf_3_sva_2;
  reg [31:0] IntSaturation_51U_32U_o_3_lpi_1_dfm_11;
  reg [31:0] IntSaturation_51U_32U_o_3_lpi_1_dfm_12;
  reg [31:0] IntSaturation_51U_32U_o_3_lpi_1_dfm_13;
  reg [31:0] IntSaturation_51U_32U_o_3_lpi_1_dfm_14;
  reg [31:0] IntSaturation_51U_32U_o_3_lpi_1_dfm_15;
  reg [31:0] IntSaturation_51U_32U_o_3_lpi_1_dfm_16;
  reg [31:0] IntSaturation_51U_32U_o_3_lpi_1_dfm_17;
  reg FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_3_sva_2;
  reg [49:0] FpAdd_8U_23U_1_int_mant_p1_3_sva_3;
  reg [7:0] FpAdd_8U_23U_o_expo_3_lpi_1_dfm_10;
  reg [48:0] FpAdd_8U_23U_int_mant_4_sva_5;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_2;
  reg [17:0] IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_7;
  wire [18:0] nl_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_7;
  reg [17:0] IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_8;
  reg [17:0] IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_9;
  reg [17:0] IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_10;
  reg [17:0] IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_11;
  reg [17:0] IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_12;
  reg [2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_2_lpi_1_dfm_9;
  reg [2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_2_lpi_1_dfm_10;
  reg [2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_2_lpi_1_dfm_11;
  reg [2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_2_lpi_1_dfm_12;
  reg [9:0] FpFractionToFloat_35U_6U_10U_1_o_mant_2_lpi_1_dfm_6;
  reg FpFractionToFloat_35U_6U_10U_1_if_else_else_if_slc_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_5_mdf_2_sva_2;
  reg [31:0] IntSaturation_51U_32U_o_2_lpi_1_dfm_11;
  reg [31:0] IntSaturation_51U_32U_o_2_lpi_1_dfm_12;
  reg [31:0] IntSaturation_51U_32U_o_2_lpi_1_dfm_13;
  reg [31:0] IntSaturation_51U_32U_o_2_lpi_1_dfm_14;
  reg [31:0] IntSaturation_51U_32U_o_2_lpi_1_dfm_15;
  reg [31:0] IntSaturation_51U_32U_o_2_lpi_1_dfm_16;
  reg [31:0] IntSaturation_51U_32U_o_2_lpi_1_dfm_17;
  reg FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_2_sva_2;
  reg [49:0] FpAdd_8U_23U_1_int_mant_p1_2_sva_3;
  reg [7:0] FpAdd_8U_23U_o_expo_2_lpi_1_dfm_10;
  reg [48:0] FpAdd_8U_23U_int_mant_3_sva_5;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_2;
  reg [17:0] IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_7;
  wire [18:0] nl_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_7;
  reg [17:0] IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_8;
  reg [17:0] IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_9;
  reg [17:0] IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_10;
  reg [17:0] IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_11;
  reg [17:0] IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_12;
  reg [2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_1_lpi_1_dfm_9;
  reg [2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_1_lpi_1_dfm_10;
  reg [2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_1_lpi_1_dfm_11;
  reg [2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_1_lpi_1_dfm_12;
  reg [9:0] FpFractionToFloat_35U_6U_10U_1_o_mant_1_lpi_1_dfm_6;
  reg FpFractionToFloat_35U_6U_10U_1_if_else_else_if_slc_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_5_mdf_1_sva_2;
  reg [31:0] IntSaturation_51U_32U_o_1_lpi_1_dfm_11;
  reg [31:0] IntSaturation_51U_32U_o_1_lpi_1_dfm_12;
  reg [31:0] IntSaturation_51U_32U_o_1_lpi_1_dfm_13;
  reg [31:0] IntSaturation_51U_32U_o_1_lpi_1_dfm_14;
  reg [31:0] IntSaturation_51U_32U_o_1_lpi_1_dfm_15;
  reg [31:0] IntSaturation_51U_32U_o_1_lpi_1_dfm_16;
  reg [31:0] IntSaturation_51U_32U_o_1_lpi_1_dfm_17;
  reg FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_1_sva_2;
  reg inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_2;
  reg [49:0] FpAdd_8U_23U_1_int_mant_p1_1_sva_3;
  reg [7:0] FpAdd_8U_23U_o_expo_1_lpi_1_dfm_10;
  reg [48:0] FpAdd_8U_23U_int_mant_2_sva_5;
  reg FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_2;
  reg [1:0] cfg_precision_1_sva_16;
  reg [1:0] cfg_precision_1_sva_17;
  reg [1:0] cfg_precision_1_sva_18;
  reg [1:0] cfg_precision_1_sva_19;
  reg [1:0] cfg_precision_1_sva_20;
  reg FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_5;
  reg [48:0] FpAdd_8U_23U_addend_larger_qr_1_lpi_1_dfm_4;
  reg [48:0] FpAdd_8U_23U_addend_smaller_qr_1_lpi_1_dfm_4;
  reg inp_lookup_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3;
  reg inp_lookup_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_4;
  reg FpAdd_8U_23U_o_sign_1_lpi_1_dfm_7;
  reg FpAdd_8U_23U_o_sign_1_lpi_1_dfm_5;
  reg FpAdd_8U_23U_o_sign_1_lpi_1_dfm_8;
  reg [22:0] FpAdd_8U_23U_o_mant_1_lpi_1_dfm_6;
  reg FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5;
  reg inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4;
  reg inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5;
  reg [7:0] FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_12;
  reg inp_lookup_1_FpMantRNE_49U_24U_1_else_and_svs_2;
  reg IsNaN_8U_23U_2_land_1_lpi_1_dfm_9;
  reg FpAdd_8U_23U_1_o_sign_1_lpi_1_dfm_5;
  reg [22:0] FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_6;
  reg inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2;
  reg inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2;
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_1_sva_2;
  wire [5:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_1_sva_2;
  reg inp_lookup_1_FpMantRNE_24U_11U_else_and_svs_2;
  reg [9:0] FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_1_lpi_1_dfm_9;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_15;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_16;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_17;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_18;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_19;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_20;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_21;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_22;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_23;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_15;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_16;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_17;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_18;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_19;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_20;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_21;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_22;
  reg FpMul_6U_10U_lor_6_lpi_1_dfm_4;
  reg [21:0] FpMul_6U_10U_p_mant_p1_1_sva_2;
  reg [5:0] FpMul_6U_10U_else_2_else_ac_int_cctor_1_sva_2;
  wire [6:0] nl_FpMul_6U_10U_else_2_else_ac_int_cctor_1_sva_2;
  reg IsNaN_6U_10U_land_1_lpi_1_dfm_5;
  reg IsNaN_6U_10U_land_1_lpi_1_dfm_6;
  reg IsNaN_6U_10U_1_land_1_lpi_1_dfm_5;
  reg IsNaN_6U_10U_1_land_1_lpi_1_dfm_6;
  reg [9:0] FpMul_6U_10U_o_mant_1_lpi_1_dfm_7;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_18;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_19;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_20;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_21;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_22;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_23;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_24;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_25;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_26;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_18;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_19;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_20;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_21;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_22;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_23;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_24;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_25;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_26;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_27;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_28;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_29;
  reg [22:0] FpAdd_6U_10U_a_int_mant_p1_1_sva_2;
  reg [22:0] FpAdd_6U_10U_b_int_mant_p1_1_sva_2;
  reg inp_lookup_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_4;
  reg inp_lookup_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_5;
  reg [23:0] FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_4;
  reg [4:0] IntLeadZero_23U_leading_sign_23_0_rtn_1_sva_2;
  reg [5:0] IntLeadZero_35U_leading_sign_35_0_rtn_1_sva_2;
  reg FpFractionToFloat_35U_6U_10U_is_zero_1_lpi_1_dfm_5;
  reg [9:0] inp_lookup_else_if_a0_9_0_1_lpi_1_dfm_10;
  reg [5:0] IntLeadZero_35U_1_leading_sign_35_0_rtn_1_sva_2;
  reg inp_lookup_1_FpMantRNE_36U_11U_1_else_and_svs_2;
  reg [9:0] FpFractionToFloat_35U_6U_10U_1_o_mant_1_lpi_1_dfm_8;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_8;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_11;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_8;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_11;
  reg FpMul_6U_10U_1_lor_6_lpi_1_dfm_5;
  reg FpMul_6U_10U_1_lor_6_lpi_1_dfm_6;
  reg IsNaN_6U_10U_5_land_1_lpi_1_dfm_5;
  reg IsNaN_6U_10U_5_land_1_lpi_1_dfm_6;
  reg [9:0] FpMul_6U_10U_1_o_mant_1_lpi_1_dfm_10;
  reg [9:0] FpMul_6U_10U_1_o_mant_1_lpi_1_dfm_11;
  reg FpMul_6U_10U_2_lor_6_lpi_1_dfm_5;
  reg FpMul_6U_10U_2_lor_6_lpi_1_dfm_6;
  reg IsNaN_6U_10U_6_land_1_lpi_1_dfm_5;
  reg IsNaN_6U_10U_7_land_1_lpi_1_dfm_5;
  reg IsNaN_6U_10U_7_land_1_lpi_1_dfm_6;
  reg [9:0] FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_8;
  reg [5:0] FpAdd_6U_10U_1_qr_2_lpi_1_dfm_5;
  reg [22:0] FpAdd_6U_10U_1_b_int_mant_p1_1_sva_2;
  reg inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4;
  reg inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5;
  reg [23:0] FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_4;
  reg FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_5;
  reg [48:0] FpAdd_8U_23U_addend_larger_qr_2_lpi_1_dfm_4;
  reg [48:0] FpAdd_8U_23U_addend_smaller_qr_2_lpi_1_dfm_4;
  reg inp_lookup_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3;
  reg inp_lookup_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_4;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_4;
  reg FpAdd_8U_23U_o_sign_2_lpi_1_dfm_7;
  reg FpAdd_8U_23U_o_sign_2_lpi_1_dfm_5;
  reg FpAdd_8U_23U_o_sign_2_lpi_1_dfm_8;
  reg [22:0] FpAdd_8U_23U_o_mant_2_lpi_1_dfm_6;
  reg FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5;
  reg inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4;
  reg inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5;
  reg [7:0] FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_13;
  reg inp_lookup_2_FpMantRNE_49U_24U_1_else_and_svs_2;
  reg IsNaN_8U_23U_2_land_2_lpi_1_dfm_9;
  reg FpAdd_8U_23U_1_o_sign_2_lpi_1_dfm_5;
  reg [22:0] FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_6;
  reg inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2;
  reg inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2;
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_2_sva_2;
  wire [5:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_2_sva_2;
  reg inp_lookup_2_FpMantRNE_24U_11U_else_and_svs_2;
  reg [9:0] FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_2_lpi_1_dfm_9;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_15;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_16;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_17;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_18;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_19;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_20;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_21;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_22;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_23;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_15;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_16;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_17;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_18;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_19;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_20;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_21;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_22;
  reg FpMul_6U_10U_lor_7_lpi_1_dfm_4;
  reg [21:0] FpMul_6U_10U_p_mant_p1_2_sva_2;
  reg [5:0] FpMul_6U_10U_else_2_else_ac_int_cctor_2_sva_2;
  wire [6:0] nl_FpMul_6U_10U_else_2_else_ac_int_cctor_2_sva_2;
  reg IsNaN_6U_10U_land_2_lpi_1_dfm_5;
  reg IsNaN_6U_10U_land_2_lpi_1_dfm_6;
  reg IsNaN_6U_10U_1_land_2_lpi_1_dfm_5;
  reg IsNaN_6U_10U_1_land_2_lpi_1_dfm_6;
  reg [9:0] FpMul_6U_10U_o_mant_2_lpi_1_dfm_7;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_18;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_19;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_20;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_21;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_22;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_23;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_24;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_25;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_26;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_18;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_19;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_20;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_21;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_22;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_23;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_24;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_25;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_26;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_27;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_28;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_29;
  reg [22:0] FpAdd_6U_10U_a_int_mant_p1_2_sva_2;
  reg [22:0] FpAdd_6U_10U_b_int_mant_p1_2_sva_2;
  reg inp_lookup_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_4;
  reg inp_lookup_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_5;
  reg [23:0] FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_4;
  reg [4:0] IntLeadZero_23U_leading_sign_23_0_rtn_2_sva_2;
  reg [5:0] IntLeadZero_35U_leading_sign_35_0_rtn_2_sva_2;
  reg FpFractionToFloat_35U_6U_10U_is_zero_2_lpi_1_dfm_5;
  reg [9:0] inp_lookup_else_if_a0_9_0_2_lpi_1_dfm_10;
  reg [5:0] IntLeadZero_35U_1_leading_sign_35_0_rtn_2_sva_2;
  reg inp_lookup_2_FpMantRNE_36U_11U_1_else_and_svs_2;
  reg [9:0] FpFractionToFloat_35U_6U_10U_1_o_mant_2_lpi_1_dfm_8;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_8;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_11;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_8;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_11;
  reg FpMul_6U_10U_1_lor_7_lpi_1_dfm_5;
  reg FpMul_6U_10U_1_lor_7_lpi_1_dfm_6;
  reg IsNaN_6U_10U_5_land_2_lpi_1_dfm_5;
  reg IsNaN_6U_10U_5_land_2_lpi_1_dfm_6;
  reg [9:0] FpMul_6U_10U_1_o_mant_2_lpi_1_dfm_10;
  reg [9:0] FpMul_6U_10U_1_o_mant_2_lpi_1_dfm_11;
  reg FpMul_6U_10U_2_lor_7_lpi_1_dfm_5;
  reg FpMul_6U_10U_2_lor_7_lpi_1_dfm_6;
  reg [5:0] FpMul_6U_10U_2_else_2_else_ac_int_cctor_2_sva_2;
  reg IsNaN_6U_10U_6_land_2_lpi_1_dfm_5;
  reg IsNaN_6U_10U_7_land_2_lpi_1_dfm_5;
  reg IsNaN_6U_10U_7_land_2_lpi_1_dfm_6;
  reg [9:0] FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_8;
  reg [5:0] FpAdd_6U_10U_1_qr_3_lpi_1_dfm_5;
  reg [22:0] FpAdd_6U_10U_1_b_int_mant_p1_2_sva_2;
  reg inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4;
  reg inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5;
  reg [23:0] FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_4;
  reg FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_5;
  reg [48:0] FpAdd_8U_23U_addend_larger_qr_3_lpi_1_dfm_4;
  reg [48:0] FpAdd_8U_23U_addend_smaller_qr_3_lpi_1_dfm_4;
  reg inp_lookup_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3;
  reg inp_lookup_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_4;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_4;
  reg FpAdd_8U_23U_o_sign_3_lpi_1_dfm_7;
  reg FpAdd_8U_23U_o_sign_3_lpi_1_dfm_8;
  reg FpAdd_8U_23U_o_sign_3_lpi_1_dfm_9;
  reg [22:0] FpAdd_8U_23U_o_mant_3_lpi_1_dfm_6;
  reg FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5;
  reg inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4;
  reg inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5;
  reg IsNaN_8U_23U_2_land_3_lpi_1_dfm_9;
  reg FpAdd_8U_23U_1_o_sign_3_lpi_1_dfm_5;
  reg [22:0] FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_6;
  reg inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2;
  reg inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2;
  reg inp_lookup_3_FpMantRNE_24U_11U_else_and_svs_2;
  reg [9:0] FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_3_lpi_1_dfm_9;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_15;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_16;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_17;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_18;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_19;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_20;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_21;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_22;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_15;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_16;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_17;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_18;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_19;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_20;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_21;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_22;
  reg FpMul_6U_10U_lor_8_lpi_1_dfm_4;
  reg [21:0] FpMul_6U_10U_p_mant_p1_3_sva_2;
  reg [5:0] FpMul_6U_10U_else_2_else_ac_int_cctor_3_sva_2;
  wire [6:0] nl_FpMul_6U_10U_else_2_else_ac_int_cctor_3_sva_2;
  reg IsNaN_6U_10U_land_3_lpi_1_dfm_5;
  reg IsNaN_6U_10U_land_3_lpi_1_dfm_6;
  reg IsNaN_6U_10U_1_land_3_lpi_1_dfm_5;
  reg IsNaN_6U_10U_1_land_3_lpi_1_dfm_6;
  reg [9:0] FpMul_6U_10U_o_mant_3_lpi_1_dfm_7;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_18;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_19;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_20;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_21;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_22;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_23;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_24;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_25;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_26;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_27;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_28;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_29;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_18;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_19;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_20;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_21;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_22;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_23;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_24;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_25;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_26;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_27;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_28;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_29;
  reg [22:0] FpAdd_6U_10U_a_int_mant_p1_3_sva_2;
  reg [22:0] FpAdd_6U_10U_b_int_mant_p1_3_sva_2;
  reg inp_lookup_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_4;
  reg inp_lookup_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_5;
  reg [23:0] FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_4;
  reg [4:0] IntLeadZero_23U_leading_sign_23_0_rtn_3_sva_2;
  reg FpNormalize_6U_23U_lor_3_lpi_1_dfm_5;
  reg [5:0] IntLeadZero_35U_leading_sign_35_0_rtn_3_sva_2;
  reg FpFractionToFloat_35U_6U_10U_is_zero_3_lpi_1_dfm_5;
  reg [9:0] inp_lookup_else_if_a0_9_0_3_lpi_1_dfm_10;
  reg [5:0] IntLeadZero_35U_1_leading_sign_35_0_rtn_3_sva_2;
  reg inp_lookup_3_FpMantRNE_36U_11U_1_else_and_svs_2;
  reg [9:0] FpFractionToFloat_35U_6U_10U_1_o_mant_3_lpi_1_dfm_8;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_8;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_10;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_11;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_8;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_11;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_3_lpi_1_dfm_8;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_3_lpi_1_dfm_9;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_3_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_3_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_3_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_3_lpi_1_dfm_11;
  reg FpMul_6U_10U_1_lor_8_lpi_1_dfm_5;
  reg FpMul_6U_10U_1_lor_8_lpi_1_dfm_6;
  reg IsNaN_6U_10U_5_land_3_lpi_1_dfm_5;
  reg IsNaN_6U_10U_5_land_3_lpi_1_dfm_6;
  reg FpMul_6U_10U_2_lor_8_lpi_1_dfm_5;
  reg FpMul_6U_10U_2_lor_8_lpi_1_dfm_6;
  reg [5:0] FpMul_6U_10U_2_else_2_else_ac_int_cctor_3_sva_2;
  reg IsNaN_6U_10U_6_land_3_lpi_1_dfm_5;
  reg IsNaN_6U_10U_7_land_3_lpi_1_dfm_5;
  reg IsNaN_6U_10U_7_land_3_lpi_1_dfm_6;
  reg [9:0] FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_8;
  reg [5:0] FpAdd_6U_10U_1_qr_4_lpi_1_dfm_5;
  reg [22:0] FpAdd_6U_10U_1_b_int_mant_p1_3_sva_2;
  reg inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4;
  reg inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5;
  reg [23:0] FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_4;
  reg [48:0] FpAdd_8U_23U_addend_larger_qr_lpi_1_dfm_4;
  reg [48:0] FpAdd_8U_23U_addend_smaller_qr_lpi_1_dfm_4;
  reg inp_lookup_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3;
  reg inp_lookup_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_4;
  reg IsNaN_8U_23U_land_lpi_1_dfm_4;
  reg FpAdd_8U_23U_o_sign_lpi_1_dfm_7;
  reg FpAdd_8U_23U_o_sign_lpi_1_dfm_8;
  reg FpAdd_8U_23U_o_sign_lpi_1_dfm_9;
  reg [22:0] FpAdd_8U_23U_o_mant_lpi_1_dfm_6;
  reg FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5;
  reg inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4;
  reg [7:0] FpAdd_8U_23U_1_o_expo_lpi_1_dfm_13;
  reg inp_lookup_4_FpMantRNE_49U_24U_1_else_and_svs_2;
  reg IsNaN_8U_23U_2_land_lpi_1_dfm_9;
  reg FpAdd_8U_23U_1_o_sign_lpi_1_dfm_5;
  reg [22:0] FpAdd_8U_23U_1_o_mant_lpi_1_dfm_6;
  reg inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2;
  reg inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2;
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva_2;
  wire [5:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva_2;
  reg inp_lookup_4_FpMantRNE_24U_11U_else_and_svs_2;
  reg [9:0] FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_lpi_1_dfm_9;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_15;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_16;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_17;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_18;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_19;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_20;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_21;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_22;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_23;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_15;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_16;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_17;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_18;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_19;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_20;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_21;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_22;
  reg FpMul_6U_10U_lor_1_lpi_1_dfm_4;
  reg [21:0] FpMul_6U_10U_p_mant_p1_sva_2;
  reg [5:0] FpMul_6U_10U_else_2_else_ac_int_cctor_sva_2;
  wire [6:0] nl_FpMul_6U_10U_else_2_else_ac_int_cctor_sva_2;
  reg IsNaN_6U_10U_land_lpi_1_dfm_5;
  reg IsNaN_6U_10U_land_lpi_1_dfm_6;
  reg IsNaN_6U_10U_1_land_lpi_1_dfm_5;
  reg IsNaN_6U_10U_1_land_lpi_1_dfm_6;
  reg [9:0] FpMul_6U_10U_o_mant_lpi_1_dfm_7;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_18;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_19;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_20;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_21;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_22;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_23;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_24;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_25;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_26;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_18;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_19;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_20;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_21;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_22;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_23;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_24;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_25;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_26;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_27;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_28;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_29;
  reg [22:0] FpAdd_6U_10U_a_int_mant_p1_sva_2;
  reg [22:0] FpAdd_6U_10U_b_int_mant_p1_sva_2;
  reg inp_lookup_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_4;
  reg inp_lookup_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_5;
  reg [23:0] FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_4;
  reg [4:0] IntLeadZero_23U_leading_sign_23_0_rtn_sva_2;
  reg [5:0] IntLeadZero_35U_leading_sign_35_0_rtn_sva_2;
  reg FpFractionToFloat_35U_6U_10U_is_zero_lpi_1_dfm_5;
  reg [9:0] inp_lookup_else_if_a0_9_0_lpi_1_dfm_10;
  reg [5:0] IntLeadZero_35U_1_leading_sign_35_0_rtn_sva_2;
  reg inp_lookup_4_FpMantRNE_36U_11U_1_else_and_svs_2;
  reg [9:0] FpFractionToFloat_35U_6U_10U_1_o_mant_lpi_1_dfm_8;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_8;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_11;
  reg [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_8;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_9;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_10;
  reg [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_11;
  reg FpMul_6U_10U_1_lor_1_lpi_1_dfm_5;
  reg FpMul_6U_10U_1_lor_1_lpi_1_dfm_6;
  reg inp_lookup_4_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs_2;
  reg IsNaN_6U_10U_4_land_lpi_1_dfm_5;
  reg IsNaN_6U_10U_5_land_lpi_1_dfm_5;
  reg IsNaN_6U_10U_5_land_lpi_1_dfm_6;
  reg [9:0] FpMul_6U_10U_1_o_mant_lpi_1_dfm_9;
  reg [9:0] FpMul_6U_10U_1_o_mant_lpi_1_dfm_10;
  reg FpMul_6U_10U_2_lor_1_lpi_1_dfm_5;
  reg FpMul_6U_10U_2_lor_1_lpi_1_dfm_6;
  reg IsNaN_6U_10U_6_land_lpi_1_dfm_5;
  reg IsNaN_6U_10U_7_land_lpi_1_dfm_5;
  reg IsNaN_6U_10U_7_land_lpi_1_dfm_6;
  reg [9:0] FpMul_6U_10U_2_o_mant_lpi_1_dfm_7;
  reg [5:0] FpAdd_6U_10U_1_qr_lpi_1_dfm_5;
  reg [22:0] FpAdd_6U_10U_1_b_int_mant_p1_sva_2;
  reg inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4;
  reg inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5;
  reg [23:0] FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_4;
  reg inp_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_2;
  reg inp_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2;
  reg IsNaN_8U_23U_1_nor_itm_2;
  reg IsNaN_8U_23U_1_IsNaN_8U_23U_1_nand_itm_2;
  reg inp_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_5;
  reg inp_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_6;
  reg inp_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_7;
  reg inp_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2;
  reg IsZero_6U_10U_1_IsZero_6U_10U_1_and_itm_7;
  reg IsZero_6U_10U_1_IsZero_6U_10U_1_and_itm_8;
  reg IsZero_6U_10U_1_IsZero_6U_10U_1_and_itm_9;
  reg IsZero_6U_10U_1_IsZero_6U_10U_1_and_itm_10;
  reg IsZero_6U_10U_1_IsZero_6U_10U_1_and_itm_11;
  reg [6:0] FpMul_6U_10U_oelse_1_acc_itm_2;
  reg inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_11;
  reg inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_12;
  reg inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_13;
  reg inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_14;
  reg inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_15;
  reg inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_16;
  reg inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_3_or_itm_2;
  reg inp_lookup_1_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_itm_2;
  reg [29:0] inp_lookup_1_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_itm_2;
  reg inp_lookup_1_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_itm_2;
  reg [9:0] FpFractionToFloat_35U_6U_10U_if_else_mux_2_itm_2;
  reg [9:0] inp_lookup_1_FpMantWidthDec_6U_21U_10U_0U_0U_1_overflow_slc_FpMantRNE_22U_11U_i_data_1_20_1_19_10_itm;
  reg IsZero_6U_10U_7_IsZero_6U_10U_7_and_itm_2;
  reg FpMul_6U_10U_2_else_2_else_and_itm_2;
  reg FpMul_6U_10U_2_FpMul_6U_10U_2_and_itm_2;
  reg inp_lookup_1_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_itm_3;
  reg FpNormalize_6U_23U_1_if_or_itm_2;
  reg [9:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_itm;
  reg [9:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_itm_2;
  reg [50:0] inp_lookup_1_else_else_b1_mul_itm_2;
  wire signed [51:0] nl_inp_lookup_1_else_else_b1_mul_itm_2;
  reg inp_lookup_1_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2;
  reg inp_lookup_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_2;
  reg inp_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_5;
  reg inp_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_6;
  reg inp_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2;
  reg inp_lookup_2_IsZero_6U_10U_1_aif_IsZero_6U_10U_1_aelse_nor_itm_2;
  reg IsZero_6U_10U_1_IsZero_6U_10U_1_and_1_itm_6;
  reg IsZero_6U_10U_1_IsZero_6U_10U_1_and_1_itm_7;
  reg IsZero_6U_10U_1_IsZero_6U_10U_1_and_1_itm_8;
  reg IsZero_6U_10U_1_IsZero_6U_10U_1_and_1_itm_9;
  reg [6:0] FpMul_6U_10U_oelse_1_acc_1_itm_2;
  reg inp_lookup_2_IsZero_6U_10U_2_aif_IsZero_6U_10U_2_aelse_nor_itm_2;
  reg inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_10;
  reg inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_11;
  reg inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_12;
  reg inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_13;
  reg inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_14;
  reg inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_15;
  reg inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_3_or_itm_2;
  reg inp_lookup_2_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_itm_2;
  reg [29:0] inp_lookup_2_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_itm_2;
  reg inp_lookup_2_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_itm_2;
  reg [9:0] FpFractionToFloat_35U_6U_10U_if_else_mux_6_itm_2;
  reg IsZero_6U_10U_5_IsZero_6U_10U_5_and_1_itm_2;
  reg IsZero_6U_10U_7_IsZero_6U_10U_7_and_1_itm_2;
  reg FpMul_6U_10U_2_else_2_else_and_1_itm_2;
  reg FpMul_6U_10U_2_FpMul_6U_10U_2_and_16_itm_2;
  reg inp_lookup_2_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_itm_3;
  reg FpNormalize_6U_23U_1_if_or_1_itm_2;
  reg [9:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_1_itm;
  reg [9:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_1_itm_2;
  reg [50:0] inp_lookup_2_else_else_b1_mul_itm_2;
  wire signed [51:0] nl_inp_lookup_2_else_else_b1_mul_itm_2;
  reg inp_lookup_2_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2;
  reg inp_lookup_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_2;
  reg inp_lookup_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2;
  reg inp_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_5;
  reg inp_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_6;
  reg inp_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_7;
  reg inp_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2;
  reg IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_itm_7;
  reg IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_itm_8;
  reg IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_itm_9;
  reg IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_itm_10;
  reg IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_itm_11;
  reg [6:0] FpMul_6U_10U_oelse_1_acc_2_itm_2;
  reg inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_11;
  reg inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_12;
  reg inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_13;
  reg inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_14;
  reg inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_15;
  reg inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_16;
  reg inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_3_or_itm_2;
  reg inp_lookup_3_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_itm_2;
  reg [29:0] inp_lookup_3_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_itm_2;
  reg inp_lookup_3_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_itm_2;
  reg [9:0] FpFractionToFloat_35U_6U_10U_if_else_mux_10_itm_2;
  reg IsZero_6U_10U_7_IsZero_6U_10U_7_and_2_itm_2;
  reg FpMul_6U_10U_2_else_2_else_and_2_itm_2;
  reg FpMul_6U_10U_2_FpMul_6U_10U_2_and_17_itm_2;
  reg inp_lookup_3_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_itm_3;
  reg FpNormalize_6U_23U_1_if_or_2_itm_2;
  reg [9:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_2_itm;
  reg [9:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_2_itm_2;
  reg [50:0] inp_lookup_3_else_else_b1_mul_itm_2;
  wire signed [51:0] nl_inp_lookup_3_else_else_b1_mul_itm_2;
  reg inp_lookup_3_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2;
  reg inp_lookup_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_2;
  reg inp_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_5;
  reg inp_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_6;
  reg inp_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2;
  reg inp_lookup_4_IsZero_6U_10U_1_aif_IsZero_6U_10U_1_aelse_nor_itm_2;
  reg IsZero_6U_10U_1_IsZero_6U_10U_1_and_3_itm_6;
  reg IsZero_6U_10U_1_IsZero_6U_10U_1_and_3_itm_7;
  reg IsZero_6U_10U_1_IsZero_6U_10U_1_and_3_itm_8;
  reg IsZero_6U_10U_1_IsZero_6U_10U_1_and_3_itm_9;
  reg [6:0] FpMul_6U_10U_oelse_1_acc_3_itm_2;
  reg inp_lookup_4_IsZero_6U_10U_2_aif_IsZero_6U_10U_2_aelse_nor_itm_2;
  reg inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_10;
  reg inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_11;
  reg inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_12;
  reg inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_13;
  reg inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_14;
  reg inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_15;
  reg inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_16;
  reg inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_3_or_itm_2;
  reg inp_lookup_4_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_itm_2;
  reg [29:0] inp_lookup_4_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_itm_2;
  reg inp_lookup_4_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_itm_2;
  reg [9:0] FpFractionToFloat_35U_6U_10U_if_else_mux_14_itm_2;
  reg IsZero_6U_10U_5_IsZero_6U_10U_5_and_3_itm_2;
  reg [9:0] inp_lookup_4_FpMantWidthDec_6U_21U_10U_0U_0U_1_overflow_slc_FpMantRNE_22U_11U_i_data_1_20_1_19_10_itm;
  reg IsZero_6U_10U_7_IsZero_6U_10U_7_and_3_itm_2;
  reg FpMul_6U_10U_2_else_2_else_and_3_itm_2;
  reg FpMul_6U_10U_2_FpMul_6U_10U_2_and_18_itm_2;
  reg inp_lookup_4_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_itm_3;
  reg FpNormalize_6U_23U_1_if_or_3_itm_2;
  reg [9:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_3_itm;
  reg [9:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_3_itm_2;
  reg [50:0] inp_lookup_4_else_else_b1_mul_itm_2;
  wire signed [51:0] nl_inp_lookup_4_else_else_b1_mul_itm_2;
  reg inp_lookup_4_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2;
  reg inp_lookup_else_mux_485_itm_6;
  reg inp_lookup_else_mux_485_itm_7;
  reg inp_lookup_else_mux_485_itm_8;
  reg inp_lookup_else_mux_485_itm_9;
  reg inp_lookup_else_mux_485_itm_10;
  reg inp_lookup_mux_1057_itm_3;
  reg inp_lookup_mux_1057_itm_4;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_19_itm_5;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_19_itm_6;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_19_itm_7;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_19_itm_8;
  reg inp_lookup_else_mux_491_itm_5;
  reg inp_lookup_else_mux_491_itm_6;
  reg inp_lookup_else_mux_491_itm_7;
  reg inp_lookup_else_mux_491_itm_8;
  reg inp_lookup_else_mux_362_itm_6;
  reg inp_lookup_else_mux_362_itm_7;
  reg inp_lookup_else_mux_362_itm_8;
  reg inp_lookup_else_mux_362_itm_9;
  reg inp_lookup_else_mux_362_itm_10;
  reg inp_lookup_mux_791_itm_3;
  reg inp_lookup_mux_791_itm_4;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_14_itm_5;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_14_itm_6;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_14_itm_7;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_14_itm_8;
  reg inp_lookup_else_mux_368_itm_5;
  reg inp_lookup_else_mux_368_itm_6;
  reg inp_lookup_else_mux_368_itm_7;
  reg inp_lookup_else_mux_368_itm_8;
  reg inp_lookup_else_mux_239_itm_6;
  reg inp_lookup_else_mux_239_itm_7;
  reg inp_lookup_else_mux_239_itm_8;
  reg inp_lookup_else_mux_239_itm_9;
  reg inp_lookup_else_mux_239_itm_10;
  reg inp_lookup_mux_525_itm_3;
  reg inp_lookup_mux_525_itm_4;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_9_itm_5;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_9_itm_6;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_9_itm_7;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_9_itm_8;
  reg inp_lookup_else_mux_245_itm_5;
  reg inp_lookup_else_mux_245_itm_6;
  reg inp_lookup_else_mux_245_itm_7;
  reg inp_lookup_else_mux_245_itm_8;
  reg inp_lookup_else_mux_116_itm_6;
  reg inp_lookup_else_mux_116_itm_7;
  reg inp_lookup_else_mux_116_itm_8;
  reg inp_lookup_else_mux_116_itm_9;
  reg inp_lookup_else_mux_116_itm_10;
  reg inp_lookup_mux_259_itm_3;
  reg inp_lookup_mux_259_itm_4;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_4_itm_5;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_4_itm_6;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_4_itm_7;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_4_itm_8;
  reg inp_lookup_else_mux_122_itm_5;
  reg inp_lookup_else_mux_122_itm_6;
  reg inp_lookup_else_mux_122_itm_7;
  reg inp_lookup_else_mux_122_itm_8;
  reg FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_st_2;
  reg [1:0] cfg_precision_1_sva_st_80;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_st_3;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_st_4;
  reg [1:0] cfg_precision_1_sva_st_81;
  reg FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_1_st_2;
  reg inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4;
  reg inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5;
  reg [1:0] cfg_precision_1_sva_st_82;
  reg [1:0] cfg_precision_1_sva_st_83;
  reg IsNaN_8U_23U_2_land_1_lpi_1_dfm_st_6;
  reg IsNaN_8U_23U_2_land_1_lpi_1_dfm_st_7;
  reg [1:0] cfg_precision_1_sva_st_84;
  reg inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2;
  reg [1:0] cfg_precision_1_sva_st_85;
  reg [1:0] cfg_precision_1_sva_st_86;
  reg FpMul_6U_10U_lor_6_lpi_1_dfm_st_2;
  reg inp_lookup_1_FpMul_6U_10U_else_2_else_slc_FpMul_6U_10U_p_mant_p1_21_itm_2;
  reg [1:0] cfg_precision_1_sva_st_87;
  reg [1:0] cfg_precision_1_sva_st_88;
  reg [1:0] cfg_precision_1_sva_st_89;
  reg inp_lookup_1_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2;
  reg FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_1_sva_st_2;
  reg IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_13;
  reg IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_14;
  reg IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_15;
  reg IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_16;
  reg IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_17;
  reg IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_18;
  reg IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_19;
  reg IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_20;
  reg IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_21;
  reg IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_22;
  reg IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_23;
  reg IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_24;
  reg [1:0] cfg_precision_1_sva_st_90;
  reg [34:0] inp_lookup_1_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_3;
  reg [1:0] cfg_precision_1_sva_st_91;
  reg [34:0] inp_lookup_1_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_4;
  reg FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_3;
  reg FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_4;
  reg FpMul_6U_10U_2_lor_6_lpi_1_dfm_st_3;
  reg FpMul_6U_10U_2_lor_6_lpi_1_dfm_st_4;
  reg inp_lookup_1_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4;
  reg inp_lookup_1_FpMul_6U_10U_2_else_2_else_slc_FpMul_6U_10U_2_p_mant_p1_21_itm_2;
  reg FpMul_6U_10U_2_else_2_else_if_if_slc_FpMul_6U_10U_2_else_2_else_if_if_acc_1_5_mdf_1_sva_st_1;
  reg inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4;
  reg inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5;
  reg inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6;
  reg IsNaN_6U_10U_8_land_1_lpi_1_dfm_st_3;
  reg FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_st_2;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_st_4;
  reg FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_1_st_2;
  reg inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4;
  reg inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5;
  reg IsNaN_8U_23U_2_land_2_lpi_1_dfm_st_6;
  reg IsNaN_8U_23U_2_land_2_lpi_1_dfm_st_7;
  reg inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2;
  reg [1:0] cfg_precision_1_sva_st_100;
  reg FpMul_6U_10U_lor_7_lpi_1_dfm_st_2;
  reg inp_lookup_2_FpMul_6U_10U_else_2_else_slc_FpMul_6U_10U_p_mant_p1_21_itm_2;
  reg [1:0] cfg_precision_1_sva_st_101;
  reg [1:0] cfg_precision_1_sva_st_102;
  reg [1:0] cfg_precision_1_sva_st_103;
  reg inp_lookup_2_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2;
  reg FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_2_sva_st_2;
  reg IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_13;
  reg IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_14;
  reg IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_15;
  reg IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_16;
  reg IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_17;
  reg IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_18;
  reg IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_19;
  reg IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_20;
  reg IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_21;
  reg IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_22;
  reg IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_23;
  reg IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_24;
  reg [34:0] inp_lookup_2_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_3;
  reg [34:0] inp_lookup_2_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_4;
  reg FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_3;
  reg FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_4;
  reg FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_3;
  reg FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_4;
  reg inp_lookup_2_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4;
  reg inp_lookup_2_FpMul_6U_10U_2_else_2_else_slc_FpMul_6U_10U_2_p_mant_p1_21_itm_2;
  reg FpMul_6U_10U_2_else_2_else_if_if_slc_FpMul_6U_10U_2_else_2_else_if_if_acc_1_5_mdf_2_sva_st_1;
  reg inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4;
  reg inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5;
  reg inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6;
  reg IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_4;
  reg IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_5;
  reg FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_st_2;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_st_4;
  reg FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_1_st_2;
  reg inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4;
  reg inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5;
  reg IsNaN_8U_23U_2_land_3_lpi_1_dfm_st_6;
  reg IsNaN_8U_23U_2_land_3_lpi_1_dfm_st_7;
  reg inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2;
  reg [1:0] cfg_precision_1_sva_st_112;
  reg FpMul_6U_10U_lor_8_lpi_1_dfm_st_2;
  reg inp_lookup_3_FpMul_6U_10U_else_2_else_slc_FpMul_6U_10U_p_mant_p1_21_itm_2;
  reg [1:0] cfg_precision_1_sva_st_113;
  reg [1:0] cfg_precision_1_sva_st_114;
  reg [1:0] cfg_precision_1_sva_st_115;
  reg inp_lookup_3_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2;
  reg FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_3_sva_st_2;
  reg IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_13;
  reg IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_14;
  reg IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_15;
  reg IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_16;
  reg IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_17;
  reg IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_18;
  reg IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_19;
  reg IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_20;
  reg IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_21;
  reg IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_22;
  reg IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_23;
  reg IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_24;
  reg [34:0] inp_lookup_3_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_3;
  reg [34:0] inp_lookup_3_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_4;
  reg FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_3;
  reg FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_4;
  reg FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_3;
  reg FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_4;
  reg inp_lookup_3_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4;
  reg inp_lookup_3_FpMul_6U_10U_2_else_2_else_slc_FpMul_6U_10U_2_p_mant_p1_21_itm_2;
  reg FpMul_6U_10U_2_else_2_else_if_if_slc_FpMul_6U_10U_2_else_2_else_if_if_acc_1_5_mdf_3_sva_st_1;
  reg inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4;
  reg inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5;
  reg inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6;
  reg IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_4;
  reg IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_5;
  reg FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2;
  reg IsNaN_8U_23U_land_lpi_1_dfm_st_4;
  reg FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_1_st_2;
  reg inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4;
  reg inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5;
  reg IsNaN_8U_23U_2_land_lpi_1_dfm_st_6;
  reg IsNaN_8U_23U_2_land_lpi_1_dfm_st_7;
  reg IsNaN_8U_23U_2_land_lpi_1_dfm_st_8;
  reg inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2;
  reg [1:0] cfg_precision_1_sva_st_124;
  reg FpMul_6U_10U_lor_1_lpi_1_dfm_st_2;
  reg inp_lookup_4_FpMul_6U_10U_else_2_else_slc_FpMul_6U_10U_p_mant_p1_21_itm_2;
  reg [1:0] cfg_precision_1_sva_st_125;
  reg [1:0] cfg_precision_1_sva_st_126;
  reg [1:0] cfg_precision_1_sva_st_127;
  reg inp_lookup_4_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2;
  reg FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_sva_st_2;
  reg IsNaN_6U_10U_2_land_lpi_1_dfm_st_13;
  reg IsNaN_6U_10U_2_land_lpi_1_dfm_st_14;
  reg IsNaN_6U_10U_2_land_lpi_1_dfm_st_15;
  reg IsNaN_6U_10U_2_land_lpi_1_dfm_st_16;
  reg IsNaN_6U_10U_2_land_lpi_1_dfm_st_17;
  reg IsNaN_6U_10U_2_land_lpi_1_dfm_st_18;
  reg IsNaN_6U_10U_2_land_lpi_1_dfm_st_19;
  reg IsNaN_6U_10U_2_land_lpi_1_dfm_st_20;
  reg IsNaN_6U_10U_2_land_lpi_1_dfm_st_21;
  reg IsNaN_6U_10U_2_land_lpi_1_dfm_st_22;
  reg IsNaN_6U_10U_2_land_lpi_1_dfm_st_23;
  reg [34:0] inp_lookup_4_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_3;
  reg [34:0] inp_lookup_4_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_4;
  reg FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_3;
  reg FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_4;
  reg FpMul_6U_10U_2_lor_1_lpi_1_dfm_st_3;
  reg FpMul_6U_10U_2_lor_1_lpi_1_dfm_st_4;
  reg inp_lookup_4_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4;
  reg inp_lookup_4_FpMul_6U_10U_2_else_2_else_slc_FpMul_6U_10U_2_p_mant_p1_21_itm_2;
  reg FpMul_6U_10U_2_else_2_else_if_if_slc_FpMul_6U_10U_2_else_2_else_if_if_acc_1_5_mdf_sva_st_2;
  reg inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4;
  reg inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5;
  reg IsNaN_6U_10U_8_land_lpi_1_dfm_st_4;
  reg IsNaN_6U_10U_8_land_lpi_1_dfm_st_5;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3_0;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_3_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_3_0;
  reg [3:0] FpAdd_6U_10U_qr_2_lpi_1_dfm_3_0;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_3_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_3_0;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3_0;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_3_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_3_0;
  reg [3:0] FpAdd_6U_10U_qr_3_lpi_1_dfm_3_0;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_3_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_3_0;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3_0;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_3_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_3_0;
  reg [3:0] FpAdd_6U_10U_qr_4_lpi_1_dfm_3_0;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_3_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_3_0;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3_0;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_3_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_3_0;
  reg [3:0] FpAdd_6U_10U_qr_lpi_1_dfm_3_0;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_3_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_3_0;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_5_4_1;
  reg [3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_5_3_0_1;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_6_4_1;
  reg [3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_6_3_0_1;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_7_4_1;
  reg [3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_7_3_0_1;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_8_4_1;
  reg [3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_8_3_0_1;
  reg inp_lookup_else_if_a0_15_10_lpi_1_dfm_6_5_1;
  reg [4:0] inp_lookup_else_if_a0_15_10_lpi_1_dfm_6_4_0_1;
  reg [30:0] IntSaturation_51U_32U_o_lpi_1_dfm_11_30_0_1;
  reg [30:0] IntSaturation_51U_32U_o_lpi_1_dfm_12_30_0_1;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_5_4_1;
  reg [3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_5_3_0_1;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_6_4_1;
  reg [3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_6_3_0_1;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_7_4_1;
  reg [3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_7_3_0_1;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_8_4_1;
  reg [3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_8_3_0_1;
  reg inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_6_5_1;
  reg [4:0] inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_6_4_0_1;
  reg [30:0] IntSaturation_51U_32U_o_3_lpi_1_dfm_11_30_0_1;
  reg [30:0] IntSaturation_51U_32U_o_3_lpi_1_dfm_12_30_0_1;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_5_4_1;
  reg [3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_5_3_0_1;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_6_4_1;
  reg [3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_6_3_0_1;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_7_4_1;
  reg [3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_7_3_0_1;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_8_4_1;
  reg [3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_8_3_0_1;
  reg inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_6_5_1;
  reg [4:0] inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_6_4_0_1;
  reg [30:0] IntSaturation_51U_32U_o_2_lpi_1_dfm_11_30_0_1;
  reg [30:0] IntSaturation_51U_32U_o_2_lpi_1_dfm_12_30_0_1;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_5_4_1;
  reg [3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_5_3_0_1;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_6_4_1;
  reg [3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_6_3_0_1;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_7_4_1;
  reg [3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_7_3_0_1;
  reg FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_8_4_1;
  reg [3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_8_3_0_1;
  reg inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_5_1;
  reg [4:0] inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_4_0_1;
  reg [30:0] IntSaturation_51U_32U_o_1_lpi_1_dfm_11_30_0_1;
  reg [30:0] IntSaturation_51U_32U_o_1_lpi_1_dfm_12_30_0_1;
  reg [344:0] chn_inp_in_crt_sva_1_739_395_1;
  reg [63:0] chn_inp_in_crt_sva_1_331_268_1;
  reg [127:0] chn_inp_in_crt_sva_1_127_0_1;
  reg [3:0] chn_inp_in_crt_sva_2_739_736_1;
  reg chn_inp_in_crt_sva_2_395_1;
  reg chn_inp_in_crt_sva_2_379_1;
  reg chn_inp_in_crt_sva_2_363_1;
  reg chn_inp_in_crt_sva_2_347_1;
  reg [63:0] chn_inp_in_crt_sva_2_331_268_1;
  reg [127:0] chn_inp_in_crt_sva_2_127_0_1;
  reg [3:0] chn_inp_in_crt_sva_3_739_736_1;
  reg [63:0] chn_inp_in_crt_sva_3_331_268_1;
  reg [127:0] chn_inp_in_crt_sva_3_127_0_1;
  reg [3:0] chn_inp_in_crt_sva_4_739_736_1;
  reg chn_inp_in_crt_sva_4_459_1;
  reg chn_inp_in_crt_sva_4_443_1;
  reg chn_inp_in_crt_sva_4_427_1;
  reg chn_inp_in_crt_sva_4_411_1;
  reg chn_inp_in_crt_sva_4_331_1;
  reg chn_inp_in_crt_sva_4_315_1;
  reg chn_inp_in_crt_sva_4_299_1;
  reg chn_inp_in_crt_sva_4_283_1;
  reg [127:0] chn_inp_in_crt_sva_4_127_0_1;
  reg [3:0] chn_inp_in_crt_sva_5_739_736_1;
  reg chn_inp_in_crt_sva_5_459_1;
  reg chn_inp_in_crt_sva_5_443_1;
  reg chn_inp_in_crt_sva_5_427_1;
  reg chn_inp_in_crt_sva_5_411_1;
  reg chn_inp_in_crt_sva_5_331_1;
  reg chn_inp_in_crt_sva_5_315_1;
  reg chn_inp_in_crt_sva_5_299_1;
  reg chn_inp_in_crt_sva_5_283_1;
  reg [3:0] chn_inp_in_crt_sva_6_739_736_1;
  reg chn_inp_in_crt_sva_6_459_1;
  reg chn_inp_in_crt_sva_6_443_1;
  reg chn_inp_in_crt_sva_6_427_1;
  reg chn_inp_in_crt_sva_6_411_1;
  reg chn_inp_in_crt_sva_6_331_1;
  reg chn_inp_in_crt_sva_6_315_1;
  reg chn_inp_in_crt_sva_6_299_1;
  reg chn_inp_in_crt_sva_6_283_1;
  reg [3:0] chn_inp_in_crt_sva_7_739_736_1;
  reg chn_inp_in_crt_sva_7_459_1;
  reg chn_inp_in_crt_sva_7_443_1;
  reg chn_inp_in_crt_sva_7_427_1;
  reg chn_inp_in_crt_sva_7_411_1;
  reg chn_inp_in_crt_sva_7_331_1;
  reg chn_inp_in_crt_sva_7_315_1;
  reg chn_inp_in_crt_sva_7_299_1;
  reg chn_inp_in_crt_sva_7_283_1;
  reg [3:0] chn_inp_in_crt_sva_8_739_736_1;
  reg chn_inp_in_crt_sva_8_331_1;
  reg chn_inp_in_crt_sva_8_315_1;
  reg chn_inp_in_crt_sva_8_299_1;
  reg chn_inp_in_crt_sva_8_283_1;
  reg [3:0] chn_inp_in_crt_sva_9_739_736_1;
  reg chn_inp_in_crt_sva_9_331_1;
  reg chn_inp_in_crt_sva_9_315_1;
  reg chn_inp_in_crt_sva_9_299_1;
  reg chn_inp_in_crt_sva_9_283_1;
  reg [3:0] chn_inp_in_crt_sva_10_739_736_1;
  reg chn_inp_in_crt_sva_10_331_1;
  reg chn_inp_in_crt_sva_10_315_1;
  reg chn_inp_in_crt_sva_10_299_1;
  reg chn_inp_in_crt_sva_10_283_1;
  reg [3:0] chn_inp_in_crt_sva_11_739_736_1;
  reg [3:0] chn_inp_in_crt_sva_12_739_736_1;
  reg [48:0] FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_3_49_1_1;
  reg FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_10_5_1;
  reg [4:0] FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_10_4_0_1;
  reg [4:0] FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_11_4_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_6_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_6_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_7_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_7_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_8_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_8_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_9_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_9_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_10_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_10_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_11_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_11_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_12_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_12_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_13_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_14_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_14_0_1;
  reg [3:0] FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_3_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_6_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_6_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_7_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_7_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_8_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_8_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_9_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_9_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_10_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_10_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_11_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_11_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_12_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_12_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_13_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_13_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_14_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_14_0_1;
  reg [3:0] FpAdd_6U_10U_qr_2_lpi_1_dfm_3_3_0_1;
  reg [3:0] FpAdd_6U_10U_qr_2_lpi_1_dfm_4_3_0_1;
  reg [66:0] IntSignedShiftRight_50U_5U_32U_mbits_fixed_1_sva_1_80_14_1;
  reg [4:0] inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_7_4_0_1;
  reg inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_8_5_1;
  reg [4:0] inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_8_4_0_1;
  reg FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_6_5_1;
  reg [4:0] FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_6_4_0_1;
  reg [4:0] FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_7_4_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_6_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_6_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_7_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_8_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_9_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_6_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_6_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_7_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_7_0_1;
  reg FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_6_5_1;
  reg [3:0] FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_6_3_0_1;
  reg FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_7_5_1;
  reg FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_7_4_1;
  reg [3:0] FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_7_3_0_1;
  reg FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_8_5_1;
  reg FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_8_4_1;
  reg FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_5_1;
  reg FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_4_1;
  reg [3:0] FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_3_0_1;
  reg FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_7_5_1;
  reg FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_7_4_1;
  reg [3:0] FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_7_3_0_1;
  reg FpAdd_6U_10U_1_qr_2_lpi_1_dfm_3_5_1;
  reg FpAdd_6U_10U_1_qr_2_lpi_1_dfm_3_4_1;
  reg [3:0] FpAdd_6U_10U_1_qr_2_lpi_1_dfm_3_3_0_1;
  reg FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_5_1;
  reg FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_4_1;
  reg [3:0] FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_3_0_1;
  reg [48:0] FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_3_49_1_1;
  reg FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_10_5_1;
  reg [4:0] FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_10_4_0_1;
  reg [4:0] FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_11_4_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_6_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_6_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_7_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_7_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_8_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_8_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_9_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_9_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_10_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_10_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_11_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_11_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_12_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_12_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_13_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_14_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_14_0_1;
  reg [3:0] FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_3_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_6_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_6_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_7_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_7_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_8_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_8_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_9_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_9_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_10_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_10_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_11_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_11_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_12_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_12_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_13_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_13_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_14_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_14_0_1;
  reg [3:0] FpAdd_6U_10U_qr_3_lpi_1_dfm_3_3_0_1;
  reg [3:0] FpAdd_6U_10U_qr_3_lpi_1_dfm_4_3_0_1;
  reg [66:0] IntSignedShiftRight_50U_5U_32U_mbits_fixed_2_sva_1_80_14_1;
  reg [4:0] inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_7_4_0_1;
  reg inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_8_5_1;
  reg [4:0] inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_8_4_0_1;
  reg FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_6_5_1;
  reg [4:0] FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_6_4_0_1;
  reg [4:0] FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_7_4_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_6_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_6_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_7_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_8_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_9_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_6_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_6_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_7_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_7_0_1;
  reg FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_6_5_1;
  reg [3:0] FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_6_3_0_1;
  reg FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_7_5_1;
  reg FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_7_4_1;
  reg [3:0] FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_7_3_0_1;
  reg FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_8_5_1;
  reg FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_8_4_1;
  reg FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_5_1;
  reg FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_4_1;
  reg [3:0] FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_3_0_1;
  reg FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_7_5_1;
  reg FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_7_4_1;
  reg [3:0] FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_7_3_0_1;
  reg FpAdd_6U_10U_1_qr_3_lpi_1_dfm_3_5_1;
  reg FpAdd_6U_10U_1_qr_3_lpi_1_dfm_3_4_1;
  reg [3:0] FpAdd_6U_10U_1_qr_3_lpi_1_dfm_3_3_0_1;
  reg FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_5_1;
  reg FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_4_1;
  reg [3:0] FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_3_0_1;
  reg [48:0] FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_3_49_1_1;
  reg FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_10_5_1;
  reg [4:0] FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_10_4_0_1;
  reg [4:0] FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_11_4_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_6_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_6_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_7_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_7_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_8_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_8_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_9_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_9_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_10_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_10_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_11_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_11_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_12_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_12_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_13_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_14_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_14_0_1;
  reg [3:0] FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_3_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_6_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_6_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_7_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_7_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_8_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_8_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_9_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_9_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_10_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_10_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_11_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_11_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_12_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_12_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_13_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_13_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_14_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_14_0_1;
  reg [3:0] FpAdd_6U_10U_qr_4_lpi_1_dfm_3_3_0_1;
  reg [3:0] FpAdd_6U_10U_qr_4_lpi_1_dfm_4_3_0_1;
  reg [66:0] IntSignedShiftRight_50U_5U_32U_mbits_fixed_3_sva_1_80_14_1;
  reg [4:0] inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_7_4_0_1;
  reg inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_8_5_1;
  reg [4:0] inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_8_4_0_1;
  reg FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_6_5_1;
  reg [4:0] FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_6_4_0_1;
  reg [4:0] FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_7_4_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_6_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_6_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_7_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_8_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_9_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_6_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_6_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_7_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_7_0_1;
  reg FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_6_5_1;
  reg [3:0] FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_6_3_0_1;
  reg FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_7_5_1;
  reg FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_7_4_1;
  reg [3:0] FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_7_3_0_1;
  reg FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_8_5_1;
  reg FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_8_4_1;
  reg FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_5_1;
  reg FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_4_1;
  reg [3:0] FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_3_0_1;
  reg FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_7_5_1;
  reg FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_7_4_1;
  reg [3:0] FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_7_3_0_1;
  reg FpAdd_6U_10U_1_qr_4_lpi_1_dfm_3_5_1;
  reg FpAdd_6U_10U_1_qr_4_lpi_1_dfm_3_4_1;
  reg [3:0] FpAdd_6U_10U_1_qr_4_lpi_1_dfm_3_3_0_1;
  reg FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_5_1;
  reg FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_4_1;
  reg [3:0] FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_3_0_1;
  reg [48:0] FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_3_49_1_1;
  reg FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_10_5_1;
  reg [4:0] FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_10_4_0_1;
  reg [4:0] FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_11_4_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_6_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_6_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_7_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_7_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_8_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_8_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_9_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_9_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_10_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_10_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_11_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_11_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_12_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_12_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_13_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_14_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_14_0_1;
  reg [3:0] FpMul_6U_10U_o_expo_lpi_1_dfm_6_3_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_6_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_6_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_7_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_7_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_8_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_8_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_9_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_9_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_10_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_10_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_11_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_11_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_12_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_12_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_13_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_13_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_14_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_14_0_1;
  reg [3:0] FpAdd_6U_10U_qr_lpi_1_dfm_3_3_0_1;
  reg [3:0] FpAdd_6U_10U_qr_lpi_1_dfm_4_3_0_1;
  reg [66:0] IntSignedShiftRight_50U_5U_32U_mbits_fixed_sva_1_80_14_1;
  reg [4:0] inp_lookup_else_if_a0_15_10_lpi_1_dfm_7_4_0_1;
  reg inp_lookup_else_if_a0_15_10_lpi_1_dfm_8_5_1;
  reg [4:0] inp_lookup_else_if_a0_15_10_lpi_1_dfm_8_4_0_1;
  reg FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_6_5_1;
  reg [4:0] FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_6_4_0_1;
  reg [4:0] FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_7_4_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_6_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_6_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_7_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_7_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_8_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_8_0;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_9_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_6_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_6_0_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_7_1_1;
  reg FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_7_0_1;
  reg FpMul_6U_10U_1_o_expo_lpi_1_dfm_6_5_1;
  reg [3:0] FpMul_6U_10U_1_o_expo_lpi_1_dfm_6_3_0_1;
  reg FpMul_6U_10U_1_o_expo_lpi_1_dfm_7_5_1;
  reg FpMul_6U_10U_1_o_expo_lpi_1_dfm_7_4_1;
  reg [3:0] FpMul_6U_10U_1_o_expo_lpi_1_dfm_7_3_0_1;
  reg FpMul_6U_10U_1_o_expo_lpi_1_dfm_8_5_1;
  reg FpMul_6U_10U_1_o_expo_lpi_1_dfm_8_4_1;
  reg FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_5_1;
  reg FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_4_1;
  reg [3:0] FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_3_0_1;
  reg FpMul_6U_10U_2_o_expo_lpi_1_dfm_7_5_1;
  reg FpMul_6U_10U_2_o_expo_lpi_1_dfm_7_4_1;
  reg [3:0] FpMul_6U_10U_2_o_expo_lpi_1_dfm_7_3_0_1;
  reg FpAdd_6U_10U_1_qr_lpi_1_dfm_3_5_1;
  reg FpAdd_6U_10U_1_qr_lpi_1_dfm_3_4_1;
  reg [3:0] FpAdd_6U_10U_1_qr_lpi_1_dfm_3_3_0_1;
  reg FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_5_1;
  reg FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_4_1;
  reg [3:0] FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_3_0_1;
  wire FpAdd_6U_10U_mux_50_tmp_23;
  wire FpAdd_6U_10U_mux_34_tmp_23;
  wire FpAdd_6U_10U_mux_18_tmp_23;
  wire FpAdd_6U_10U_mux_2_tmp_23;
  wire FpFractionToFloat_35U_6U_10U_1_and_2_cse;
  wire FpFractionToFloat_35U_6U_10U_1_and_1_cse;
  wire main_stage_en_1;
  wire IsZero_5U_10U_IsZero_5U_10U_nor_cse_sva;
  wire IsZero_5U_10U_3_IsZero_5U_10U_3_nor_cse_sva;
  wire IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_sva;
  wire IsZero_5U_10U_IsZero_5U_10U_nor_cse_3_sva;
  wire IsZero_5U_10U_3_IsZero_5U_10U_3_nor_cse_3_sva;
  wire IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_3_sva;
  wire IsZero_5U_10U_IsZero_5U_10U_nor_cse_2_sva;
  wire IsZero_5U_10U_3_IsZero_5U_10U_3_nor_cse_2_sva;
  wire IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_2_sva;
  wire IsZero_5U_10U_IsZero_5U_10U_nor_cse_1_sva;
  wire IsZero_5U_10U_3_IsZero_5U_10U_3_nor_cse_1_sva;
  wire IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_1_sva;
  wire FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_3_5_mx0w0;
  wire FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_3_5_mx0w0;
  wire FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_3_5_mx0w0;
  wire FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_3_5_mx0w0;
  wire FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0;
  wire FpMul_6U_10U_2_FpMul_6U_10U_2_nor_3_ssc;
  wire FpAdd_8U_23U_is_inf_lpi_1_dfm;
  wire FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0;
  wire FpMul_6U_10U_2_FpMul_6U_10U_2_nor_2_ssc;
  wire FpAdd_8U_23U_is_inf_3_lpi_1_dfm;
  wire FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0;
  wire FpMul_6U_10U_2_FpMul_6U_10U_2_nor_1_ssc;
  wire FpAdd_8U_23U_is_inf_2_lpi_1_dfm;
  wire FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0;
  wire FpMul_6U_10U_2_FpMul_6U_10U_2_nor_ssc;
  wire FpAdd_8U_23U_is_inf_1_lpi_1_dfm;
  wire [5:0] FpMul_6U_10U_1_p_expo_lpi_1_dfm_1_mx0;
  wire [5:0] FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_sva_1;
  wire [6:0] nl_FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_sva_1;
  wire FpMantWidthDec_6U_21U_10U_0U_0U_1_if_1_unequal_tmp_3;
  wire [5:0] FpMul_6U_10U_1_p_expo_3_lpi_1_dfm_1_mx0;
  wire [5:0] FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_3_sva_1;
  wire [6:0] nl_FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_3_sva_1;
  wire FpMantWidthDec_6U_21U_10U_0U_0U_1_if_1_unequal_tmp_2;
  wire [5:0] FpMul_6U_10U_1_p_expo_2_lpi_1_dfm_1_mx0;
  wire [5:0] FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_2_sva_1;
  wire [6:0] nl_FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_2_sva_1;
  wire FpMantWidthDec_6U_21U_10U_0U_0U_1_if_1_unequal_tmp_1;
  wire [5:0] FpMul_6U_10U_1_p_expo_1_lpi_1_dfm_1_mx0;
  wire [5:0] FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_1_sva_1;
  wire [6:0] nl_FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_1_sva_1;
  wire FpMantWidthDec_6U_21U_10U_0U_0U_1_if_1_unequal_tmp;
  wire FpAdd_8U_23U_1_is_inf_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_11_m1c;
  wire FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_9_m1c;
  wire FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_7_m1c;
  wire FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_5_m1c;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_else_and_3_tmp;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_lpi_1_dfm_3;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_else_and_2_tmp;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_3_lpi_1_dfm_3;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_else_and_1_tmp;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_2_lpi_1_dfm_3;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_else_and_tmp;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_1_lpi_1_dfm_3;
  wire FpMantRNE_22U_11U_else_carry_sva;
  wire FpMantRNE_22U_11U_else_carry_3_sva;
  wire FpMantRNE_22U_11U_else_carry_2_sva;
  wire FpMantRNE_22U_11U_else_carry_1_sva;
  wire IsNaN_6U_23U_IsNaN_6U_23U_nand_3_cse;
  wire FpAdd_6U_10U_and_34_ssc;
  wire FpAdd_6U_10U_is_inf_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_FpAdd_6U_10U_nor_11_m1c;
  wire FpAdd_6U_10U_and_3_tmp;
  wire FpAdd_6U_10U_and_22_ssc;
  wire IsNaN_6U_23U_IsNaN_6U_23U_nand_2_cse;
  wire FpAdd_6U_10U_and_32_ssc;
  wire FpAdd_6U_10U_is_inf_3_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_FpAdd_6U_10U_nor_9_m1c;
  wire FpAdd_6U_10U_and_2_tmp;
  wire FpAdd_6U_10U_and_16_ssc;
  wire IsNaN_6U_23U_IsNaN_6U_23U_nand_1_cse;
  wire FpAdd_6U_10U_and_30_ssc;
  wire FpAdd_6U_10U_is_inf_2_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_FpAdd_6U_10U_nor_7_m1c;
  wire FpAdd_6U_10U_and_1_tmp;
  wire FpAdd_6U_10U_and_10_ssc;
  wire IsNaN_6U_23U_IsNaN_6U_23U_nand_cse;
  wire FpAdd_6U_10U_and_28_ssc;
  wire FpAdd_6U_10U_is_inf_1_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_FpAdd_6U_10U_nor_5_m1c;
  wire FpAdd_6U_10U_and_tmp;
  wire FpAdd_6U_10U_and_4_ssc;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_3_0_mx0w0;
  wire IsDenorm_5U_10U_3_land_lpi_1_dfm;
  wire IsInf_5U_10U_3_land_lpi_1_dfm;
  wire IsInf_5U_10U_3_IsInf_5U_10U_3_and_cse_sva;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_3_0_mx0w0;
  wire IsDenorm_5U_10U_3_land_3_lpi_1_dfm;
  wire IsInf_5U_10U_3_land_3_lpi_1_dfm;
  wire IsInf_5U_10U_3_IsInf_5U_10U_3_and_cse_3_sva;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_3_0_mx0w0;
  wire IsDenorm_5U_10U_3_land_2_lpi_1_dfm;
  wire IsInf_5U_10U_3_land_2_lpi_1_dfm;
  wire IsInf_5U_10U_3_IsInf_5U_10U_3_and_cse_2_sva;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_3_0_mx0w0;
  wire IsDenorm_5U_10U_3_land_1_lpi_1_dfm;
  wire IsInf_5U_10U_3_land_1_lpi_1_dfm;
  wire IsInf_5U_10U_3_IsInf_5U_10U_3_and_cse_1_sva;
  wire FpFractionToFloat_35U_6U_10U_is_zero_lpi_1_dfm_mx0w0;
  wire FpFractionToFloat_35U_6U_10U_is_zero_3_lpi_1_dfm_mx0w0;
  wire FpFractionToFloat_35U_6U_10U_is_zero_2_lpi_1_dfm_mx0w0;
  wire FpFractionToFloat_35U_6U_10U_is_zero_1_lpi_1_dfm_mx0w0;
  wire [5:0] FpMul_6U_10U_2_p_expo_lpi_1_dfm_1_mx0;
  wire [5:0] FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_sva_1;
  wire [6:0] nl_FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_sva_1;
  wire FpMantWidthDec_6U_21U_10U_0U_0U_2_if_1_unequal_tmp_3;
  wire [5:0] FpMul_6U_10U_2_p_expo_3_lpi_1_dfm_1_mx0;
  wire [5:0] FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_3_sva_1;
  wire [6:0] nl_FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_3_sva_1;
  wire FpMantWidthDec_6U_21U_10U_0U_0U_2_if_1_unequal_tmp_2;
  wire [5:0] FpMul_6U_10U_2_p_expo_2_lpi_1_dfm_1_mx0;
  wire [5:0] FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_2_sva_1;
  wire [6:0] nl_FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_2_sva_1;
  wire FpMantWidthDec_6U_21U_10U_0U_0U_2_if_1_unequal_tmp_1;
  wire [5:0] FpMul_6U_10U_2_p_expo_1_lpi_1_dfm_1_mx0;
  wire [5:0] FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_1_sva_1;
  wire [6:0] nl_FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_1_sva_1;
  wire FpMantWidthDec_6U_21U_10U_0U_0U_2_if_1_unequal_tmp;
  wire FpMantRNE_24U_11U_else_carry_sva_mx0w1;
  wire FpAdd_8U_23U_1_and_3_tmp;
  wire FpMantRNE_24U_11U_else_carry_3_sva_mx0w1;
  wire FpAdd_8U_23U_1_and_2_tmp;
  wire FpMantRNE_24U_11U_else_carry_2_sva_mx0w1;
  wire FpAdd_8U_23U_1_and_1_tmp;
  wire FpMantRNE_24U_11U_else_carry_1_sva;
  wire FpAdd_8U_23U_1_and_tmp;
  wire FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_5_mx0w0;
  wire FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_4_mx0w0;
  wire FpAdd_6U_10U_1_and_34_ssc;
  wire FpAdd_6U_10U_1_and_3_tmp;
  wire FpAdd_6U_10U_1_is_inf_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_11_m1c;
  wire FpAdd_6U_10U_1_and_22_ssc;
  wire FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_5_mx0w0;
  wire FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_4_mx0w0;
  wire FpAdd_6U_10U_1_and_32_ssc;
  wire FpAdd_6U_10U_1_and_2_tmp;
  wire FpAdd_6U_10U_1_is_inf_3_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_9_m1c;
  wire FpAdd_6U_10U_1_and_16_ssc;
  wire FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_5_mx0w0;
  wire FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_4_mx0w0;
  wire FpAdd_6U_10U_1_and_30_ssc;
  wire FpAdd_6U_10U_1_and_1_tmp;
  wire FpAdd_6U_10U_1_is_inf_2_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_7_m1c;
  wire FpAdd_6U_10U_1_and_10_ssc;
  wire FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_5_mx0w0;
  wire FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_4_mx0w0;
  wire FpAdd_6U_10U_1_and_28_ssc;
  wire FpAdd_6U_10U_1_and_tmp;
  wire FpAdd_6U_10U_1_is_inf_1_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_1_and_4_ssc;
  wire [5:0] FpMul_6U_10U_p_expo_lpi_1_dfm_1_mx0;
  wire [5:0] FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_sva_1;
  wire [6:0] nl_FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_sva_1;
  wire inp_lookup_4_FpMantRNE_22U_11U_else_and_svs;
  wire FpMul_6U_10U_is_inf_lpi_1_dfm_2;
  wire FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp_3;
  wire [5:0] FpMul_6U_10U_p_expo_3_lpi_1_dfm_1_mx0;
  wire [5:0] FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_3_sva_1;
  wire [6:0] nl_FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_3_sva_1;
  wire inp_lookup_3_FpMantRNE_22U_11U_else_and_svs;
  wire FpMul_6U_10U_is_inf_3_lpi_1_dfm_2;
  wire FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp_2;
  wire [5:0] FpMul_6U_10U_p_expo_2_lpi_1_dfm_1_mx0;
  wire [5:0] FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_2_sva_1;
  wire [6:0] nl_FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_2_sva_1;
  wire inp_lookup_2_FpMantRNE_22U_11U_else_and_svs;
  wire FpMul_6U_10U_is_inf_2_lpi_1_dfm_2;
  wire FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp_1;
  wire [5:0] FpMul_6U_10U_p_expo_1_lpi_1_dfm_1_mx0;
  wire [5:0] FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_1_sva_1;
  wire [6:0] nl_FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_1_sva_1;
  wire inp_lookup_1_FpMantRNE_22U_11U_else_and_svs;
  wire FpMul_6U_10U_is_inf_1_lpi_1_dfm_2;
  wire FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp;
  wire inp_lookup_4_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_mx0w0;
  wire inp_lookup_4_IsZero_6U_10U_5_IsZero_6U_10U_5_nor_mx0w1;
  wire inp_lookup_3_IsZero_6U_10U_2_aif_IsZero_6U_10U_2_aelse_nor_2;
  wire inp_lookup_3_IsZero_6U_10U_5_IsZero_6U_10U_5_nor_2;
  wire inp_lookup_2_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_mx0w0;
  wire inp_lookup_2_IsZero_6U_10U_5_IsZero_6U_10U_5_nor_mx0w1;
  wire inp_lookup_1_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_2;
  wire inp_lookup_1_IsZero_6U_10U_5_IsZero_6U_10U_5_nor_2;
  wire FpMul_6U_10U_o_expo_lpi_1_dfm_3_5_mx0w0;
  wire FpMul_6U_10U_o_expo_lpi_1_dfm_3_4_mx0w0;
  wire FpMul_6U_10U_o_expo_3_lpi_1_dfm_3_5_mx0w0;
  wire FpMul_6U_10U_o_expo_3_lpi_1_dfm_3_4_mx0w0;
  wire FpMul_6U_10U_o_expo_2_lpi_1_dfm_3_5_mx0w0;
  wire FpMul_6U_10U_o_expo_2_lpi_1_dfm_3_4_mx0w0;
  wire FpMul_6U_10U_o_expo_1_lpi_1_dfm_3_5_mx0w0;
  wire FpMul_6U_10U_o_expo_1_lpi_1_dfm_3_4_mx0w0;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_3_cse;
  wire IsNaN_5U_10U_3_land_lpi_1_dfm;
  wire IsZero_5U_10U_3_land_lpi_1_dfm;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_3_cse;
  wire IsInf_5U_10U_1_land_lpi_1_dfm;
  wire IsNaN_5U_10U_1_land_lpi_1_dfm;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_2_cse;
  wire IsNaN_5U_10U_3_land_3_lpi_1_dfm;
  wire IsZero_5U_10U_3_land_3_lpi_1_dfm;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_2_cse;
  wire IsInf_5U_10U_1_land_3_lpi_1_dfm;
  wire IsNaN_5U_10U_1_land_3_lpi_1_dfm;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_1_cse;
  wire IsNaN_5U_10U_3_land_2_lpi_1_dfm;
  wire IsZero_5U_10U_3_land_2_lpi_1_dfm;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_1_cse;
  wire IsInf_5U_10U_1_land_2_lpi_1_dfm;
  wire IsNaN_5U_10U_1_land_2_lpi_1_dfm;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_cse;
  wire IsNaN_5U_10U_3_land_1_lpi_1_dfm;
  wire IsZero_5U_10U_3_land_1_lpi_1_dfm;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_cse;
  wire IsInf_5U_10U_1_land_1_lpi_1_dfm;
  wire IsNaN_5U_10U_1_land_1_lpi_1_dfm;
  wire FpMul_6U_10U_1_o_sign_lpi_1_dfm_mx0w0;
  wire FpMul_6U_10U_2_o_sign_lpi_1_dfm_mx0w0;
  wire FpMul_6U_10U_1_o_sign_3_lpi_1_dfm_mx0w0;
  wire FpMul_6U_10U_2_o_sign_3_lpi_1_dfm_mx0w0;
  wire FpMul_6U_10U_1_o_sign_2_lpi_1_dfm_mx0w0;
  wire FpMul_6U_10U_2_o_sign_2_lpi_1_dfm_mx0w0;
  wire FpMul_6U_10U_1_o_sign_1_lpi_1_dfm_mx0w0;
  wire FpMul_6U_10U_2_o_sign_1_lpi_1_dfm_mx0w0;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_nor_3_ssc;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_lpi_1_dfm_2;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_and_7_m1c;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_nor_2_ssc;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_3_lpi_1_dfm_2;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_and_5_m1c;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_nor_1_ssc;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_2_lpi_1_dfm_2;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_and_3_m1c;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_nor_ssc;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_1_lpi_1_dfm_2;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_and_1_m1c;
  wire IsDenorm_5U_10U_land_lpi_1_dfm;
  wire IsInf_5U_10U_land_lpi_1_dfm;
  wire IsInf_5U_10U_IsInf_5U_10U_and_cse_sva;
  wire IsDenorm_5U_10U_land_3_lpi_1_dfm;
  wire IsInf_5U_10U_land_3_lpi_1_dfm;
  wire IsInf_5U_10U_IsInf_5U_10U_and_cse_3_sva;
  wire IsDenorm_5U_10U_land_2_lpi_1_dfm;
  wire IsInf_5U_10U_land_2_lpi_1_dfm;
  wire IsInf_5U_10U_IsInf_5U_10U_and_cse_2_sva;
  wire IsDenorm_5U_10U_land_1_lpi_1_dfm;
  wire IsInf_5U_10U_land_1_lpi_1_dfm;
  wire IsInf_5U_10U_IsInf_5U_10U_and_cse_1_sva;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_3_0_mx0w0;
  wire IsDenorm_5U_10U_2_land_lpi_1_dfm;
  wire IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_sva;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_3_0_mx0w0;
  wire IsDenorm_5U_10U_2_land_3_lpi_1_dfm;
  wire IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_3_sva;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_3_0_mx0w0;
  wire IsDenorm_5U_10U_2_land_2_lpi_1_dfm;
  wire IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_2_sva;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_3_0_mx0w0;
  wire IsDenorm_5U_10U_2_land_1_lpi_1_dfm;
  wire IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_1_sva;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_3_cse;
  wire IsNaN_5U_10U_land_lpi_1_dfm;
  wire IsZero_5U_10U_land_lpi_1_dfm;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_2_cse;
  wire IsNaN_5U_10U_land_3_lpi_1_dfm;
  wire IsZero_5U_10U_land_3_lpi_1_dfm;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_1_cse;
  wire IsNaN_5U_10U_land_2_lpi_1_dfm;
  wire IsZero_5U_10U_land_2_lpi_1_dfm;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_cse;
  wire IsNaN_5U_10U_land_1_lpi_1_dfm;
  wire IsZero_5U_10U_land_1_lpi_1_dfm;
  wire FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_5;
  wire FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_4;
  wire FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_5;
  wire FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_4;
  wire FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_5;
  wire FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_4;
  wire FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_5;
  wire FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_4;
  wire [1:0] FpAdd_6U_10U_o_expo_lpi_1_dfm_2_5_4;
  wire [1:0] FpAdd_6U_10U_o_expo_3_lpi_1_dfm_2_5_4;
  wire [1:0] FpAdd_6U_10U_o_expo_2_lpi_1_dfm_2_5_4;
  wire [1:0] FpAdd_6U_10U_o_expo_1_lpi_1_dfm_2_5_4;
  wire FpFractionToFloat_35U_6U_10U_1_is_zero_lpi_1_dfm_1;
  wire FpFractionToFloat_35U_6U_10U_1_is_zero_3_lpi_1_dfm_1;
  wire FpFractionToFloat_35U_6U_10U_1_is_zero_2_lpi_1_dfm_1;
  wire FpFractionToFloat_35U_6U_10U_1_is_zero_1_lpi_1_dfm_1;
  wire inp_lookup_else_if_a0_15_10_lpi_1_dfm_3_5_mx0w1;
  wire inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_3_5_mx0w1;
  wire inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_3_5_mx0w1;
  wire inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_3_5_mx0w1;
  wire FpMul_6U_10U_1_o_expo_lpi_1_dfm_3_5_mx0w1;
  wire FpMul_6U_10U_1_o_expo_lpi_1_dfm_3_4_mx0w1;
  wire FpMul_6U_10U_1_lor_2_lpi_1_dfm;
  wire FpMul_6U_10U_1_and_6_ssc;
  wire [5:0] FpMul_6U_10U_1_o_expo_lpi_1_dfm;
  wire FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_5_mx1w1;
  wire FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_4_mx1w1;
  wire FpMul_6U_10U_1_lor_11_lpi_1_dfm;
  wire FpMul_6U_10U_1_and_4_ssc;
  wire [5:0] FpMul_6U_10U_1_o_expo_3_lpi_1_dfm;
  wire FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_3_5_mx1w1;
  wire FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_3_4_mx1w1;
  wire FpMul_6U_10U_1_lor_10_lpi_1_dfm;
  wire FpMul_6U_10U_1_and_2_ssc;
  wire [5:0] FpMul_6U_10U_1_o_expo_2_lpi_1_dfm;
  wire FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_3_5_mx1w1;
  wire FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_3_4_mx1w1;
  wire FpMul_6U_10U_1_lor_9_lpi_1_dfm;
  wire FpMul_6U_10U_1_and_ssc;
  wire [5:0] FpMul_6U_10U_1_o_expo_1_lpi_1_dfm;
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva;
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva;
  wire [5:0] FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_sva_3;
  wire [6:0] nl_FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_sva_3;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_sva;
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_3_sva;
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_3_sva;
  wire [5:0] FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_sva_3;
  wire [6:0] nl_FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_sva_3;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_3_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_3_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_3_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_3_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_3_sva;
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_2_sva;
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_2_sva;
  wire [5:0] FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_sva_3;
  wire [6:0] nl_FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_sva_3;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_2_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_2_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_2_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_2_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_2_sva;
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_1_sva;
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_1_sva;
  wire [5:0] FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_sva_3;
  wire [6:0] nl_FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_sva_3;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_1_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_1_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_1_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_1_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_1_sva;
  wire [19:0] FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0;
  wire [19:0] FpMul_6U_10U_p_mant_20_1_3_lpi_1_dfm_3_mx0;
  wire [19:0] FpMul_6U_10U_p_mant_20_1_2_lpi_1_dfm_3_mx0;
  wire [19:0] FpMul_6U_10U_p_mant_20_1_1_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_3_mx1;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_3_mx0w0;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_3_lpi_1_dfm_3_mx1;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_3_lpi_1_dfm_3_mx0w0;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_3_mx1;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_3_mx0w0;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_3_mx1;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_3_mx0w0;
  wire [5:0] FpMul_6U_10U_2_o_expo_lpi_1_dfm;
  wire [5:0] FpMul_6U_10U_2_o_expo_3_lpi_1_dfm;
  wire [5:0] FpMul_6U_10U_2_o_expo_2_lpi_1_dfm;
  wire [5:0] FpMul_6U_10U_2_o_expo_1_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_1_o_expo_lpi_1_dfm_7;
  wire [23:0] FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_mx0;
  wire [7:0] FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_7;
  wire [23:0] FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_mx0;
  wire [7:0] FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_7;
  wire [23:0] FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_mx0;
  wire [7:0] FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_7_mx0w0;
  wire [23:0] FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_mx0;
  wire [5:0] FpMul_6U_10U_o_expo_lpi_1_dfm;
  wire [5:0] FpMul_6U_10U_o_expo_3_lpi_1_dfm;
  wire [5:0] FpMul_6U_10U_o_expo_2_lpi_1_dfm;
  wire [5:0] FpMul_6U_10U_o_expo_1_lpi_1_dfm;
  wire [23:0] FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_mx0;
  wire [23:0] FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_mx0;
  wire [23:0] FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_mx0;
  wire [23:0] FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_mx0;
  wire [34:0] inp_lookup_else_if_a0_frac_sva_mx0w0;
  wire [35:0] nl_inp_lookup_else_if_a0_frac_sva_mx0w0;
  wire [34:0] inp_lookup_else_if_a0_frac_3_sva_mx0w0;
  wire [35:0] nl_inp_lookup_else_if_a0_frac_3_sva_mx0w0;
  wire [34:0] inp_lookup_else_if_a0_frac_2_sva_mx0w0;
  wire [35:0] nl_inp_lookup_else_if_a0_frac_2_sva_mx0w0;
  wire [34:0] inp_lookup_else_if_a0_frac_1_sva_mx0w0;
  wire [35:0] nl_inp_lookup_else_if_a0_frac_1_sva_mx0w0;
  wire FpAdd_8U_23U_else_6_mux_9_mx0w1;
  wire FpAdd_8U_23U_else_6_mux_6_mx0w1;
  wire FpAdd_8U_23U_else_6_mux_3_mx0w1;
  wire FpAdd_8U_23U_else_6_mux_mx0w1;
  wire [3:0] FpMul_6U_10U_o_expo_lpi_1_dfm_3_3_0_mx0w0;
  wire FpMul_6U_10U_lor_2_lpi_1_dfm;
  wire FpMul_6U_10U_and_6_ssc;
  wire [3:0] FpMul_6U_10U_o_expo_3_lpi_1_dfm_3_3_0_mx0w0;
  wire FpMul_6U_10U_lor_11_lpi_1_dfm;
  wire FpMul_6U_10U_and_4_ssc;
  wire [3:0] FpMul_6U_10U_o_expo_2_lpi_1_dfm_3_3_0_mx0w0;
  wire FpMul_6U_10U_lor_10_lpi_1_dfm;
  wire FpMul_6U_10U_and_2_ssc;
  wire [3:0] FpMul_6U_10U_o_expo_1_lpi_1_dfm_3_3_0_mx0w0;
  wire FpMul_6U_10U_lor_9_lpi_1_dfm;
  wire FpMul_6U_10U_and_ssc;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_sva;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_3_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_3_sva;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_2_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_2_sva;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_1_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_1_sva;
  wire FpMul_6U_10U_2_and_6_ssc;
  wire FpMul_6U_10U_2_and_4_ssc;
  wire FpMul_6U_10U_2_and_2_ssc;
  wire FpMul_6U_10U_2_and_ssc;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_sva;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_3_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_3_sva;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_2_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_2_sva;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_1_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_1_sva;
  wire [23:0] FpAdd_6U_10U_1_int_mant_p1_sva;
  wire [24:0] nl_FpAdd_6U_10U_1_int_mant_p1_sva;
  wire [23:0] FpAdd_6U_10U_1_int_mant_p1_3_sva;
  wire [24:0] nl_FpAdd_6U_10U_1_int_mant_p1_3_sva;
  wire [23:0] FpAdd_6U_10U_1_int_mant_p1_2_sva;
  wire [24:0] nl_FpAdd_6U_10U_1_int_mant_p1_2_sva;
  wire [23:0] FpAdd_6U_10U_1_int_mant_p1_1_sva;
  wire [24:0] nl_FpAdd_6U_10U_1_int_mant_p1_1_sva;
  wire [3:0] FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_3_0;
  wire [3:0] FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_3_0;
  wire [3:0] FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_3_0;
  wire [3:0] FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_3_0;
  wire [3:0] FpAdd_6U_10U_o_expo_lpi_1_dfm_2_3_0;
  wire [3:0] FpAdd_6U_10U_o_expo_3_lpi_1_dfm_2_3_0;
  wire [3:0] FpAdd_6U_10U_o_expo_2_lpi_1_dfm_2_3_0;
  wire [3:0] FpAdd_6U_10U_o_expo_1_lpi_1_dfm_2_3_0;
  wire [9:0] FpMul_6U_10U_1_o_mant_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpMul_6U_10U_1_o_expo_lpi_1_dfm_3_3_0_mx0w1;
  wire [9:0] FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_3_mx0w1;
  wire [3:0] FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_3_0_mx1w1;
  wire [9:0] FpMul_6U_10U_1_o_mant_2_lpi_1_dfm_3;
  wire [3:0] FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_3_3_0_mx1w1;
  wire [9:0] FpMul_6U_10U_1_o_mant_1_lpi_1_dfm_3;
  wire [3:0] FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_3_3_0_mx1w1;
  wire [9:0] FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_22_13_lpi_1_dfm_mx0w1;
  wire [9:0] FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_22_13_3_lpi_1_dfm_mx0w1;
  wire [9:0] FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_22_13_2_lpi_1_dfm_mx0w1;
  wire [9:0] FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_22_13_1_lpi_1_dfm_mx0w1;
  wire [1:0] FpAdd_6U_10U_o_expo_lpi_1_dfm_7_5_4;
  wire [1:0] FpAdd_6U_10U_o_expo_3_lpi_1_dfm_7_5_4;
  wire [1:0] FpAdd_6U_10U_o_expo_2_lpi_1_dfm_7_5_4;
  wire [1:0] FpAdd_6U_10U_o_expo_1_lpi_1_dfm_7_5_4;
  wire [22:0] FpAdd_8U_23U_1_o_mant_lpi_1_dfm_2_mx1;
  wire [22:0] FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx1;
  wire [22:0] FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_2_mx1;
  wire [22:0] FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_2_mx1;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_sva;
  wire IsZero_5U_10U_2_land_lpi_1_dfm;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_3_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_3_sva;
  wire IsZero_5U_10U_2_land_3_lpi_1_dfm;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_2_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_2_sva;
  wire IsZero_5U_10U_2_land_2_lpi_1_dfm;
  wire [4:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_1_sva;
  wire [5:0] nl_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_1_sva;
  wire IsZero_5U_10U_2_land_1_lpi_1_dfm;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_3_mx1;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_2_lpi_1_dfm_3_mx0;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_1_lpi_1_dfm_3_mx0;
  wire IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0;
  wire FpMul_6U_10U_1_FpMul_6U_10U_1_nor_2_ssc;
  wire FpMul_6U_10U_1_FpMul_6U_10U_1_nor_1_ssc;
  wire FpMul_6U_10U_1_FpMul_6U_10U_1_nor_ssc;
  wire FpMul_6U_10U_2_lor_2_lpi_1_dfm;
  wire FpMul_6U_10U_2_lor_11_lpi_1_dfm;
  wire FpMul_6U_10U_2_lor_10_lpi_1_dfm;
  wire FpMul_6U_10U_2_lor_9_lpi_1_dfm;
  wire [23:0] FpAdd_6U_10U_1_int_mant_p1_sva_1;
  wire [25:0] nl_FpAdd_6U_10U_1_int_mant_p1_sva_1;
  wire [23:0] FpAdd_6U_10U_1_int_mant_p1_3_sva_1;
  wire [25:0] nl_FpAdd_6U_10U_1_int_mant_p1_3_sva_1;
  wire [23:0] FpAdd_6U_10U_1_int_mant_p1_2_sva_1;
  wire [25:0] nl_FpAdd_6U_10U_1_int_mant_p1_2_sva_1;
  wire [23:0] FpAdd_6U_10U_1_int_mant_p1_1_sva_1;
  wire [25:0] nl_FpAdd_6U_10U_1_int_mant_p1_1_sva_1;
  wire FpMul_6U_10U_1_p_mant_p1_sva_mx2_21;
  wire FpMul_6U_10U_1_p_mant_p1_3_sva_mx2_21;
  wire FpMul_6U_10U_1_p_mant_p1_2_sva_mx2_21;
  wire FpMul_6U_10U_1_p_mant_p1_1_sva_mx2_21;
  wire FpMul_6U_10U_2_p_mant_p1_sva_mx2_21;
  wire FpMul_6U_10U_2_p_mant_p1_3_sva_mx2_21;
  wire FpMul_6U_10U_2_p_mant_p1_2_sva_mx2_21;
  wire FpMul_6U_10U_2_p_mant_p1_1_sva_mx2_21;
  wire FpMul_6U_10U_FpMul_6U_10U_nor_3_ssc;
  wire FpMul_6U_10U_FpMul_6U_10U_nor_2_ssc;
  wire FpMul_6U_10U_FpMul_6U_10U_nor_1_ssc;
  wire FpMul_6U_10U_FpMul_6U_10U_nor_ssc;
  wire [32:0] inp_lookup_if_else_o_acc_psp_sva;
  wire [33:0] nl_inp_lookup_if_else_o_acc_psp_sva;
  wire [32:0] inp_lookup_if_else_o_acc_psp_3_sva;
  wire [33:0] nl_inp_lookup_if_else_o_acc_psp_3_sva;
  wire [32:0] inp_lookup_if_else_o_acc_psp_2_sva;
  wire [33:0] nl_inp_lookup_if_else_o_acc_psp_2_sva;
  wire [32:0] inp_lookup_if_else_o_acc_psp_1_sva;
  wire [33:0] nl_inp_lookup_if_else_o_acc_psp_1_sva;
  wire [3:0] FpAdd_6U_10U_o_expo_lpi_1_dfm_7_3_0;
  wire [3:0] FpAdd_6U_10U_o_expo_3_lpi_1_dfm_7_3_0;
  wire [3:0] FpAdd_6U_10U_o_expo_2_lpi_1_dfm_7_3_0;
  wire [3:0] FpAdd_6U_10U_o_expo_1_lpi_1_dfm_7_3_0;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_3_mx0w0;
  wire [3:0] FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_3_0_mx0w0;
  wire [3:0] FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_3_0_mx0w0;
  wire [3:0] FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_3_0_mx0w0;
  wire [3:0] FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_3_0_mx0w0;
  wire [4:0] FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_3_4_0_mx0w0;
  wire [4:0] FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_3_4_0_mx0w0;
  wire [4:0] FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_3_4_0_mx0w0;
  wire [4:0] FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_3_4_0_mx0w0;
  wire [4:0] inp_lookup_else_if_a0_15_10_lpi_1_dfm_3_4_0_mx0w0;
  wire [4:0] inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_3_4_0_mx0w0;
  wire [4:0] inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_3_4_0_mx0w0;
  wire [4:0] inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_3_4_0_mx0w0;
  wire [9:0] FpFractionToFloat_35U_6U_10U_1_o_mant_lpi_1_dfm_3_mx0w0;
  wire [9:0] FpFractionToFloat_35U_6U_10U_1_o_mant_3_lpi_1_dfm_3_mx0w0;
  wire [9:0] FpFractionToFloat_35U_6U_10U_1_o_mant_2_lpi_1_dfm_3_mx0w0;
  wire [9:0] FpFractionToFloat_35U_6U_10U_1_o_mant_1_lpi_1_dfm_3_mx0w0;
  wire [9:0] inp_lookup_else_if_a0_9_0_lpi_1_dfm_3_mx0w0;
  wire [9:0] inp_lookup_else_if_a0_9_0_3_lpi_1_dfm_3_mx0w0;
  wire [9:0] inp_lookup_else_if_a0_9_0_2_lpi_1_dfm_3_mx0w0;
  wire [9:0] inp_lookup_else_if_a0_9_0_1_lpi_1_dfm_3_mx0w0;
  wire [9:0] FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_9_0_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_9_0_3_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_9_0_2_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_9_0_1_lpi_1_dfm;
  wire [9:0] FpMul_6U_10U_o_mant_lpi_1_dfm_3_mx0w0;
  wire [9:0] FpMul_6U_10U_o_mant_3_lpi_1_dfm_3_mx0w0;
  wire [9:0] FpMul_6U_10U_o_mant_2_lpi_1_dfm_3_mx0w0;
  wire [9:0] FpMul_6U_10U_o_mant_1_lpi_1_dfm_3_mx0w0;
  wire [9:0] FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_22_13_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_22_13_3_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_22_13_2_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_22_13_1_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_9_0_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_9_0_3_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_9_0_2_lpi_1_dfm;
  wire [9:0] FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_9_0_1_lpi_1_dfm;
  wire [66:0] IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_sva;
  wire [67:0] nl_IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_sva;
  wire [66:0] IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_3_sva;
  wire [67:0] nl_IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_3_sva;
  wire [66:0] IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_2_sva;
  wire [67:0] nl_IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_2_sva;
  wire [66:0] IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_1_sva;
  wire [67:0] nl_IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_1_sva;
  wire IntShiftRight_69U_6U_32U_obits_fixed_and_m1c;
  wire IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_1;
  wire IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_2;
  wire IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_3;
  wire IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_4;
  wire IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_5;
  wire and_2321_m1c;
  wire IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_6;
  wire IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_7;
  wire and_2319_m1c;
  wire and_m1c;
  wire and_2315_m1c;
  wire and_m1c_1;
  wire and_2311_m1c;
  wire and_m1c_2;
  wire and_2307_m1c;
  wire and_m1c_3;
  wire inp_lookup_if_and_m1c;
  wire inp_lookup_if_and_m1c_1;
  wire inp_lookup_if_and_m1c_2;
  wire and_1944_m1c;
  wire inp_lookup_if_and_m1c_3;
  wire inp_lookup_if_and_m1c_4;
  wire inp_lookup_if_and_m1c_5;
  wire and_1942_m1c;
  wire inp_lookup_if_and_m1c_6;
  wire inp_lookup_if_and_m1c_7;
  wire inp_lookup_if_and_m1c_8;
  wire inp_lookup_if_and_m1c_9;
  wire inp_lookup_if_and_m1c_10;
  wire inp_lookup_if_and_m1c_11;
  reg [9:0] reg_FpMantRNE_36U_11U_1_else_ac_int_cctor_tmp;
  reg [9:0] reg_FpMantRNE_36U_11U_1_else_ac_int_cctor_4_tmp;
  reg [9:0] reg_FpMantRNE_36U_11U_1_else_ac_int_cctor_3_tmp;
  reg [9:0] reg_FpMantRNE_36U_11U_1_else_ac_int_cctor_2_tmp;
  wire or_4591_tmp;
  wire chn_inp_out_and_cse;
  wire or_11_cse;
  wire or_82_cse;
  wire nor_1713_cse;
  wire or_356_cse;
  wire FpAdd_8U_23U_o_expo_and_cse;
  wire or_461_cse;
  wire or_683_cse;
  wire or_471_cse;
  wire or_523_cse;
  wire or_740_cse;
  wire or_597_cse;
  wire or_792_cse;
  wire or_801_cse;
  wire or_802_cse;
  wire mux_500_cse;
  wire nor_1584_cse;
  wire nor_126_cse;
  wire nor_136_cse;
  wire nor_1546_cse;
  wire nor_1517_cse;
  wire IsInf_6U_23U_aelse_and_cse;
  wire IsInf_6U_23U_aelse_and_1_cse;
  wire IsInf_6U_23U_aelse_and_2_cse;
  wire IsInf_6U_23U_aelse_and_3_cse;
  reg reg_chn_inp_out_rsci_ld_core_psct_cse;
  wire nor_44_cse;
  wire nor_67_cse;
  wire IntLeadZero_35U_1_leading_sign_35_0_rtn_and_cse;
  wire IntLeadZero_35U_1_leading_sign_35_0_rtn_and_1_cse;
  wire IntLeadZero_35U_1_leading_sign_35_0_rtn_and_2_cse;
  wire IntLeadZero_35U_1_leading_sign_35_0_rtn_and_3_cse;
  wire nor_1340_cse;
  wire and_3358_cse;
  wire and_3355_cse;
  wire and_3351_cse;
  wire and_3345_cse;
  wire and_3393_cse;
  wire and_3246_cse;
  wire and_3391_cse;
  wire and_3244_cse;
  wire and_3401_cse;
  wire and_3242_cse;
  wire nor_35_cse;
  wire or_507_cse;
  wire nor_1264_cse;
  wire nor_55_cse;
  wire nor_1251_cse;
  wire and_3240_cse;
  wire mux_1015_cse;
  wire mux_1031_cse;
  wire nand_661_cse;
  wire nand_579_cse;
  wire mux_476_cse;
  wire mux_485_cse;
  wire FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_1_cse;
  wire FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_2_cse;
  wire nor_1397_cse;
  wire nor_1407_cse;
  wire FpAdd_6U_10U_and_35_cse;
  wire FpAdd_6U_10U_and_37_cse;
  wire FpAdd_6U_10U_and_39_cse;
  wire and_3389_cse;
  wire and_3249_cse;
  wire nor_268_cse;
  wire nor_267_cse;
  wire or_763_cse;
  wire or_3291_cse;
  wire mux_1061_cse;
  wire or_3384_cse;
  wire or_3379_cse;
  wire nor_956_cse;
  wire or_3484_cse;
  wire or_3489_cse;
  wire FpAdd_6U_10U_and_41_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_3_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_6_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_9_cse;
  wire nor_1593_cse;
  wire nor_1587_cse;
  wire mux_1140_cse;
  wire nor_1130_cse;
  wire nor_1210_cse;
  wire nor_1221_cse;
  wire nor_1193_cse;
  wire or_5689_cse;
  wire and_2320_cse;
  wire nor_1217_cse;
  wire nor_905_cse;
  wire nor_908_cse;
  wire nor_898_cse;
  wire nor_901_cse;
  wire nor_605_cse;
  wire nor_894_cse;
  wire or_3722_cse;
  wire or_3720_cse;
  wire or_3718_cse;
  wire or_3716_cse;
  wire FpAdd_8U_23U_o_sign_and_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_3_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_6_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_9_cse;
  wire and_3149_cse;
  wire or_79_cse;
  wire or_457_cse;
  wire or_519_cse;
  wire FpAdd_8U_23U_or_2_cse;
  wire or_593_cse;
  wire or_648_cse;
  wire FpAdd_6U_10U_1_or_12_cse;
  wire FpAdd_6U_10U_1_or_16_cse;
  wire FpAdd_6U_10U_1_or_18_cse;
  wire or_5020_cse;
  wire or_5021_cse;
  wire or_5022_cse;
  wire or_5023_cse;
  wire FpAdd_8U_23U_or_cse;
  wire FpAdd_8U_23U_or_1_cse;
  wire FpAdd_8U_23U_or_3_cse;
  wire nor_1225_cse;
  wire nor_1208_cse;
  wire nor_1191_cse;
  wire nor_1180_cse;
  wire nor_1727_cse;
  wire FpAdd_6U_10U_or_16_cse;
  wire FpAdd_6U_10U_or_17_cse;
  wire FpAdd_6U_10U_or_18_cse;
  wire FpAdd_6U_10U_or_19_cse;
  wire nor_1274_cse;
  wire or_3779_cse;
  wire nor_1238_cse;
  wire nand_694_cse;
  wire or_2176_cse;
  wire nor_1380_cse;
  wire nand_358_cse;
  wire nand_693_cse;
  wire nor_1354_cse;
  wire nor_301_cse;
  wire nand_616_cse;
  wire nor_29_cse;
  wire or_5372_cse;
  wire and_348_cse;
  wire nor_275_cse;
  wire or_604_cse;
  wire or_2282_cse;
  wire or_2010_cse;
  wire nor_572_cse;
  wire or_3850_cse;
  wire or_3167_cse;
  wire or_2663_cse;
  wire or_2797_cse;
  wire and_3374_cse;
  wire or_2810_cse;
  wire or_2822_cse;
  wire nand_653_cse;
  wire nand_652_cse;
  wire nor_884_cse;
  wire or_5369_cse;
  wire nor_257_cse;
  wire nor_880_cse;
  wire or_504_cse;
  wire nor_584_cse;
  wire nor_266_cse;
  wire nor_875_cse;
  wire nor_586_cse;
  wire or_114_cse;
  wire nor_5_cse;
  wire or_178_cse;
  wire nor_13_cse;
  wire nor_74_cse;
  wire or_2444_cse;
  wire or_2445_cse;
  wire nand_570_cse;
  wire and_3113_cse;
  wire and_3111_cse;
  wire and_3110_cse;
  wire and_3112_cse;
  wire nor_1371_cse;
  wire or_3558_cse;
  wire and_3118_cse;
  wire and_3120_cse;
  wire and_3124_cse;
  wire and_3106_cse;
  wire or_3885_cse;
  wire or_3913_cse;
  wire or_3941_cse;
  wire or_3969_cse;
  wire or_2_cse;
  wire and_3056_cse;
  wire nor_1017_cse;
  wire and_3054_cse;
  wire and_3346_cse;
  wire nand_544_cse;
  wire nand_557_cse;
  wire FpAdd_6U_10U_1_is_a_greater_oelse_FpAdd_6U_10U_1_is_a_greater_oelse_and_cse;
  wire FpAdd_6U_10U_1_is_a_greater_oelse_FpAdd_6U_10U_1_is_a_greater_oelse_and_1_cse;
  wire FpAdd_6U_10U_1_is_a_greater_oelse_FpAdd_6U_10U_1_is_a_greater_oelse_and_2_cse;
  wire or_1970_cse;
  wire [30:0] mux_1993_rgt;
  wire [9:0] FpMul_6U_10U_2_o_mant_FpMul_6U_10U_2_o_mant_mux_rgt;
  wire [7:0] FpAdd_8U_23U_o_expo_FpAdd_8U_23U_o_expo_mux_rgt;
  wire [7:0] FpAdd_8U_23U_o_expo_FpAdd_8U_23U_o_expo_mux_1_rgt;
  wire [7:0] FpAdd_8U_23U_o_expo_FpAdd_8U_23U_o_expo_mux_2_rgt;
  wire [7:0] FpAdd_8U_23U_o_expo_FpAdd_8U_23U_o_expo_mux_3_rgt;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_mux1h_11_rgt;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_mux1h_16_rgt;
  wire [35:0] inp_lookup_else_else_a0_mux1h_rgt;
  wire [35:0] inp_lookup_else_else_a0_mux1h_1_rgt;
  wire [35:0] inp_lookup_else_else_a0_mux1h_2_rgt;
  wire [35:0] inp_lookup_else_else_a0_mux1h_3_rgt;
  reg [7:0] reg_chn_inp_in_crt_sva_3_510_480_reg;
  reg [22:0] reg_chn_inp_in_crt_sva_3_510_480_1_reg;
  reg [7:0] reg_chn_inp_in_crt_sva_3_542_512_reg;
  reg [22:0] reg_chn_inp_in_crt_sva_3_542_512_1_reg;
  reg [7:0] reg_chn_inp_in_crt_sva_3_574_544_reg;
  reg [22:0] reg_chn_inp_in_crt_sva_3_574_544_1_reg;
  reg [7:0] reg_chn_inp_in_crt_sva_3_606_576_reg;
  reg [22:0] reg_chn_inp_in_crt_sva_3_606_576_1_reg;
  reg [1:0] reg_FpMul_6U_10U_2_o_mant_lpi_1_dfm_7_reg;
  reg [7:0] reg_FpMul_6U_10U_2_o_mant_lpi_1_dfm_7_1_reg;
  reg [7:0] reg_chn_inp_in_crt_sva_6_30_0_reg;
  reg [22:0] reg_chn_inp_in_crt_sva_6_30_0_1_reg;
  reg [7:0] reg_chn_inp_in_crt_sva_6_62_32_reg;
  reg [22:0] reg_chn_inp_in_crt_sva_6_62_32_1_reg;
  reg [7:0] reg_chn_inp_in_crt_sva_6_94_64_reg;
  reg [22:0] reg_chn_inp_in_crt_sva_6_94_64_1_reg;
  reg [7:0] reg_chn_inp_in_crt_sva_6_126_96_reg;
  reg [22:0] reg_chn_inp_in_crt_sva_6_126_96_1_reg;
  reg [1:0] reg_FpAdd_8U_23U_o_expo_1_lpi_1_dfm_11_reg;
  reg [5:0] reg_FpAdd_8U_23U_o_expo_1_lpi_1_dfm_11_1_reg;
  reg [1:0] reg_FpAdd_8U_23U_o_expo_2_lpi_1_dfm_11_reg;
  reg [5:0] reg_FpAdd_8U_23U_o_expo_2_lpi_1_dfm_11_1_reg;
  reg [1:0] reg_FpAdd_8U_23U_o_expo_3_lpi_1_dfm_11_reg;
  reg [5:0] reg_FpAdd_8U_23U_o_expo_3_lpi_1_dfm_11_1_reg;
  reg [1:0] reg_FpAdd_8U_23U_o_expo_lpi_1_dfm_11_reg;
  reg [5:0] reg_FpAdd_8U_23U_o_expo_lpi_1_dfm_11_1_reg;
  reg [3:0] reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_8_reg;
  reg [5:0] reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_8_1_reg;
  reg [3:0] reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_8_reg;
  reg [5:0] reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_8_1_reg;
  reg reg_inp_lookup_1_else_else_a0_acc_reg;
  reg reg_inp_lookup_1_else_else_a0_acc_1_reg;
  reg [33:0] reg_inp_lookup_1_else_else_a0_acc_2_reg;
  reg reg_inp_lookup_2_else_else_a0_acc_reg;
  reg reg_inp_lookup_2_else_else_a0_acc_1_reg;
  reg [33:0] reg_inp_lookup_2_else_else_a0_acc_2_reg;
  reg reg_inp_lookup_3_else_else_a0_acc_reg;
  reg reg_inp_lookup_3_else_else_a0_acc_1_reg;
  reg [33:0] reg_inp_lookup_3_else_else_a0_acc_2_reg;
  reg reg_inp_lookup_4_else_else_a0_acc_reg;
  reg reg_inp_lookup_4_else_else_a0_acc_1_reg;
  reg [33:0] reg_inp_lookup_4_else_else_a0_acc_2_reg;
  wire FpAdd_6U_10U_1_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0;
  wire [48:0] FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0;
  wire [48:0] FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0;
  wire [48:0] FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_1_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0;
  wire FpAdd_6U_10U_1_is_a_greater_lor_lpi_1_dfm_1_mx0w0;
  wire [48:0] FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0;
  wire [5:0] FpMul_6U_10U_1_else_2_else_ac_int_cctor_1_sva_mx0w0;
  wire [6:0] nl_FpMul_6U_10U_1_else_2_else_ac_int_cctor_1_sva_mx0w0;
  wire [5:0] FpMul_6U_10U_1_else_2_else_ac_int_cctor_2_sva_mx0w0;
  wire [6:0] nl_FpMul_6U_10U_1_else_2_else_ac_int_cctor_2_sva_mx0w0;
  wire [5:0] FpMul_6U_10U_1_else_2_else_ac_int_cctor_3_sva_mx0w0;
  wire [6:0] nl_FpMul_6U_10U_1_else_2_else_ac_int_cctor_3_sva_mx0w0;
  wire [5:0] FpMul_6U_10U_1_else_2_else_ac_int_cctor_sva_mx0w0;
  wire [6:0] nl_FpMul_6U_10U_1_else_2_else_ac_int_cctor_sva_mx0w0;
  wire [5:0] FpMul_6U_10U_2_else_2_else_ac_int_cctor_1_sva_mx0w0;
  wire [6:0] nl_FpMul_6U_10U_2_else_2_else_ac_int_cctor_1_sva_mx0w0;
  wire [5:0] FpMul_6U_10U_2_else_2_else_ac_int_cctor_sva_mx0w0;
  wire [6:0] nl_FpMul_6U_10U_2_else_2_else_ac_int_cctor_sva_mx0w0;
  wire and_3463_cse;
  wire or_5800_cse;
  wire mux_400_cse;
  wire nor_1800_cse;
  wire or_5809_cse;
  wire nor_1113_cse;
  wire nor_959_cse;
  wire nor_960_cse;
  wire mux_1480_cse;
  wire nor_950_cse;
  wire nor_952_cse;
  wire mux_1493_cse;
  wire nor_941_cse;
  wire nor_943_cse;
  wire mux_1506_cse;
  wire nor_1124_cse;
  wire nor_932_cse;
  wire mux_1519_cse;
  wire nor_1798_cse;
  wire or_5680_cse;
  wire nor_1224_cse;
  wire nor_1207_cse;
  wire nor_1190_cse;
  wire nor_1273_cse;
  wire nor_1790_cse;
  wire nor_1789_cse;
  wire nor_1237_cse;
  wire nand_701_cse;
  wire and_3483_cse;
  wire [10:0] FpMantRNE_36U_11U_1_else_ac_int_cctor_2_sva_mx0w0;
  wire [11:0] nl_FpMantRNE_36U_11U_1_else_ac_int_cctor_2_sva_mx0w0;
  wire [10:0] FpMantRNE_36U_11U_1_else_ac_int_cctor_3_sva_mx0w0;
  wire [11:0] nl_FpMantRNE_36U_11U_1_else_ac_int_cctor_3_sva_mx0w0;
  wire [10:0] FpMantRNE_36U_11U_1_else_ac_int_cctor_4_sva_mx0w0;
  wire [11:0] nl_FpMantRNE_36U_11U_1_else_ac_int_cctor_4_sva_mx0w0;
  wire [10:0] FpMantRNE_36U_11U_1_else_ac_int_cctor_sva_mx0w0;
  wire [11:0] nl_FpMantRNE_36U_11U_1_else_ac_int_cctor_sva_mx0w0;
  wire [19:0] FpMul_6U_10U_1_p_mant_20_1_3_lpi_1_dfm_3_mx0;
  wire [19:0] FpMul_6U_10U_1_p_mant_20_1_1_lpi_1_dfm_3_mx0;
  wire [19:0] FpMul_6U_10U_1_p_mant_20_1_lpi_1_dfm_3_mx0;
  wire inp_lookup_asn_106;
  wire inp_lookup_and_8_m1c;
  wire IsInf_6U_23U_land_1_lpi_1_dfm_mx0w0;
  wire IsNaN_6U_23U_land_1_lpi_1_dfm_mx2;
  wire inp_lookup_and_10_m1c;
  wire inp_lookup_asn_122;
  wire inp_lookup_and_28_m1c;
  wire IsInf_6U_23U_land_2_lpi_1_dfm_mx0w0;
  wire IsNaN_6U_23U_land_2_lpi_1_dfm_mx2;
  wire inp_lookup_and_30_m1c;
  wire inp_lookup_asn_114;
  wire inp_lookup_and_48_m1c;
  wire IsInf_6U_23U_land_3_lpi_1_dfm_mx0w0;
  wire IsNaN_6U_23U_land_3_lpi_1_dfm_mx1;
  wire inp_lookup_and_50_m1c;
  wire inp_lookup_asn_98;
  wire inp_lookup_and_68_m1c;
  wire IsInf_6U_23U_land_lpi_1_dfm_mx0w0;
  wire IsNaN_6U_23U_land_lpi_1_dfm_mx1;
  wire inp_lookup_and_70_m1c;
  wire IsInf_6U_23U_1_land_lpi_1_dfm_mx0w0;
  wire IsInf_6U_23U_1_land_3_lpi_1_dfm_mx0w0;
  wire IsInf_6U_23U_1_land_2_lpi_1_dfm_mx0w0;
  wire IsInf_6U_23U_1_land_1_lpi_1_dfm_mx0w0;
  wire [9:0] FpExpoWidthInc_6U_8U_23U_0U_1U_o_mant_9_0_1_lpi_1_dfm_2_mx0;
  wire inp_lookup_asn_110;
  wire [9:0] FpExpoWidthInc_6U_8U_23U_0U_1U_o_mant_9_0_2_lpi_1_dfm_2_mx0;
  wire inp_lookup_asn_126;
  wire [9:0] FpExpoWidthInc_6U_8U_23U_0U_1U_o_mant_9_0_3_lpi_1_dfm_2_mx0;
  wire inp_lookup_asn_118;
  wire [9:0] FpExpoWidthInc_6U_8U_23U_0U_1U_o_mant_9_0_lpi_1_dfm_2_mx0;
  wire inp_lookup_asn_102;
  wire and_3548_tmp;
  wire or_5842_tmp;
  wire and_3547_tmp;
  wire or_5840_tmp;
  wire and_3546_tmp;
  wire or_5838_tmp;
  wire and_3545_tmp;
  wire or_5836_tmp;
  wire and_3588_cse;
  wire and_3587_cse;
  wire and_3586_cse;
  wire and_3585_cse;
  wire and_861_rgt;
  wire IsZero_6U_10U_6_IsZero_6U_10U_6_nor_tmp;
  wire not_tmp_2674;
  wire or_tmp_4611;
  wire or_tmp_4615;
  wire or_tmp_4620;
  wire and_869_rgt;
  wire IsZero_6U_10U_6_IsZero_6U_10U_6_nor_1_tmp;
  wire nor_tmp_708;
  wire or_tmp_4625;
  wire and_877_rgt;
  wire and_883_rgt;
  wire IsZero_6U_10U_6_IsZero_6U_10U_6_nor_3_tmp;
  wire or_tmp_4637;
  wire and_899_rgt;
  wire and_901_rgt;
  wire and_903_rgt;
  wire and_907_rgt;
  wire and_912_rgt;
  wire and_915_rgt;
  wire and_918_rgt;
  wire and_920_rgt;
  wire and_936_rgt;
  wire and_939_rgt;
  wire and_941_rgt;
  wire and_945_rgt;
  wire and_950_rgt;
  wire and_953_rgt;
  wire and_956_rgt;
  wire and_973_rgt;
  wire and_976_rgt;
  wire and_978_rgt;
  wire and_982_rgt;
  wire and_987_rgt;
  wire and_990_rgt;
  wire and_993_rgt;
  wire nor_1743_rgt;
  wire and_1012_rgt;
  wire and_1014_rgt;
  wire and_1018_rgt;
  wire and_1023_rgt;
  wire and_1026_rgt;
  wire and_1029_rgt;
  wire and_1049_rgt;
  wire and_1052_rgt;
  wire and_1068_rgt;
  wire and_1071_rgt;
  wire and_1099_rgt;
  wire and_1102_rgt;
  wire and_1131_rgt;
  wire and_dcpl_2185;
  wire or_tmp_4675;
  wire and_1139_rgt;
  wire or_tmp_4685;
  wire and_1147_rgt;
  wire or_tmp_4698;
  wire or_tmp_4703;
  wire and_1155_rgt;
  wire and_1163_rgt;
  wire and_1174_rgt;
  wire and_1192_rgt;
  wire and_1209_rgt;
  wire and_1211_rgt;
  wire and_1213_rgt;
  wire FpAdd_6U_10U_1_and_47_rgt;
  wire and_1217_rgt;
  wire and_1221_rgt;
  wire and_1223_rgt;
  wire and_1225_rgt;
  wire and_1229_rgt;
  wire and_1233_rgt;
  wire and_1235_rgt;
  wire and_1237_rgt;
  wire and_1241_rgt;
  wire and_1245_rgt;
  wire and_1247_rgt;
  wire and_1249_rgt;
  wire and_1253_rgt;
  wire and_1270_rgt;
  wire and_1273_rgt;
  wire and_1277_rgt;
  wire and_1279_rgt;
  wire and_1280_rgt;
  wire and_1293_rgt;
  wire and_1296_rgt;
  wire nor_1733_rgt;
  wire and_1303_rgt;
  wire and_1304_rgt;
  wire and_1317_rgt;
  wire and_1320_rgt;
  wire nor_1732_rgt;
  wire and_1327_rgt;
  wire and_1329_rgt;
  wire and_1342_rgt;
  wire and_1345_rgt;
  wire and_1349_rgt;
  wire and_1351_rgt;
  wire and_1352_rgt;
  wire and_1360_rgt;
  wire and_1364_rgt;
  wire and_1368_rgt;
  wire and_1372_rgt;
  wire and_1386_rgt;
  wire and_1388_rgt;
  wire and_1390_rgt;
  wire and_1392_rgt;
  wire and_dcpl_2279;
  wire and_1468_rgt;
  wire and_1471_rgt;
  wire and_1474_rgt;
  wire and_1477_rgt;
  wire and_1537_rgt;
  wire and_1538_rgt;
  wire and_1588_rgt;
  wire and_1589_rgt;
  wire and_1639_rgt;
  wire and_1640_rgt;
  wire and_1690_rgt;
  wire and_1691_rgt;
  wire and_dcpl_2318;
  wire or_tmp_4714;
  wire or_tmp_4721;
  wire or_tmp_4726;
  wire or_tmp_4730;
  wire and_1717_rgt;
  wire and_1725_rgt;
  wire and_1726_rgt;
  wire and_1734_rgt;
  wire and_1735_rgt;
  wire and_1743_rgt;
  wire and_1744_rgt;
  wire and_1752_rgt;
  wire and_1754_rgt;
  wire and_1755_rgt;
  wire and_1757_rgt;
  wire and_1758_rgt;
  wire and_1760_rgt;
  wire and_1761_rgt;
  wire and_1764_rgt;
  wire and_1768_rgt;
  wire and_1772_rgt;
  wire and_1776_rgt;
  wire and_1780_rgt;
  wire and_1794_rgt;
  wire and_1796_rgt;
  wire and_1798_rgt;
  wire and_1800_rgt;
  wire and_1802_rgt;
  wire and_1804_rgt;
  wire and_1806_rgt;
  wire and_1808_rgt;
  wire and_1816_rgt;
  wire and_1821_rgt;
  wire and_1829_rgt;
  wire and_1834_rgt;
  wire and_1842_rgt;
  wire and_1847_rgt;
  wire and_1855_rgt;
  wire and_1860_rgt;
  wire or_tmp_4737;
  wire or_tmp_4741;
  wire or_tmp_4745;
  wire or_tmp_4753;
  wire and_1871_rgt;
  wire and_1873_rgt;
  wire and_1875_rgt;
  wire and_1877_rgt;
  wire and_1881_rgt;
  wire nor_1765_rgt;
  wire and_1888_rgt;
  wire and_1892_rgt;
  wire nor_1764_rgt;
  wire and_1899_rgt;
  wire and_1903_rgt;
  wire nor_1763_rgt;
  wire and_1910_rgt;
  wire and_1914_rgt;
  wire nor_1762_rgt;
  wire and_1921_rgt;
  wire and_dcpl_2461;
  wire inp_lookup_if_or_6_rgt;
  wire inp_lookup_if_or_7_rgt;
  wire inp_lookup_if_and_31_rgt;
  wire and_1941_rgt;
  wire inp_lookup_if_or_4_rgt;
  wire inp_lookup_if_or_5_rgt;
  wire inp_lookup_if_and_23_rgt;
  wire and_1943_rgt;
  wire inp_lookup_if_or_2_rgt;
  wire inp_lookup_if_or_3_rgt;
  wire inp_lookup_if_and_15_rgt;
  wire and_1945_rgt;
  wire inp_lookup_if_or_rgt;
  wire inp_lookup_if_or_1_rgt;
  wire inp_lookup_if_and_7_rgt;
  wire and_1947_rgt;
  wire and_1975_rgt;
  wire and_1978_rgt;
  wire and_1982_rgt;
  wire and_1985_rgt;
  wire and_2012_rgt;
  wire and_2013_rgt;
  wire and_2022_rgt;
  wire and_2023_rgt;
  wire and_2033_rgt;
  wire and_2034_rgt;
  wire and_2043_rgt;
  wire and_2044_rgt;
  wire and_2054_rgt;
  wire and_2065_rgt;
  wire and_2067_rgt;
  wire and_2069_rgt;
  wire and_2073_rgt;
  wire and_2076_rgt;
  wire and_2078_rgt;
  wire and_2097_rgt;
  wire and_2104_rgt;
  wire and_dcpl_2487;
  wire and_2112_rgt;
  wire and_2119_rgt;
  wire and_dcpl_2500;
  wire and_2125_rgt;
  wire and_2130_rgt;
  wire and_2135_rgt;
  wire and_2140_rgt;
  wire and_dcpl_2528;
  wire and_2194_rgt;
  wire and_2284_rgt;
  wire and_2287_rgt;
  wire and_2289_rgt;
  wire and_2291_rgt;
  wire and_2294_rgt;
  wire and_2296_rgt;
  wire and_2298_rgt;
  wire and_2301_rgt;
  wire and_2303_rgt;
  wire or_5766_rgt;
  wire or_5767_rgt;
  wire or_5764_rgt;
  wire or_5765_rgt;
  wire or_5762_rgt;
  wire or_5763_rgt;
  wire or_5760_rgt;
  wire or_5761_rgt;
  wire IntShiftRight_69U_6U_32U_obits_fixed_or_6_rgt;
  wire IntShiftRight_69U_6U_32U_obits_fixed_or_7_rgt;
  wire IntShiftRight_69U_6U_32U_obits_fixed_or_4_rgt;
  wire IntShiftRight_69U_6U_32U_obits_fixed_or_5_rgt;
  wire IntShiftRight_69U_6U_32U_obits_fixed_or_2_rgt;
  wire IntShiftRight_69U_6U_32U_obits_fixed_or_3_rgt;
  wire IntShiftRight_69U_6U_32U_obits_fixed_or_rgt;
  wire IntShiftRight_69U_6U_32U_obits_fixed_or_1_rgt;
  wire and_2342_rgt;
  wire and_2345_rgt;
  wire and_2348_rgt;
  wire and_2350_rgt;
  wire and_2351_rgt;
  wire and_2358_rgt;
  wire and_2359_rgt;
  wire and_2367_rgt;
  wire and_2368_rgt;
  wire and_2375_rgt;
  wire and_2376_rgt;
  wire and_2384_rgt;
  wire and_2385_rgt;
  wire IntSaturation_51U_32U_o_IntSaturation_51U_32U_o_nor_rgt;
  wire IntSaturation_51U_32U_and_7_rgt;
  wire IntSaturation_51U_32U_o_and_7_rgt;
  wire IntSaturation_51U_32U_o_IntSaturation_51U_32U_o_nor_1_rgt;
  wire IntSaturation_51U_32U_and_5_rgt;
  wire IntSaturation_51U_32U_o_and_5_rgt;
  wire IntSaturation_51U_32U_o_IntSaturation_51U_32U_o_nor_2_rgt;
  wire IntSaturation_51U_32U_and_3_rgt;
  wire IntSaturation_51U_32U_o_and_3_rgt;
  wire IntSaturation_51U_32U_o_IntSaturation_51U_32U_o_nor_3_rgt;
  wire IntSaturation_51U_32U_and_1_rgt;
  wire IntSaturation_51U_32U_o_and_1_rgt;
  wire and_2392_rgt;
  wire and_2399_rgt;
  wire and_2404_rgt;
  wire and_2405_rgt;
  wire and_2412_rgt;
  wire and_2414_rgt;
  wire and_2416_rgt;
  wire and_2417_rgt;
  wire and_2418_rgt;
  wire and_2419_rgt;
  wire and_2497_rgt;
  wire and_2499_rgt;
  wire and_2501_rgt;
  wire and_2503_rgt;
  wire and_2505_rgt;
  wire and_2507_rgt;
  wire and_2509_rgt;
  wire and_2511_rgt;
  wire and_2513_rgt;
  wire and_2515_rgt;
  wire and_2517_rgt;
  wire and_2519_rgt;
  wire [35:0] inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp;
  wire [35:0] inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp;
  wire [35:0] inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp;
  wire [35:0] inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_mux1h_1_itm;
  reg [1:0] reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_7_itm;
  reg [7:0] reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_7_1_itm;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_mux1h_3_itm;
  reg [1:0] reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_7_itm;
  reg [7:0] reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_7_1_itm;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_mux1h_6_itm;
  reg [1:0] reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_7_itm;
  reg [7:0] reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_7_1_itm;
  wire [48:0] inp_lookup_1_FpNormalize_8U_49U_else_lshift_itm;
  wire [48:0] inp_lookup_2_FpNormalize_8U_49U_else_lshift_itm;
  wire [48:0] inp_lookup_3_FpNormalize_8U_49U_else_lshift_itm;
  wire [48:0] inp_lookup_4_FpNormalize_8U_49U_else_lshift_itm;
  wire [9:0] FpMul_6U_10U_2_o_mant_mux1h_1_itm;
  reg [1:0] reg_FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_7_itm;
  reg [7:0] reg_FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_7_1_itm;
  wire [9:0] FpMul_6U_10U_2_o_mant_mux1h_3_itm;
  reg [1:0] reg_FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_7_itm;
  reg [7:0] reg_FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_7_1_itm;
  wire [9:0] FpMul_6U_10U_1_o_mant_mux1h_1_itm;
  reg [1:0] reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_6_itm;
  reg [7:0] reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_6_1_itm;
  wire [9:0] FpMul_6U_10U_2_o_mant_mux1h_5_itm;
  reg [1:0] reg_FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_7_itm;
  reg [7:0] reg_FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_7_1_itm;
  wire [22:0] inp_lookup_1_FpAdd_6U_10U_1_a_int_mant_p1_lshift_itm;
  wire [22:0] inp_lookup_1_FpAdd_6U_10U_1_b_int_mant_p1_lshift_itm;
  wire [22:0] inp_lookup_2_FpAdd_6U_10U_1_a_int_mant_p1_lshift_itm;
  wire [22:0] inp_lookup_2_FpAdd_6U_10U_1_b_int_mant_p1_lshift_itm;
  wire [22:0] inp_lookup_3_FpAdd_6U_10U_1_a_int_mant_p1_lshift_itm;
  wire [22:0] inp_lookup_3_FpAdd_6U_10U_1_b_int_mant_p1_lshift_itm;
  wire [22:0] inp_lookup_4_FpAdd_6U_10U_1_a_int_mant_p1_lshift_itm;
  wire [22:0] inp_lookup_4_FpAdd_6U_10U_1_b_int_mant_p1_lshift_itm;
  wire [22:0] inp_lookup_1_FpAdd_6U_10U_a_int_mant_p1_lshift_itm;
  wire [22:0] inp_lookup_1_FpAdd_6U_10U_b_int_mant_p1_lshift_itm;
  wire [22:0] inp_lookup_2_FpAdd_6U_10U_a_int_mant_p1_lshift_itm;
  wire [22:0] inp_lookup_2_FpAdd_6U_10U_b_int_mant_p1_lshift_itm;
  wire [22:0] inp_lookup_3_FpAdd_6U_10U_a_int_mant_p1_lshift_itm;
  wire [22:0] inp_lookup_3_FpAdd_6U_10U_b_int_mant_p1_lshift_itm;
  wire [22:0] inp_lookup_4_FpAdd_6U_10U_a_int_mant_p1_lshift_itm;
  wire [22:0] inp_lookup_4_FpAdd_6U_10U_b_int_mant_p1_lshift_itm;
  reg [7:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_10_17_1_itm;
  reg [8:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_10_17_1_1_itm;
  reg [7:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_10_17_1_itm;
  reg [8:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_10_17_1_1_itm;
  reg [7:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_10_17_1_itm;
  reg [8:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_10_17_1_1_itm;
  reg [7:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_10_17_1_itm;
  reg [8:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_10_17_1_1_itm;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_mux1h_4_itm;
  reg [1:0] reg_FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_7_itm;
  reg [7:0] reg_FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_7_1_itm;
  wire or_5695_itm;
  wire [30:0] mux1h_34_itm;
  reg [11:0] reg_chn_inp_in_crt_sva_2_606_576_itm;
  reg [18:0] reg_chn_inp_in_crt_sva_2_606_576_1_itm;
  wire or_5694_itm;
  wire [30:0] mux1h_36_itm;
  reg [11:0] reg_chn_inp_in_crt_sva_2_574_544_itm;
  reg [18:0] reg_chn_inp_in_crt_sva_2_574_544_1_itm;
  wire [30:0] mux1h_38_itm;
  reg [11:0] reg_chn_inp_in_crt_sva_2_510_480_itm;
  reg [18:0] reg_chn_inp_in_crt_sva_2_510_480_1_itm;
  wire or_5693_itm;
  wire [30:0] mux1h_40_itm;
  reg [11:0] reg_chn_inp_in_crt_sva_2_542_512_itm;
  reg [18:0] reg_chn_inp_in_crt_sva_2_542_512_1_itm;
  wire [30:0] mux1h_47_itm;
  reg [7:0] reg_chn_inp_in_crt_sva_5_30_0_itm;
  reg [22:0] reg_chn_inp_in_crt_sva_5_30_0_1_itm;
  wire [30:0] mux1h_49_itm;
  reg [7:0] reg_chn_inp_in_crt_sva_5_62_32_itm;
  reg [22:0] reg_chn_inp_in_crt_sva_5_62_32_1_itm;
  wire [30:0] mux1h_51_itm;
  reg [7:0] reg_chn_inp_in_crt_sva_5_94_64_itm;
  reg [22:0] reg_chn_inp_in_crt_sva_5_94_64_1_itm;
  wire [30:0] mux1h_53_itm;
  reg [7:0] reg_chn_inp_in_crt_sva_5_126_96_itm;
  reg [22:0] reg_chn_inp_in_crt_sva_5_126_96_1_itm;
  reg [4:0] reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_8_1_itm;
  wire [3:0] FpMul_6U_10U_1_o_expo_mux1h_23_itm;
  reg reg_FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_8_3_0_itm;
  reg [2:0] reg_FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_8_3_0_1_itm;
  wire [3:0] FpMul_6U_10U_1_o_expo_mux1h_29_itm;
  reg reg_FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_8_3_0_itm;
  reg [2:0] reg_FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_8_3_0_1_itm;
  wire [3:0] FpMul_6U_10U_1_o_expo_mux1h_35_itm;
  reg reg_FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_8_3_0_itm;
  reg [2:0] reg_FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_8_3_0_1_itm;
  wire [3:0] FpMul_6U_10U_1_o_expo_mux1h_41_itm;
  reg reg_FpMul_6U_10U_1_o_expo_lpi_1_dfm_8_3_0_itm;
  reg [2:0] reg_FpMul_6U_10U_1_o_expo_lpi_1_dfm_8_3_0_1_itm;
  reg [7:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_9_17_1_itm;
  reg [8:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_9_17_1_1_itm;
  reg [7:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_9_17_1_itm;
  reg [8:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_9_17_1_1_itm;
  reg [7:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_9_17_1_itm;
  reg [8:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_9_17_1_1_itm;
  reg [7:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_9_17_1_itm;
  reg [8:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_9_17_1_1_itm;
  reg [1:0] reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_7_itm;
  reg [7:0] reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_7_1_itm;
  reg [7:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_8_17_1_itm;
  reg [8:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_8_17_1_1_itm;
  reg [7:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_8_17_1_itm;
  reg [8:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_8_17_1_1_itm;
  reg [7:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_8_17_1_itm;
  reg [8:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_8_17_1_1_itm;
  reg [7:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_8_17_1_itm;
  reg [8:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_8_17_1_1_itm;
  wire [16:0] IntShiftRight_69U_6U_32U_obits_fixed_mux1h_25_itm;
  reg [7:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_7_17_1_itm;
  reg [8:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_7_17_1_1_itm;
  wire [16:0] IntShiftRight_69U_6U_32U_obits_fixed_mux1h_27_itm;
  reg [7:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_7_17_1_itm;
  reg [8:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_7_17_1_1_itm;
  wire [16:0] IntShiftRight_69U_6U_32U_obits_fixed_mux1h_29_itm;
  reg [7:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_7_17_1_itm;
  reg [8:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_7_17_1_1_itm;
  wire [16:0] IntShiftRight_69U_6U_32U_obits_fixed_mux1h_31_itm;
  reg [7:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_7_17_1_itm;
  reg [8:0] reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_7_17_1_1_itm;
  wire [9:0] inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_itm;
  wire [9:0] inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_itm;
  wire [22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_7_itm;
  wire [9:0] inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_itm;
  wire [9:0] FpMul_6U_10U_1_FpMul_6U_10U_1_FpMul_6U_10U_1_nor_4_itm;
  wire FpMul_6U_10U_1_or_11_itm;
  wire [9:0] FpMul_6U_10U_1_FpMul_6U_10U_1_FpMul_6U_10U_1_nor_5_itm;
  wire FpMul_6U_10U_1_or_10_itm;
  wire [9:0] FpMul_6U_10U_1_FpMul_6U_10U_1_FpMul_6U_10U_1_nor_7_itm;
  wire FpMul_6U_10U_1_or_8_itm;
  wire [9:0] inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_itm;
  wire [9:0] inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_itm;
  wire [9:0] inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_itm;
  wire [9:0] inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_itm;
  wire [9:0] inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_itm;
  wire [48:0] inp_lookup_1_FpNormalize_8U_49U_1_else_lshift_itm;
  wire [48:0] inp_lookup_2_FpNormalize_8U_49U_1_else_lshift_itm;
  wire [48:0] inp_lookup_3_FpNormalize_8U_49U_1_else_lshift_itm;
  wire [48:0] inp_lookup_4_FpNormalize_8U_49U_1_else_lshift_itm;
  wire [23:0] inp_lookup_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_itm;
  wire [22:0] inp_lookup_1_FpNormalize_6U_23U_1_else_lshift_itm;
  wire [23:0] inp_lookup_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_itm;
  wire [22:0] inp_lookup_2_FpNormalize_6U_23U_1_else_lshift_itm;
  wire [23:0] inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_itm;
  wire [22:0] inp_lookup_3_FpNormalize_6U_23U_1_else_lshift_itm;
  wire [23:0] inp_lookup_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_itm;
  wire [22:0] inp_lookup_4_FpNormalize_6U_23U_1_else_lshift_itm;
  wire [22:0] inp_lookup_1_FpNormalize_6U_23U_else_lshift_itm;
  wire [22:0] inp_lookup_2_FpNormalize_6U_23U_else_lshift_itm;
  wire [22:0] inp_lookup_3_FpNormalize_6U_23U_else_lshift_itm;
  wire [22:0] inp_lookup_4_FpNormalize_6U_23U_else_lshift_itm;
  wire mux_81_itm;
  wire mux_87_itm;
  wire mux_95_itm;
  wire mux_100_itm;
  wire mux_115_itm;
  wire mux_197_itm;
  wire mux_516_itm;
  wire mux_530_itm;
  wire mux_540_itm;
  wire mux_559_itm;
  wire mux_573_itm;
  wire mux_586_itm;
  wire mux_587_itm;
  wire mux_599_itm;
  wire mux_623_itm;
  wire mux_632_itm;
  wire mux_659_itm;
  wire mux_666_itm;
  wire mux_673_itm;
  wire mux_680_itm;
  wire mux_782_itm;
  wire mux_799_itm;
  wire mux_816_itm;
  wire mux_829_itm;
  wire mux_1066_itm;
  wire mux_1067_itm;
  wire mux_1172_itm;
  wire or_5684_itm;
  wire mux_1179_itm;
  wire or_5683_itm;
  wire mux_1182_itm;
  wire mux_1347_itm;
  wire mux_1362_itm;
  wire mux_1367_itm;
  wire mux_1558_itm;
  wire mux_1559_itm;
  wire mux_1560_itm;
  wire mux_1561_itm;
  wire FpAdd_8U_23U_else_2_and_tmp;
  wire [49:0] z_out;
  wire FpAdd_8U_23U_else_2_and_tmp_1;
  wire [49:0] z_out_1;
  wire FpAdd_8U_23U_else_2_and_tmp_2;
  wire [49:0] z_out_2;
  wire FpAdd_8U_23U_else_2_and_tmp_3;
  wire [49:0] z_out_3;
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp;
  wire [7:0] z_out_4;
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp_1;
  wire [7:0] z_out_5;
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp_2;
  wire [7:0] z_out_6;
  wire FpAdd_8U_23U_a_right_shift_qelse_and_tmp_3;
  wire [7:0] z_out_7;
  wire FpAdd_6U_10U_1_if_4_if_and_tmp;
  wire [6:0] z_out_8;
  wire [7:0] nl_z_out_8;
  wire FpAdd_6U_10U_1_if_4_if_and_tmp_1;
  wire [6:0] z_out_9;
  wire [7:0] nl_z_out_9;
  wire FpAdd_6U_10U_1_if_4_if_and_tmp_2;
  wire [6:0] z_out_10;
  wire [7:0] nl_z_out_10;
  wire FpAdd_6U_10U_1_if_4_if_and_tmp_3;
  wire [6:0] z_out_11;
  wire [7:0] nl_z_out_11;
  wire FpAdd_6U_10U_b_right_shift_qif_and_tmp;
  wire [5:0] z_out_12;
  wire FpAdd_6U_10U_b_right_shift_qif_and_tmp_1;
  wire [5:0] z_out_13;
  wire FpAdd_6U_10U_b_right_shift_qif_and_tmp_2;
  wire [5:0] z_out_14;
  wire FpAdd_6U_10U_b_right_shift_qif_and_tmp_3;
  wire [5:0] z_out_15;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_and_tmp;
  wire [9:0] z_out_16;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_and_tmp_1;
  wire [9:0] z_out_17;
  wire chn_inp_in_rsci_ld_core_psct_mx0c0;
  wire chn_inp_out_rsci_d_0_mx0c1;
  wire chn_inp_out_rsci_d_32_mx0c1;
  wire chn_inp_out_rsci_d_64_mx0c1;
  wire chn_inp_out_rsci_d_96_mx0c1;
  wire inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
  wire inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
  wire inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
  wire inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
  wire inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
  wire inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
  wire inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
  wire inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
  wire main_stage_v_1_mx0c1;
  wire FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0;
  wire inp_lookup_else_if_unequal_tmp_mx0w1;
  wire FpFractionToFloat_35U_6U_10U_1_o_mant_1_lpi_1_dfm_6_mx0c1;
  wire FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0;
  wire inp_lookup_else_if_unequal_tmp_1_mx0w1;
  wire FpFractionToFloat_35U_6U_10U_1_o_mant_2_lpi_1_dfm_6_mx0c1;
  wire FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0;
  wire FpFractionToFloat_35U_6U_10U_1_o_mant_3_lpi_1_dfm_6_mx0c1;
  wire inp_lookup_else_if_unequal_tmp_3_mx0w1;
  wire FpFractionToFloat_35U_6U_10U_1_o_mant_lpi_1_dfm_6_mx0c1;
  wire main_stage_v_2_mx0c1;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_19_mx0w1;
  wire inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_13_mx0w1;
  wire inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_7_mx0w1;
  wire inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_mx0w1;
  wire [48:0] FpAdd_8U_23U_addend_larger_asn_1_mx0w1;
  wire inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_mx0w1;
  wire main_stage_v_3_mx0c1;
  wire [7:0] FpAdd_8U_23U_o_expo_1_lpi_1_dfm_7_mx1w1;
  wire FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_3_5_mx1w1;
  wire [7:0] FpAdd_8U_23U_o_expo_2_lpi_1_dfm_7_mx1w1;
  wire FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_3_5_mx1w1;
  wire [7:0] FpAdd_8U_23U_o_expo_3_lpi_1_dfm_7_mx1w1;
  wire [9:0] FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_3_mx1w1;
  wire FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_3_5_mx1w1;
  wire [7:0] FpAdd_8U_23U_o_expo_lpi_1_dfm_7_mx1w1;
  wire main_stage_v_4_mx0c1;
  wire FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0;
  wire FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_3_4_mx0w0;
  wire [3:0] FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_3_3_0_mx0w0;
  wire FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0;
  wire FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_3_4_mx0w0;
  wire [3:0] FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_3_3_0_mx0w0;
  wire FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0;
  wire FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_3_4_mx0w0;
  wire [3:0] FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_3_3_0_mx0w0;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_9_mx0c0;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_9_mx0c2;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_9_mx0c3;
  wire FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_1_mx0w0;
  wire FpMul_6U_10U_2_o_expo_lpi_1_dfm_3_5_mx0w0;
  wire FpMul_6U_10U_2_o_expo_lpi_1_dfm_3_4_mx0w0;
  wire [3:0] FpMul_6U_10U_2_o_expo_lpi_1_dfm_3_3_0_mx0w0;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_9_1_mx0c0;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_9_1_mx0c2;
  wire main_stage_v_5_mx0c1;
  wire main_stage_v_6_mx0c1;
  wire [7:0] FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_2_mx0w0;
  wire [7:0] FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_2_mx0w0;
  wire [7:0] FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_2_mx0w0;
  wire [7:0] FpAdd_8U_23U_1_o_expo_lpi_1_dfm_2_mx0w0;
  wire main_stage_v_7_mx0c1;
  wire inp_lookup_1_FpMantRNE_24U_11U_else_and_svs_mx0w0;
  wire [2:0] FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_2_sva_mx0w0;
  wire [3:0] nl_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_2_sva_mx0w0;
  wire inp_lookup_2_FpMantRNE_24U_11U_else_and_svs_mx0w0;
  wire [2:0] FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_3_sva_mx0w0;
  wire [3:0] nl_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_3_sva_mx0w0;
  wire inp_lookup_3_FpMantRNE_24U_11U_else_and_svs_mx0w0;
  wire [22:0] FpAdd_8U_23U_1_asn_40_mx0w1;
  wire [2:0] FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_4_sva_mx0w0;
  wire [3:0] nl_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_4_sva_mx0w0;
  wire inp_lookup_4_FpMantRNE_24U_11U_else_and_svs_mx0w0;
  wire [2:0] FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_1_sva_mx0w0;
  wire [3:0] nl_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_1_sva_mx0w0;
  wire main_stage_v_8_mx0c1;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_7_5_mx0w0;
  wire [4:0] FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_7_4_0_mx0w0;
  wire [9:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_itm_mx0w0;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_7_5_mx0w0;
  wire [4:0] FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_7_4_0_mx0w0;
  wire [9:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_1_itm_mx0w0;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_7_5_mx0w0;
  wire [4:0] FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_7_4_0_mx0w0;
  wire [9:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_2_itm_mx0w0;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_7_5_mx0w0;
  wire [4:0] FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_7_4_0_mx0w0;
  wire [9:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_3_itm_mx0w0;
  wire main_stage_v_9_mx0c1;
  wire main_stage_v_10_mx0c1;
  wire main_stage_v_11_mx0c1;
  wire FpAdd_6U_10U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0;
  wire FpAdd_6U_10U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0;
  wire FpAdd_6U_10U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0;
  wire FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_1_mx0w0;
  wire main_stage_v_12_mx0c1;
  wire IsInf_6U_23U_land_1_lpi_1_dfm_mx1;
  wire [23:0] FpAdd_6U_10U_asn_23_mx0w1;
  wire [25:0] nl_FpAdd_6U_10U_asn_23_mx0w1;
  wire IsInf_6U_23U_land_2_lpi_1_dfm_mx1;
  wire [23:0] FpAdd_6U_10U_asn_20_mx0w1;
  wire [25:0] nl_FpAdd_6U_10U_asn_20_mx0w1;
  wire IsInf_6U_23U_land_3_lpi_1_dfm_mx1;
  wire [23:0] FpAdd_6U_10U_asn_17_mx0w1;
  wire [25:0] nl_FpAdd_6U_10U_asn_17_mx0w1;
  wire IsInf_6U_23U_land_lpi_1_dfm_mx1;
  wire [23:0] FpAdd_6U_10U_asn_mx0w1;
  wire [25:0] nl_FpAdd_6U_10U_asn_mx0w1;
  wire FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx0c0;
  wire FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx0c1;
  wire FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx0c2;
  wire [9:0] FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_3_mx0w0;
  wire [9:0] FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_3_mx0w0;
  wire [9:0] FpMul_6U_10U_2_o_mant_lpi_1_dfm_3_mx0w0;
  wire FpMantRNE_22U_11U_1_else_carry_1_sva;
  wire FpMantRNE_22U_11U_2_else_carry_1_sva_mx1w1;
  wire FpMantRNE_22U_11U_1_else_carry_3_sva;
  wire FpMantRNE_22U_11U_2_else_carry_3_sva_mx1w1;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_or_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_or_4_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_or_8_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_or_12_mx0w1;
  wire [21:0] FpMul_6U_10U_2_p_mant_p1_1_sva_mx3;
  wire [21:0] FpMul_6U_10U_2_p_mant_p1_2_sva_mx3;
  wire [21:0] FpMul_6U_10U_2_p_mant_p1_3_sva_mx3;
  wire [21:0] FpMul_6U_10U_2_p_mant_p1_sva_mx3;
  wire [21:0] FpMul_6U_10U_1_p_mant_p1_1_sva_mx3;
  wire [21:0] FpMul_6U_10U_1_p_mant_p1_2_sva_mx3;
  wire [5:0] FpMul_6U_10U_2_else_2_else_ac_int_cctor_2_sva_mx0w0;
  wire [6:0] nl_FpMul_6U_10U_2_else_2_else_ac_int_cctor_2_sva_mx0w0;
  wire [21:0] FpMul_6U_10U_1_p_mant_p1_3_sva_mx3;
  wire [5:0] FpMul_6U_10U_2_else_2_else_ac_int_cctor_3_sva_mx0w0;
  wire [6:0] nl_FpMul_6U_10U_2_else_2_else_ac_int_cctor_3_sva_mx0w0;
  wire [21:0] FpMul_6U_10U_1_p_mant_p1_sva_mx3;
  wire FpMantRNE_49U_24U_1_else_carry_1_sva_mx0w2;
  wire FpMantRNE_49U_24U_1_else_carry_2_sva_mx0w2;
  wire FpMantRNE_49U_24U_1_else_carry_3_sva_mx0w2;
  wire FpMantRNE_49U_24U_1_else_carry_sva_mx0w2;
  wire [9:0] FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_mx0w1;
  wire [9:0] FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_1_mx0w1;
  wire [9:0] FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_2_mx0w1;
  wire [9:0] FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_3_mx0w1;
  wire inp_lookup_if_unequal_tmp_1_mx0w0;
  wire FpMantRNE_22U_11U_1_else_carry_2_sva;
  wire FpMantRNE_22U_11U_2_else_carry_2_sva_mx1w1;
  wire FpMantRNE_22U_11U_1_else_carry_sva_mx0w1;
  wire FpMantRNE_22U_11U_2_else_carry_sva_mx0w2;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_or_8_mx0w1;
  wire IsNaN_6U_10U_1_land_1_lpi_1_dfm_mx0w0;
  wire IsNaN_6U_10U_1_land_2_lpi_1_dfm_mx0w0;
  wire IsNaN_6U_10U_1_land_3_lpi_1_dfm_mx0w0;
  wire IsNaN_6U_10U_1_land_lpi_1_dfm_mx0w0;
  wire [9:0] FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_1_lpi_1_dfm_5_mx1;
  wire inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0;
  wire inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0;
  wire inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0;
  wire inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0;
  wire [22:0] FpAdd_8U_23U_o_mant_1_lpi_1_dfm_2_mx2;
  wire [22:0] FpAdd_8U_23U_o_mant_2_lpi_1_dfm_2_mx2;
  wire [22:0] FpAdd_8U_23U_o_mant_3_lpi_1_dfm_2_mx2;
  wire [22:0] FpAdd_8U_23U_o_mant_lpi_1_dfm_2_mx2;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_3_mx0c1;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_3_mx0c1;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_3_lpi_1_dfm_3_mx0c1;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_3_mx0c1;
  wire IsNaN_6U_10U_4_land_1_lpi_1_dfm_mx0w1;
  wire IsNaN_6U_10U_4_land_2_lpi_1_dfm_mx0w1;
  wire IsNaN_6U_10U_4_land_3_lpi_1_dfm_mx0w1;
  wire IsNaN_6U_10U_4_land_lpi_1_dfm_mx0w1;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3_0_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w0;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3_0_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w0;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3_0_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w0;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3_0_mx0w0;
  wire [3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w0;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_4_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_8_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_12_mx0w1;
  wire IsNaN_6U_10U_2_land_1_lpi_1_dfm_mx0w0;
  wire IsNaN_6U_10U_2_land_2_lpi_1_dfm_mx0w0;
  wire IsNaN_6U_10U_2_land_3_lpi_1_dfm_mx0w0;
  wire IsNaN_6U_10U_2_land_lpi_1_dfm_mx0w0;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_or_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_or_4_mx0w1;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_or_12_mx0w1;
  wire FpAdd_8U_23U_o_sign_lpi_1_dfm_1_mx0c0;
  wire FpAdd_8U_23U_o_sign_lpi_1_dfm_1_mx0c1;
  wire FpAdd_8U_23U_o_sign_lpi_1_dfm_1_mx0c2;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_3_mx0c1;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_3_mx1;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_3_mx0c1;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_3_mx1;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_3_mx0c1;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_3_mx1;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_3_mx0c1;
  wire [9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_3_mx1;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_3_mx0c1;
  wire FpMantRNE_36U_11U_1_else_carry_1_sva;
  wire FpMantRNE_36U_11U_1_else_carry_2_sva;
  wire FpMantRNE_36U_11U_1_else_carry_3_sva;
  wire FpMantRNE_36U_11U_1_else_carry_sva;
  wire FpMantRNE_36U_11U_else_carry_1_sva;
  wire [35:0] FpMantRNE_36U_11U_i_data_2_sva;
  wire FpMantRNE_36U_11U_else_carry_2_sva;
  wire [35:0] FpMantRNE_36U_11U_i_data_3_sva;
  wire FpMantRNE_36U_11U_else_carry_3_sva;
  wire [35:0] FpMantRNE_36U_11U_i_data_4_sva;
  wire FpMantRNE_36U_11U_else_carry_sva;
  wire [35:0] FpMantRNE_36U_11U_i_data_sva;
  wire FpAdd_8U_23U_and_tmp;
  wire FpMantRNE_49U_24U_else_carry_1_sva;
  wire [48:0] FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_and_1_tmp;
  wire FpMantRNE_49U_24U_else_carry_2_sva;
  wire [48:0] FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_and_2_tmp;
  wire FpMantRNE_49U_24U_else_carry_3_sva;
  wire [48:0] FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0;
  wire FpAdd_8U_23U_and_3_tmp;
  wire FpMantRNE_49U_24U_else_carry_sva;
  wire [48:0] FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0;
  wire [22:0] FpAdd_6U_10U_1_addend_larger_qr_1_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_1_addend_smaller_qr_1_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_1_addend_larger_qr_2_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_1_addend_smaller_qr_2_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_1_addend_larger_qr_3_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_1_addend_smaller_qr_3_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_1_addend_larger_qr_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_1_addend_smaller_qr_lpi_1_dfm_mx0;
  wire [5:0] FpAdd_6U_10U_1_o_expo_1_sva_1;
  wire [6:0] nl_FpAdd_6U_10U_1_o_expo_1_sva_1;
  wire [22:0] FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_1;
  wire FpMantRNE_23U_11U_1_else_carry_1_sva;
  wire [21:0] FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0;
  wire [9:0] FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_2_lpi_1_dfm_5_mx0;
  wire [5:0] FpAdd_6U_10U_1_o_expo_2_sva_1;
  wire [6:0] nl_FpAdd_6U_10U_1_o_expo_2_sva_1;
  wire [22:0] FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_1;
  wire FpMantRNE_23U_11U_1_else_carry_2_sva;
  wire [21:0] FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0;
  wire [9:0] FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_3_lpi_1_dfm_5_mx0;
  wire [5:0] FpAdd_6U_10U_1_o_expo_3_sva_1;
  wire [6:0] nl_FpAdd_6U_10U_1_o_expo_3_sva_1;
  wire [22:0] FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_1;
  wire FpMantRNE_23U_11U_1_else_carry_3_sva;
  wire [21:0] FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0;
  wire [9:0] FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_lpi_1_dfm_5_mx0;
  wire [5:0] FpAdd_6U_10U_1_o_expo_sva_1;
  wire [6:0] nl_FpAdd_6U_10U_1_o_expo_sva_1;
  wire [22:0] FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_1_o_expo_lpi_1_dfm_1;
  wire FpMantRNE_23U_11U_1_else_carry_sva;
  wire [21:0] FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0;
  wire IsNaN_6U_23U_2_land_1_lpi_1_dfm;
  wire IsNaN_6U_23U_2_land_2_lpi_1_dfm;
  wire IsNaN_6U_23U_2_land_3_lpi_1_dfm;
  wire IsNaN_6U_23U_2_land_lpi_1_dfm;
  wire [23:0] FpAdd_6U_10U_int_mant_p1_1_sva;
  wire [24:0] nl_FpAdd_6U_10U_int_mant_p1_1_sva;
  wire [22:0] FpAdd_6U_10U_addend_larger_qr_1_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_addend_smaller_qr_1_lpi_1_dfm_mx0;
  wire [23:0] FpAdd_6U_10U_int_mant_p1_2_sva;
  wire [24:0] nl_FpAdd_6U_10U_int_mant_p1_2_sva;
  wire [22:0] FpAdd_6U_10U_addend_larger_qr_2_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_addend_smaller_qr_2_lpi_1_dfm_mx0;
  wire [23:0] FpAdd_6U_10U_int_mant_p1_3_sva;
  wire [24:0] nl_FpAdd_6U_10U_int_mant_p1_3_sva;
  wire [22:0] FpAdd_6U_10U_addend_larger_qr_3_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_addend_smaller_qr_3_lpi_1_dfm_mx0;
  wire [23:0] FpAdd_6U_10U_int_mant_p1_sva;
  wire [24:0] nl_FpAdd_6U_10U_int_mant_p1_sva;
  wire [22:0] FpAdd_6U_10U_addend_larger_qr_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_addend_smaller_qr_lpi_1_dfm_mx0;
  wire [5:0] FpAdd_6U_10U_o_expo_1_sva_1;
  wire [6:0] nl_FpAdd_6U_10U_o_expo_1_sva_1;
  wire [22:0] FpAdd_6U_10U_int_mant_2_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_o_expo_1_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_o_expo_1_sva_4;
  wire [6:0] nl_FpAdd_6U_10U_o_expo_1_sva_4;
  wire [21:0] FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_else_carry_1_sva;
  wire [9:0] FpAdd_6U_10U_o_mant_1_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_and_ssc;
  wire FpAdd_6U_10U_and_6_ssc;
  wire [5:0] FpAdd_6U_10U_o_expo_2_sva_1;
  wire [6:0] nl_FpAdd_6U_10U_o_expo_2_sva_1;
  wire [22:0] FpAdd_6U_10U_int_mant_3_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_o_expo_2_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_o_expo_2_sva_4;
  wire [6:0] nl_FpAdd_6U_10U_o_expo_2_sva_4;
  wire [21:0] FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_else_carry_2_sva;
  wire [9:0] FpAdd_6U_10U_o_mant_2_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_and_29_ssc;
  wire FpAdd_6U_10U_and_13_ssc;
  wire [5:0] FpAdd_6U_10U_o_expo_3_sva_1;
  wire [6:0] nl_FpAdd_6U_10U_o_expo_3_sva_1;
  wire [22:0] FpAdd_6U_10U_int_mant_4_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_o_expo_3_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_o_expo_3_sva_4;
  wire [6:0] nl_FpAdd_6U_10U_o_expo_3_sva_4;
  wire [21:0] FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_else_carry_3_sva;
  wire [9:0] FpAdd_6U_10U_o_mant_3_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_and_31_ssc;
  wire FpAdd_6U_10U_and_19_ssc;
  wire [5:0] FpAdd_6U_10U_o_expo_sva_1;
  wire [6:0] nl_FpAdd_6U_10U_o_expo_sva_1;
  wire [22:0] FpAdd_6U_10U_int_mant_1_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_o_expo_lpi_1_dfm_1;
  wire [5:0] FpAdd_6U_10U_o_expo_sva_4;
  wire [6:0] nl_FpAdd_6U_10U_o_expo_sva_4;
  wire [21:0] FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0;
  wire FpMantRNE_23U_11U_else_carry_sva;
  wire [9:0] FpAdd_6U_10U_o_mant_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_and_33_ssc;
  wire FpAdd_6U_10U_and_25_ssc;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_1_sva;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm;
  wire [10:0] FpMantRNE_36U_11U_else_ac_int_cctor_2_sva;
  wire [11:0] nl_FpMantRNE_36U_11U_else_ac_int_cctor_2_sva;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_2_sva;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm;
  wire [10:0] FpMantRNE_36U_11U_else_ac_int_cctor_3_sva;
  wire [11:0] nl_FpMantRNE_36U_11U_else_ac_int_cctor_3_sva;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_3_sva;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm;
  wire [10:0] FpMantRNE_36U_11U_else_ac_int_cctor_4_sva;
  wire [11:0] nl_FpMantRNE_36U_11U_else_ac_int_cctor_4_sva;
  wire [48:0] FpAdd_8U_23U_a_int_mant_p1_sva;
  wire [7:0] FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm;
  wire [10:0] FpMantRNE_36U_11U_else_ac_int_cctor_sva;
  wire [11:0] nl_FpMantRNE_36U_11U_else_ac_int_cctor_sva;
  wire IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_ovfl_1_sva;
  wire IntSignedShiftRight_50U_5U_32U_obits_fixed_and_unfl_1_sva;
  wire [19:0] FpMul_6U_10U_2_p_mant_20_1_1_lpi_1_dfm_3_mx0;
  wire IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_ovfl_2_sva;
  wire IntSignedShiftRight_50U_5U_32U_obits_fixed_and_unfl_2_sva;
  wire [19:0] FpMul_6U_10U_2_p_mant_20_1_2_lpi_1_dfm_3_mx0;
  wire IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_ovfl_3_sva;
  wire IntSignedShiftRight_50U_5U_32U_obits_fixed_and_unfl_3_sva;
  wire [19:0] FpMul_6U_10U_2_p_mant_20_1_3_lpi_1_dfm_3_mx0;
  wire IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_ovfl_sva;
  wire IntSignedShiftRight_50U_5U_32U_obits_fixed_and_unfl_sva;
  wire [19:0] FpMul_6U_10U_2_p_mant_20_1_lpi_1_dfm_3_mx0;
  wire [19:0] FpMul_6U_10U_1_p_mant_20_1_2_lpi_1_dfm_3_mx0;
  wire [48:0] FpAdd_8U_23U_1_addend_larger_asn_19_mx0w1;
  wire [48:0] FpAdd_8U_23U_1_addend_larger_qr_1_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_1_addend_smaller_qr_1_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_1_a_int_mant_p1_1_sva;
  wire [7:0] FpAdd_8U_23U_1_b_right_shift_qr_1_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_1_a_right_shift_qr_1_lpi_1_dfm;
  wire [48:0] FpAdd_8U_23U_1_addend_larger_asn_13_mx0w1;
  wire [48:0] FpAdd_8U_23U_1_addend_larger_qr_2_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_1_addend_smaller_qr_2_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_1_a_int_mant_p1_2_sva;
  wire [7:0] FpAdd_8U_23U_1_b_right_shift_qr_2_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_1_a_right_shift_qr_2_lpi_1_dfm;
  wire [48:0] FpAdd_8U_23U_1_addend_larger_asn_7_mx0w1;
  wire [48:0] FpAdd_8U_23U_1_addend_larger_qr_3_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_1_addend_smaller_qr_3_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_1_a_int_mant_p1_3_sva;
  wire [7:0] FpAdd_8U_23U_1_b_right_shift_qr_3_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_1_a_right_shift_qr_3_lpi_1_dfm;
  wire [48:0] FpAdd_8U_23U_1_addend_larger_asn_1_mx0w1;
  wire [48:0] FpAdd_8U_23U_1_addend_larger_qr_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_1_addend_smaller_qr_lpi_1_dfm_mx0;
  wire [48:0] FpAdd_8U_23U_1_a_int_mant_p1_sva;
  wire [7:0] FpAdd_8U_23U_1_b_right_shift_qr_lpi_1_dfm;
  wire [7:0] FpAdd_8U_23U_1_a_right_shift_qr_lpi_1_dfm;
  wire [5:0] FpAdd_6U_10U_1_o_expo_1_sva_4;
  wire [6:0] nl_FpAdd_6U_10U_1_o_expo_1_sva_4;
  wire FpAdd_6U_10U_1_and_ssc;
  wire FpAdd_6U_10U_1_and_6_ssc;
  wire [5:0] FpAdd_6U_10U_1_o_expo_2_sva_4;
  wire [6:0] nl_FpAdd_6U_10U_1_o_expo_2_sva_4;
  wire FpAdd_6U_10U_1_and_29_ssc;
  wire FpAdd_6U_10U_1_and_13_ssc;
  wire [5:0] FpAdd_6U_10U_1_o_expo_3_sva_4;
  wire [6:0] nl_FpAdd_6U_10U_1_o_expo_3_sva_4;
  wire FpAdd_6U_10U_1_and_31_ssc;
  wire FpAdd_6U_10U_1_and_19_ssc;
  wire [5:0] FpAdd_6U_10U_1_o_expo_sva_4;
  wire [6:0] nl_FpAdd_6U_10U_1_o_expo_sva_4;
  wire FpAdd_6U_10U_1_and_33_ssc;
  wire FpAdd_6U_10U_1_and_25_ssc;
  wire [80:0] IntSignedShiftRight_50U_5U_32U_mbits_fixed_1_sva;
  wire [80:0] IntSignedShiftRight_50U_5U_32U_mbits_fixed_2_sva;
  wire [80:0] IntSignedShiftRight_50U_5U_32U_mbits_fixed_3_sva;
  wire [80:0] IntSignedShiftRight_50U_5U_32U_mbits_fixed_sva;
  wire [9:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_9_0_1_lpi_1_dfm_2_mx0;
  wire [9:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_9_0_2_lpi_1_dfm_2_mx0;
  wire [9:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_9_0_3_lpi_1_dfm_2_mx0;
  wire [9:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_9_0_lpi_1_dfm_2_mx0;
  wire [52:0] inp_lookup_else_else_o_acc_psp_1_sva;
  wire [53:0] nl_inp_lookup_else_else_o_acc_psp_1_sva;
  wire [52:0] inp_lookup_else_else_o_acc_psp_2_sva;
  wire [53:0] nl_inp_lookup_else_else_o_acc_psp_2_sva;
  wire [52:0] inp_lookup_else_else_o_acc_psp_3_sva;
  wire [53:0] nl_inp_lookup_else_else_o_acc_psp_3_sva;
  wire [52:0] inp_lookup_else_else_o_acc_psp_sva;
  wire [53:0] nl_inp_lookup_else_else_o_acc_psp_sva;
  wire FpNormalize_8U_49U_1_oelse_not_9;
  wire FpNormalize_8U_49U_1_oelse_not_11;
  wire FpNormalize_8U_49U_1_oelse_not_13;
  wire FpNormalize_8U_49U_1_oelse_not_15;
  wire FpAdd_6U_10U_1_asn_124;
  wire FpNormalize_6U_23U_1_oelse_not_9;
  wire FpAdd_6U_10U_1_asn_126;
  wire FpNormalize_6U_23U_1_oelse_not_11;
  wire FpAdd_6U_10U_1_asn_128;
  wire FpNormalize_6U_23U_1_oelse_not_13;
  wire FpAdd_6U_10U_1_asn_130;
  wire FpNormalize_6U_23U_1_oelse_not_15;
  wire FpAdd_6U_10U_asn_87;
  wire FpAdd_6U_10U_asn_89;
  wire FpAdd_6U_10U_asn_91;
  wire FpAdd_6U_10U_asn_93;
  wire [20:0] FpMul_6U_10U_2_p_mant_p1_1_sva_mx1_20_0;
  wire [20:0] FpMul_6U_10U_2_p_mant_p1_2_sva_mx1_20_0;
  wire [20:0] FpMul_6U_10U_2_p_mant_p1_3_sva_mx1_20_0;
  wire [20:0] FpMul_6U_10U_2_p_mant_p1_sva_mx1_20_0;
  wire [20:0] FpMul_6U_10U_1_p_mant_p1_1_sva_mx1_20_0;
  wire [20:0] FpMul_6U_10U_1_p_mant_p1_2_sva_mx1_20_0;
  wire [20:0] FpMul_6U_10U_1_p_mant_p1_3_sva_mx1_20_0;
  wire [20:0] FpMul_6U_10U_1_p_mant_p1_sva_mx1_20_0;
  wire [5:0] libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_8;
  wire [5:0] libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_9;
  wire [5:0] libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_10;
  wire [5:0] libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_11;
  wire [5:0] libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_12;
  wire [5:0] libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_13;
  wire [5:0] libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_14;
  wire [5:0] libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_15;
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_8;
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_9;
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_10;
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_11;
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_12;
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_13;
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_14;
  wire [5:0] libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_15;
  wire [4:0] libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_8;
  wire [4:0] libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_9;
  wire [4:0] libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_10;
  wire [4:0] libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_11;
  wire [3:0] libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_16;
  wire [3:0] libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_17;
  wire [3:0] libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_18;
  wire [3:0] libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_19;
  wire [4:0] libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_12;
  wire [4:0] libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_13;
  wire [4:0] libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_14;
  wire [4:0] libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_15;
  wire [3:0] libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_20;
  wire [3:0] libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_21;
  wire [3:0] libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_22;
  wire [3:0] libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_23;
  wire [3:0] libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_24;
  wire [3:0] libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_25;
  wire [3:0] libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_26;
  wire [3:0] libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_27;
  wire FpAdd_8U_23U_o_expo_and_14_ssc;
  reg [1:0] reg_FpAdd_8U_23U_o_expo_1_lpi_1_dfm_12_tmp;
  reg [5:0] reg_FpAdd_8U_23U_o_expo_1_lpi_1_dfm_12_tmp_1;
  wire FpAdd_8U_23U_o_expo_and_13_ssc;
  reg [1:0] reg_FpAdd_8U_23U_o_expo_2_lpi_1_dfm_12_tmp;
  reg [5:0] reg_FpAdd_8U_23U_o_expo_2_lpi_1_dfm_12_tmp_1;
  wire FpAdd_8U_23U_o_expo_and_12_ssc;
  reg [1:0] reg_FpAdd_8U_23U_o_expo_lpi_1_dfm_12_tmp;
  reg [5:0] reg_FpAdd_8U_23U_o_expo_lpi_1_dfm_12_tmp_1;
  reg reg_FpMul_6U_10U_o_expo_lpi_1_dfm_6_5_4_tmp;
  reg reg_FpMul_6U_10U_o_expo_lpi_1_dfm_6_5_4_tmp_1;
  reg reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_15_tmp;
  reg reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_15_tmp_1;
  reg reg_FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_5_4_tmp;
  reg reg_FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_5_4_tmp_1;
  reg reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_15_tmp;
  reg reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_15_tmp_1;
  reg reg_FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_5_4_tmp;
  reg reg_FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_5_4_tmp_1;
  reg reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_15_tmp;
  reg reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_15_tmp_1;
  reg reg_FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_5_4_tmp;
  reg reg_FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_5_4_tmp_1;
  reg reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_15_tmp;
  reg reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_15_tmp_1;
  reg reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_16_tmp;
  reg reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_16_tmp_1;
  reg reg_FpAdd_6U_10U_qr_lpi_1_dfm_5_4_tmp;
  reg reg_FpAdd_6U_10U_qr_lpi_1_dfm_5_4_tmp_1;
  reg reg_FpAdd_6U_10U_qr_lpi_1_dfm_3_5_4_tmp;
  reg reg_FpAdd_6U_10U_qr_lpi_1_dfm_3_5_4_tmp_1;
  reg reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_16_tmp;
  reg reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_16_tmp_1;
  reg reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_5_4_tmp;
  reg reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_5_4_tmp_1;
  reg reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_3_5_4_tmp;
  reg reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_3_5_4_tmp_1;
  reg reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_16_tmp;
  reg reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_16_tmp_1;
  reg reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_5_4_tmp;
  reg reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_5_4_tmp_1;
  reg reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_3_5_4_tmp;
  reg reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_3_5_4_tmp_1;
  reg reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_16_tmp;
  reg reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_16_tmp_1;
  reg reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_5_4_tmp;
  reg reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_5_4_tmp_1;
  reg reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_3_5_4_tmp;
  reg reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_3_5_4_tmp_1;
  reg reg_FpAdd_6U_10U_qr_lpi_1_dfm_4_5_4_tmp;
  reg reg_FpAdd_6U_10U_qr_lpi_1_dfm_4_5_4_tmp_1;
  reg reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_4_5_4_tmp;
  reg reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_4_5_4_tmp_1;
  reg reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_4_5_4_tmp;
  reg reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_4_5_4_tmp_1;
  reg reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_4_5_4_tmp;
  reg reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_4_5_4_tmp_1;
  reg reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_17_tmp;
  reg reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_17_tmp_1;
  reg reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_17_tmp;
  reg reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_17_tmp_1;
  reg reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_17_tmp;
  reg reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_17_tmp_1;
  reg reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_17_tmp;
  reg reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_17_tmp_1;
  wire and_1185_tmp;
  wire mux_1958_m1c;
  wire mux_1904_tmp;
  wire mux_1903_tmp;
  wire mux_1902_tmp;
  wire mux_1901_tmp;
  wire and_3875_ssc;
  reg [1:0] reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_8_itm_4_3;
  reg [2:0] reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_8_itm_2_0;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_12_cse;
  wire FpAdd_8U_23U_is_a_greater_oelse_and_cse;
  wire IntLeadZero_35U_1_leading_sign_35_0_rtn_and_4_cse;
  wire FpFractionToFloat_35U_6U_10U_1_if_else_else_and_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_15_cse;
  wire FpAdd_8U_23U_is_a_greater_oelse_FpAdd_8U_23U_is_a_greater_oelse_or_19_cse;
  wire IntLeadZero_35U_1_leading_sign_35_0_rtn_and_5_cse;
  wire FpFractionToFloat_35U_6U_10U_1_if_else_else_and_1_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_18_cse;
  wire FpAdd_8U_23U_is_a_greater_oelse_and_2_cse;
  wire IntLeadZero_35U_1_leading_sign_35_0_rtn_and_6_cse;
  wire FpFractionToFloat_35U_6U_10U_1_if_else_else_and_2_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_21_cse;
  wire FpAdd_8U_23U_is_a_greater_oelse_FpAdd_8U_23U_is_a_greater_oelse_or_17_cse;
  wire IntLeadZero_35U_1_leading_sign_35_0_rtn_and_7_cse;
  wire FpFractionToFloat_35U_6U_10U_1_if_else_else_and_3_cse;
  wire cfg_precision_and_cse;
  wire FpAdd_8U_23U_addend_larger_and_cse;
  wire FpAdd_8U_23U_is_addition_and_cse;
  wire FpFractionToFloat_35U_6U_10U_is_zero_FpFractionToFloat_35U_6U_10U_is_zero_or_3_cse;
  wire or_5873_cse;
  wire nor_1896_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_17_cse;
  wire FpAdd_8U_23U_addend_larger_and_1_cse;
  wire FpAdd_8U_23U_is_addition_and_2_cse;
  wire cfg_precision_and_4_cse;
  wire FpFractionToFloat_35U_6U_10U_is_zero_FpFractionToFloat_35U_6U_10U_is_zero_or_2_cse;
  wire or_5889_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_19_cse;
  wire FpAdd_8U_23U_addend_larger_and_2_cse;
  wire FpAdd_8U_23U_is_addition_and_4_cse;
  wire FpFractionToFloat_35U_6U_10U_is_zero_FpFractionToFloat_35U_6U_10U_is_zero_or_1_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_21_cse;
  wire FpAdd_8U_23U_addend_larger_and_3_cse;
  wire FpAdd_8U_23U_is_addition_and_6_cse;
  wire FpFractionToFloat_35U_6U_10U_is_zero_FpFractionToFloat_35U_6U_10U_is_zero_or_cse;
  wire or_6160_cse;
  wire or_5904_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_24_cse;
  wire nand_602_cse_1;
  wire IntSignedShiftRight_50U_5U_32U_obits_fixed_and_cse;
  wire and_3624_cse;
  wire FpMul_6U_10U_2_oelse_1_and_4_cse;
  wire IntSignedShiftRight_50U_5U_32U_obits_fixed_and_3_cse;
  wire IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_2_cse;
  wire IntSignedShiftRight_50U_5U_32U_obits_fixed_and_6_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_or_cse;
  wire IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_1_cse;
  wire IntSignedShiftRight_50U_5U_32U_obits_fixed_and_9_cse;
  wire IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_cse;
  wire FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_or_6_cse;
  wire FpMul_6U_10U_2_o_expo_and_cse;
  wire inp_lookup_else_if_a0_and_12_cse;
  wire FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_or_5_cse;
  wire cfg_precision_and_12_cse;
  wire FpMul_6U_10U_2_o_expo_and_3_cse;
  wire inp_lookup_else_if_a0_and_14_cse;
  wire FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_or_4_cse;
  wire FpMul_6U_10U_2_o_expo_and_6_cse;
  wire inp_lookup_else_if_a0_and_16_cse;
  wire FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_4_cse;
  wire FpMul_6U_10U_2_o_expo_and_9_cse;
  wire inp_lookup_else_if_a0_and_18_cse;
  wire or_5950_cse;
  wire and_4141_cse;
  wire and_3637_cse;
  wire xnor_6_cse;
  wire cfg_precision_and_16_cse;
  wire or_5967_cse;
  wire and_4136_cse;
  wire and_3663_cse;
  wire xnor_4_cse;
  wire or_5985_cse;
  wire and_3689_cse;
  wire xnor_2_cse;
  wire and_4126_cse;
  wire IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_4_cse;
  wire cfg_precision_and_20_cse;
  wire IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_3_cse;
  reg reg_inp_lookup_3_FpMantRNE_49U_24U_1_else_and_svs_1_cse;
  wire IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_2_cse;
  wire IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_1_cse;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_and_cse;
  wire cfg_precision_and_24_cse;
  wire FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_14_cse;
  wire FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_13_cse;
  wire FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_12_cse;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_and_cse;
  reg reg_FpMul_6U_10U_lor_3_lpi_1_dfm_3_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_12_cse;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_and_2_cse;
  reg reg_FpMul_6U_10U_lor_4_lpi_1_dfm_3_cse;
  wire cfg_precision_and_28_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_13_cse;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_and_4_cse;
  reg reg_FpMul_6U_10U_lor_5_lpi_1_dfm_3_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_14_cse;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_and_6_cse;
  reg reg_FpMul_6U_10U_lor_lpi_1_dfm_3_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_15_cse;
  wire IsNaN_6U_10U_2_aelse_and_cse;
  wire IsNaN_6U_10U_2_aelse_and_1_cse;
  wire IsNaN_6U_10U_2_aelse_and_2_cse;
  wire IsNaN_6U_10U_2_aelse_and_3_cse;
  wire chn_inp_in_flow_and_32_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_cse;
  wire FpMul_6U_10U_o_expo_and_8_cse;
  reg reg_inp_lookup_1_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_13_cse;
  wire FpMul_6U_10U_o_expo_and_10_cse;
  reg reg_inp_lookup_2_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_15_cse;
  wire FpMul_6U_10U_o_expo_and_12_cse;
  reg reg_inp_lookup_3_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_17_cse;
  wire FpMul_6U_10U_o_expo_and_14_cse;
  reg reg_inp_lookup_4_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse;
  wire chn_inp_in_flow_and_36_cse;
  wire FpAdd_6U_10U_is_addition_and_cse;
  wire FpAdd_6U_10U_is_addition_and_2_cse;
  wire FpAdd_6U_10U_is_addition_and_4_cse;
  wire FpAdd_6U_10U_is_addition_and_6_cse;
  wire chn_inp_in_flow_and_40_cse;
  wire FpAdd_6U_10U_and_43_cse;
  reg reg_FpNormalize_6U_23U_lor_1_lpi_1_dfm_4_cse;
  wire IsNaN_6U_10U_3_aelse_and_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_19_cse;
  wire FpAdd_6U_10U_and_45_cse;
  reg reg_FpNormalize_6U_23U_lor_2_lpi_1_dfm_4_cse;
  wire IsNaN_6U_10U_3_aelse_and_1_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_21_cse;
  wire FpAdd_6U_10U_and_47_cse;
  wire IsNaN_6U_10U_3_aelse_and_2_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_23_cse;
  wire FpAdd_6U_10U_and_49_cse;
  reg reg_FpNormalize_6U_23U_lor_lpi_1_dfm_4_cse;
  wire IsNaN_6U_10U_3_aelse_and_3_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_25_cse;
  wire inp_lookup_and_cse;
  wire FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_and_cse;
  wire FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_cse;
  wire FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_and_6_cse;
  wire FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_2_cse;
  wire FpAdd_6U_10U_and_51_cse;
  wire FpAdd_6U_10U_and_53_cse;
  wire FpAdd_6U_10U_and_55_cse;
  wire FpAdd_6U_10U_and_57_cse;
  wire FpNormalize_6U_23U_1_if_FpNormalize_6U_23U_1_if_or_3_cse;
  wire FpMul_6U_10U_2_else_2_else_if_FpMul_6U_10U_2_else_2_else_if_or_3_cse;
  wire inp_lookup_else_if_a0_and_8_cse;
  wire FpMul_6U_10U_2_else_2_else_if_FpMul_6U_10U_2_else_2_else_if_or_2_cse;
  wire inp_lookup_else_if_a0_and_9_cse;
  wire inp_lookup_else_if_a0_and_10_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_37_cse;
  wire inp_lookup_else_if_a0_and_11_cse;
  wire IsNaN_8U_23U_aelse_and_cse;
  wire IsZero_8U_23U_1_and_cse;
  wire IsZero_8U_23U_1_and_1_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_24_cse;
  wire FpFractionToFloat_35U_6U_10U_1_o_mant_and_12_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_27_cse;
  wire FpFractionToFloat_35U_6U_10U_1_o_mant_and_13_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_and_cse;
  wire FpFractionToFloat_35U_6U_10U_1_o_mant_and_14_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_33_cse;
  wire FpFractionToFloat_35U_6U_10U_1_o_mant_and_15_cse;
  wire FpMul_6U_10U_2_oelse_1_FpMul_6U_10U_2_oelse_1_or_11_cse;
  wire IsZero_8U_23U_3_and_3_cse;
  wire IsNaN_8U_23U_2_aelse_IsNaN_8U_23U_2_aelse_or_cse;
  wire FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_1_cse;
  wire FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_2_cse;
  wire FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_3_cse;
  wire FpAdd_6U_10U_1_is_addition_and_cse;
  wire FpAdd_6U_10U_1_is_addition_and_1_cse;
  wire FpAdd_6U_10U_1_is_addition_and_2_cse;
  wire FpAdd_6U_10U_1_is_addition_and_3_cse;
  wire FpMul_6U_10U_2_o_expo_and_12_cse;
  wire FpMul_6U_10U_2_o_expo_and_15_cse;
  wire FpMul_6U_10U_2_o_expo_and_18_cse;
  wire FpMul_6U_10U_2_o_expo_and_21_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_or_15_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_or_14_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_or_13_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_or_12_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_28_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_31_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_34_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_37_cse;
  wire FpAdd_6U_10U_is_a_greater_and_cse;
  wire FpAdd_6U_10U_is_a_greater_and_2_cse;
  wire IsZero_6U_10U_3_and_cse;
  wire IsZero_6U_10U_3_and_1_cse;
  wire IsZero_6U_10U_3_and_2_cse;
  wire IsZero_6U_10U_3_and_3_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_9_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_8_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_7_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_6_cse;
  wire FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_4_cse;
  wire FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_5_cse;
  wire FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_6_cse;
  wire FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_7_cse;
  wire FpAdd_8U_23U_is_addition_and_11_cse;
  wire FpAdd_8U_23U_is_addition_and_10_cse;
  wire FpAdd_8U_23U_is_addition_and_9_cse;
  wire IsNaN_8U_23U_1_and_cse;
  wire FpMul_6U_10U_1_o_expo_FpMul_6U_10U_1_o_expo_or_7_cse;
  wire FpMul_6U_10U_1_o_expo_FpMul_6U_10U_1_o_expo_or_5_cse;
  wire FpMul_6U_10U_1_o_expo_FpMul_6U_10U_1_o_expo_or_3_cse;
  wire FpMul_6U_10U_1_o_expo_FpMul_6U_10U_1_o_expo_or_1_cse;
  wire FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_8_cse;
  wire FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_9_cse;
  wire FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_10_cse;
  wire FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_11_cse;
  wire inp_lookup_else_and_23_cse;
  wire inp_lookup_else_and_22_cse;
  wire inp_lookup_else_and_21_cse;
  wire inp_lookup_else_and_20_cse;
  wire FpMul_6U_10U_oelse_and_cse;
  wire FpMul_6U_10U_oelse_and_2_cse;
  wire FpMul_6U_10U_oelse_and_4_cse;
  wire FpMul_6U_10U_oelse_and_6_cse;
  wire FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_12_cse;
  wire FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_13_cse;
  wire FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_14_cse;
  wire FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_15_cse;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_if_and_2_cse;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_if_and_4_cse;
  wire FpWidthDec_8U_23U_6U_10U_0U_1U_if_and_6_cse;
  wire IsNaN_6U_10U_5_aelse_and_4_cse;
  wire FpMantRNE_49U_24U_1_else_and_6_cse;
  wire FpMantRNE_49U_24U_1_else_and_4_cse;
  wire FpMantRNE_49U_24U_1_else_and_2_cse;
  wire FpMantRNE_49U_24U_1_else_and_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_100_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_103_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_106_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_109_cse;
  wire IsZero_6U_10U_1_and_12_cse;
  wire or_5890_cse;
  wire or_5882_cse;
  wire nor_1869_cse;
  wire or_5896_cse;
  wire or_2676_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_18_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_20_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_22_cse;
  wire and_3361_cse_1;
  wire FpMul_6U_10U_2_oelse_1_and_5_cse;
  wire FpMul_6U_10U_2_oelse_1_and_6_cse;
  wire FpMul_6U_10U_2_oelse_1_and_7_cse;
  wire FpAdd_8U_23U_1_is_a_greater_oelse_and_cse;
  wire FpAdd_8U_23U_1_is_a_greater_oelse_and_1_cse;
  wire FpAdd_8U_23U_1_is_a_greater_oelse_and_2_cse;
  wire IsNaN_6U_10U_4_aelse_and_cse;
  wire FpAdd_8U_23U_1_is_a_greater_oelse_and_3_cse;
  wire IsNaN_8U_23U_2_aelse_and_cse;
  wire and_4164_cse;
  wire and_4165_cse;
  wire and_4159_cse;
  wire and_4160_cse;
  wire nor_1877_cse;
  wire and_4154_cse;
  wire and_4155_cse;
  wire nor_1493_cse;
  wire IsNaN_6U_10U_8_aelse_and_3_cse;
  wire IsNaN_6U_10U_8_aelse_and_cse;
  wire IsNaN_6U_10U_8_aelse_and_1_cse;
  wire IsNaN_6U_10U_8_aelse_and_2_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_31_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_33_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_and_cse;
  wire FpAdd_8U_23U_is_a_greater_oelse_and_1_cse;
  wire FpAdd_8U_23U_is_a_greater_oelse_and_3_cse;
  wire nor_1318_cse;
  wire FpMul_6U_10U_2_oelse_1_and_8_cse;
  wire FpMul_6U_10U_2_oelse_1_and_9_cse;
  wire FpMul_6U_10U_2_oelse_1_and_10_cse;
  wire FpMul_6U_10U_2_oelse_1_and_11_cse;
  wire FpMul_6U_10U_1_oelse_1_and_5_cse;
  wire FpMul_6U_10U_1_oelse_1_and_7_cse;
  wire FpMul_6U_10U_1_oelse_1_and_9_cse;
  wire IsNaN_8U_23U_3_aelse_and_cse;
  wire IsNaN_8U_23U_3_aelse_and_1_cse;
  wire IsNaN_8U_23U_3_aelse_and_2_cse;
  wire IsNaN_8U_23U_3_aelse_and_3_cse;
  wire and_3880_cse;
  wire mux_615_cse;
  wire nor_1490_cse;
  wire nor_1488_cse;
  wire mux_635_cse;
  wire mux_645_cse;
  wire nor_1469_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_39_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_41_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_43_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_45_cse;
  wire and_4145_cse;
  wire IsZero_6U_10U_9_and_cse;
  wire IsZero_6U_10U_9_and_1_cse;
  wire IsZero_6U_10U_9_and_2_cse;
  wire IsZero_6U_10U_9_and_3_cse;
  wire IsNaN_6U_10U_2_aelse_and_12_cse;
  wire IsNaN_6U_10U_2_aelse_and_13_cse;
  wire IsNaN_6U_10U_2_aelse_and_14_cse;
  wire IsNaN_6U_10U_2_aelse_and_15_cse;
  wire IsNaN_8U_23U_3_aelse_and_7_cse;
  wire IsNaN_8U_23U_3_aelse_and_6_cse;
  wire IsNaN_8U_23U_3_aelse_and_5_cse;
  wire IsNaN_8U_23U_3_aelse_and_4_cse;
  wire or_6042_cse;
  wire and_4178_cse;
  wire and_4177_cse;
  wire and_4176_cse;
  wire and_4175_cse;
  wire nor_1336_cse_1;
  wire nor_1697_cse;
  wire mux_93_cse;
  wire nor_1913_cse;
  wire nand_326_cse;
  wire nor_758_cse;
  wire nor_756_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_5_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_6_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_7_cse;
  wire FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_8_cse;
  reg reg_inp_lookup_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse;
  reg reg_inp_lookup_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse;
  reg reg_inp_lookup_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse;
  reg reg_inp_lookup_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse;
  wire nand_772_cse;
  wire nand_774_cse;
  wire nand_773_cse;
  wire nor_1883_cse;
  wire nand_332_cse;
  wire or_1621_cse;
  wire or_1632_cse;
  wire or_1645_cse;
  wire or_1658_cse;
  wire IsNaN_6U_10U_7_aelse_and_4_cse;
  wire mux_1963_cse;
  wire IntShiftRight_69U_6U_32U_obits_fixed_inp_lookup_else_or_7_cse;
  wire nor_623_cse;
  wire mux_461_cse;
  wire mux_854_cse;
  wire IsNaN_6U_10U_2_aelse_and_30_cse;
  wire mux_1541_cse;
  wire or_5152_cse;
  wire mux_1476_cse;
  wire mux_1483_cse;
  wire or_5154_cse;
  wire or_5155_cse;
  wire and_3286_cse;
  wire and_3285_cse;
  wire and_307_cse;
  wire and_312_cse;
  wire and_152_cse;
  wire and_144_cse;
  wire and_137_cse;
  wire and_131_cse;
  wire and_3169_cse;
  wire and_3283_cse;
  wire and_3281_cse;
  wire and_310_cse;
  wire and_4210_cse;
  wire cfg_precision_and_32_cse;
  wire cfg_precision_and_35_cse;
  wire cfg_precision_and_33_cse;
  wire cfg_precision_and_34_cse;
  wire nor_962_itm;
  wire [22:0] FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_4_itm;
  wire [22:0] FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_5_itm;
  wire [22:0] FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_7_itm;
  wire [9:0] FpMul_6U_10U_2_FpMul_6U_10U_2_FpMul_6U_10U_2_nor_5_itm;
  wire [22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_4_itm;
  wire [22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_5_itm;
  wire [22:0] FpAdd_8U_23U_FpAdd_8U_23U_or_6_itm;
  wire inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_itm_5;
  wire inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_itm_5;
  wire inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_itm_5;
  wire inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_itm_5;
  wire inp_lookup_1_FpMul_6U_10U_2_else_2_if_acc_itm_6;
  wire inp_lookup_1_FpMul_6U_10U_2_oelse_1_acc_itm_7;
  wire inp_lookup_2_FpMul_6U_10U_2_else_2_if_acc_itm_6;
  wire inp_lookup_2_FpMul_6U_10U_2_oelse_1_acc_itm_7;
  wire inp_lookup_3_FpMul_6U_10U_2_else_2_if_acc_itm_6_1;
  wire inp_lookup_4_FpMul_6U_10U_2_else_2_if_acc_itm_6;
  wire inp_lookup_4_FpMul_6U_10U_2_oelse_1_acc_itm_7;
  wire inp_lookup_1_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1;
  wire inp_lookup_1_FpMul_6U_10U_1_else_2_if_acc_itm_6_1;
  wire inp_lookup_1_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1;
  wire inp_lookup_2_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1;
  wire inp_lookup_2_FpMul_6U_10U_1_else_2_if_acc_itm_6_1;
  wire inp_lookup_2_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1;
  wire inp_lookup_3_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1;
  wire inp_lookup_3_FpMul_6U_10U_1_else_2_if_acc_itm_6_1;
  wire inp_lookup_3_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1;
  wire inp_lookup_4_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1;
  wire inp_lookup_4_FpMul_6U_10U_1_else_2_if_acc_itm_6_1;
  wire inp_lookup_4_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1;
  wire inp_lookup_1_FpMul_6U_10U_1_else_2_else_if_if_acc_1_itm_5_1;
  wire inp_lookup_2_FpMul_6U_10U_1_else_2_else_if_if_acc_1_itm_5_1;
  wire inp_lookup_3_FpMul_6U_10U_1_else_2_else_if_if_acc_1_itm_5_1;
  wire inp_lookup_4_FpMul_6U_10U_1_else_2_else_if_if_acc_1_itm_5_1;
  wire inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8;
  wire inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7;
  wire inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8;
  wire inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8;
  wire inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7;
  wire inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8;
  wire inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8;
  wire inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7;
  wire inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8;
  wire inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8;
  wire inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7;
  wire inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8;
  wire inp_lookup_1_FpMul_6U_10U_else_2_if_acc_itm_6_1;
  wire inp_lookup_2_FpMul_6U_10U_else_2_if_acc_itm_6_1;
  wire inp_lookup_3_FpMul_6U_10U_else_2_if_acc_itm_6_1;
  wire inp_lookup_4_FpMul_6U_10U_else_2_if_acc_itm_6_1;
  wire FpAdd_6U_10U_is_a_greater_acc_itm_6_1;
  wire FpAdd_6U_10U_is_a_greater_acc_1_itm_6_1;
  wire FpAdd_6U_10U_is_a_greater_acc_2_itm_6_1;
  wire FpAdd_6U_10U_is_a_greater_acc_3_itm_6_1;
  wire inp_lookup_1_FpAdd_6U_10U_if_3_if_acc_1_itm_5;
  wire inp_lookup_2_FpAdd_6U_10U_if_3_if_acc_1_itm_5;
  wire inp_lookup_3_FpAdd_6U_10U_if_3_if_acc_1_itm_5;
  wire inp_lookup_4_FpAdd_6U_10U_if_3_if_acc_1_itm_5;
  wire FpAdd_6U_10U_1_is_a_greater_acc_3_itm_6_1;
  wire FpAdd_6U_10U_1_is_a_greater_acc_2_itm_6;
  wire FpAdd_6U_10U_1_is_a_greater_acc_1_itm_6;
  wire FpAdd_6U_10U_1_is_a_greater_acc_itm_6;
  wire inp_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_1_itm_7_1;
  wire inp_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_1_itm_7;
  wire inp_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_1_itm_7_1;
  wire inp_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_1_itm_7_1;
  wire inp_lookup_1_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_itm_5_1;
  wire inp_lookup_2_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_itm_5_1;
  wire inp_lookup_3_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_itm_5_1;
  wire inp_lookup_4_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_itm_5_1;
  wire inp_lookup_1_FpMul_6U_10U_1_oelse_1_acc_itm_7_1;
  wire inp_lookup_2_FpMul_6U_10U_1_oelse_1_acc_itm_7_1;
  wire inp_lookup_3_FpMul_6U_10U_1_oelse_1_acc_itm_7_1;
  wire inp_lookup_4_FpMul_6U_10U_1_oelse_1_acc_itm_7_1;
  wire inp_lookup_1_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1;
  wire FpAdd_8U_23U_1_is_a_greater_acc_itm_8_1;
  wire inp_lookup_1_IntSaturation_51U_32U_if_acc_itm_2_1;
  wire inp_lookup_2_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1;
  wire FpAdd_8U_23U_1_is_a_greater_acc_1_itm_8_1;
  wire inp_lookup_2_IntSaturation_51U_32U_if_acc_itm_2_1;
  wire inp_lookup_3_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1;
  wire FpAdd_8U_23U_1_is_a_greater_acc_2_itm_8_1;
  wire inp_lookup_3_IntSaturation_51U_32U_if_acc_itm_2_1;
  wire inp_lookup_4_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1;
  wire FpAdd_8U_23U_1_is_a_greater_acc_3_itm_8_1;
  wire inp_lookup_4_IntSaturation_51U_32U_if_acc_itm_2_1;
  wire inp_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_1_itm_7_1;
  wire FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_itm_10;
  wire inp_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_1_itm_7_1;
  wire FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_1_itm_10;
  wire inp_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_1_itm_7;
  wire FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_2_itm_10;
  wire inp_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_1_itm_7_1;
  wire FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_3_itm_10;
  wire inp_lookup_1_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1;
  wire inp_lookup_2_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1;
  wire inp_lookup_3_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1;
  wire inp_lookup_4_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1;
  wire inp_lookup_1_FpMul_6U_10U_oelse_1_acc_itm_7_1;
  wire inp_lookup_2_FpMul_6U_10U_oelse_1_acc_itm_7_1;
  wire inp_lookup_3_FpMul_6U_10U_oelse_1_acc_itm_7_1;
  wire inp_lookup_4_FpMul_6U_10U_oelse_1_acc_itm_7_1;
  wire inp_lookup_1_FpMul_6U_10U_else_2_else_if_if_acc_1_itm_5_1;
  wire inp_lookup_2_FpMul_6U_10U_else_2_else_if_if_acc_1_itm_5_1;
  wire inp_lookup_3_FpMul_6U_10U_else_2_else_if_if_acc_1_itm_5_1;
  wire inp_lookup_4_FpMul_6U_10U_else_2_else_if_if_acc_1_itm_5_1;
  wire inp_lookup_1_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1;
  wire inp_lookup_2_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1;
  wire inp_lookup_3_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1;
  wire inp_lookup_4_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1;
  wire inp_lookup_1_IntSaturation_51U_32U_else_if_acc_itm_2_1;
  wire inp_lookup_2_IntSaturation_51U_32U_else_if_acc_itm_2_1;
  wire inp_lookup_3_IntSaturation_51U_32U_else_if_acc_itm_2_1;
  wire inp_lookup_4_IntSaturation_51U_32U_else_if_acc_itm_2_1;
  wire FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_itm_23_1;
  wire FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_1_itm_23_1;
  wire FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_2_itm_23_1;
  wire FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_3_itm_23_1;
  wire FpAdd_6U_10U_is_a_greater_oif_aelse_acc_itm_10_1;
  wire FpAdd_6U_10U_is_a_greater_oif_aelse_acc_1_itm_10_1;
  wire FpAdd_6U_10U_is_a_greater_oif_aelse_acc_2_itm_10_1;
  wire FpAdd_6U_10U_is_a_greater_oif_aelse_acc_3_itm_10_1;
  wire or_tmp_4811;
  wire or_tmp_4815;
  wire mux_tmp;
  wire not_tmp_3015;
  wire or_tmp_4829;
  wire or_tmp_4830;
  wire mux_tmp_2075;
  wire or_tmp_4831;
  wire or_tmp_4843;
  wire or_tmp_4845;
  wire or_tmp_4846;
  wire mux_tmp_2091;
  wire or_6231_cse;
  wire or_6230_cse;
  wire or_6229_cse;
  wire nor_1961_cse;
  wire or_6241_cse;
  wire nand_728_cse_1;
  wire or_6252_cse;
  wire or_6257_cse;
  wire nand_598_cse;
  wire nor_1967_cse;
  wire or_6272_cse;
  wire nor_1978_cse;
  wire or_4340_cse;
  wire[0:0] shift_0_prb;
  wire[0:0] and_44;
  wire[0:0] shift_0_prb_1;
  wire[0:0] and_51;
  wire[0:0] shift_0_prb_2;
  wire[0:0] and_58;
  wire[0:0] shift_0_prb_3;
  wire[0:0] and_65;
  wire[0:0] iMantWidth_oMantWidth_prb;
  wire[0:0] iExpoWidth_oExpoWidth_prb;
  wire[0:0] iExpoWidth_oExpoWidth_prb_1;
  wire[0:0] iMantWidth_oMantWidth_prb_1;
  wire[0:0] iExpoWidth_oExpoWidth_prb_2;
  wire[0:0] iExpoWidth_oExpoWidth_prb_3;
  wire[0:0] iMantWidth_oMantWidth_prb_2;
  wire[0:0] iMantWidth_oMantWidth_prb_3;
  wire[0:0] iExpoWidth_oExpoWidth_prb_4;
  wire[0:0] oWidth_iWidth_prb;
  wire[0:0] or_4171;
  wire[0:0] iExpoWidth_oExpoWidth_prb_5;
  wire[0:0] iExpoWidth_oExpoWidth_prb_6;
  wire[0:0] iMantWidth_oMantWidth_prb_4;
  wire[0:0] iMantWidth_oMantWidth_prb_5;
  wire[0:0] iExpoWidth_oExpoWidth_prb_7;
  wire[0:0] iMantWidth_oMantWidth_prb_6;
  wire[0:0] iMantWidth_oMantWidth_prb_7;
  wire[0:0] iExpoWidth_oExpoWidth_prb_8;
  wire[0:0] iMantWidth_oMantWidth_prb_8;
  wire[0:0] iExpoWidth_oExpoWidth_prb_9;
  wire[0:0] iExpoWidth_oExpoWidth_prb_10;
  wire[0:0] iMantWidth_oMantWidth_prb_9;
  wire[0:0] iExpoWidth_oExpoWidth_prb_11;
  wire[0:0] iExpoWidth_oExpoWidth_prb_12;
  wire[0:0] iMantWidth_oMantWidth_prb_10;
  wire[0:0] iMantWidth_oMantWidth_prb_11;
  wire[0:0] iExpoWidth_oExpoWidth_prb_13;
  wire[0:0] oWidth_iWidth_prb_1;
  wire[0:0] or_4174;
  wire[0:0] iExpoWidth_oExpoWidth_prb_14;
  wire[0:0] iExpoWidth_oExpoWidth_prb_15;
  wire[0:0] iMantWidth_oMantWidth_prb_12;
  wire[0:0] iMantWidth_oMantWidth_prb_13;
  wire[0:0] iExpoWidth_oExpoWidth_prb_16;
  wire[0:0] iMantWidth_oMantWidth_prb_14;
  wire[0:0] iMantWidth_oMantWidth_prb_15;
  wire[0:0] iExpoWidth_oExpoWidth_prb_17;
  wire[0:0] iMantWidth_oMantWidth_prb_16;
  wire[0:0] iExpoWidth_oExpoWidth_prb_18;
  wire[0:0] iExpoWidth_oExpoWidth_prb_19;
  wire[0:0] iMantWidth_oMantWidth_prb_17;
  wire[0:0] iExpoWidth_oExpoWidth_prb_20;
  wire[0:0] iExpoWidth_oExpoWidth_prb_21;
  wire[0:0] iMantWidth_oMantWidth_prb_18;
  wire[0:0] iMantWidth_oMantWidth_prb_19;
  wire[0:0] iExpoWidth_oExpoWidth_prb_22;
  wire[0:0] oWidth_iWidth_prb_2;
  wire[0:0] or_4177;
  wire[0:0] iExpoWidth_oExpoWidth_prb_23;
  wire[0:0] iExpoWidth_oExpoWidth_prb_24;
  wire[0:0] iMantWidth_oMantWidth_prb_20;
  wire[0:0] iMantWidth_oMantWidth_prb_21;
  wire[0:0] iExpoWidth_oExpoWidth_prb_25;
  wire[0:0] iMantWidth_oMantWidth_prb_22;
  wire[0:0] iMantWidth_oMantWidth_prb_23;
  wire[0:0] iExpoWidth_oExpoWidth_prb_26;
  wire[0:0] iMantWidth_oMantWidth_prb_24;
  wire[0:0] iExpoWidth_oExpoWidth_prb_27;
  wire[0:0] iExpoWidth_oExpoWidth_prb_28;
  wire[0:0] iMantWidth_oMantWidth_prb_25;
  wire[0:0] iExpoWidth_oExpoWidth_prb_29;
  wire[0:0] iExpoWidth_oExpoWidth_prb_30;
  wire[0:0] iMantWidth_oMantWidth_prb_26;
  wire[0:0] iMantWidth_oMantWidth_prb_27;
  wire[0:0] iExpoWidth_oExpoWidth_prb_31;
  wire[0:0] oWidth_iWidth_prb_3;
  wire[0:0] or_4180;
  wire[0:0] iExpoWidth_oExpoWidth_prb_32;
  wire[0:0] iExpoWidth_oExpoWidth_prb_33;
  wire[0:0] iMantWidth_oMantWidth_prb_28;
  wire[0:0] iMantWidth_oMantWidth_prb_29;
  wire[0:0] iExpoWidth_oExpoWidth_prb_34;
  wire[0:0] iMantWidth_oMantWidth_prb_30;
  wire[0:0] iMantWidth_oMantWidth_prb_31;
  wire[0:0] iExpoWidth_oExpoWidth_prb_35;
  wire[3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_4_nl;
  wire[3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_mux_5_nl;
  wire[0:0] FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_20_nl;
  wire[3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_9_nl;
  wire[3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_mux_18_nl;
  wire[0:0] FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_21_nl;
  wire[3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_14_nl;
  wire[3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_mux_31_nl;
  wire[0:0] FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_22_nl;
  wire[3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_19_nl;
  wire[3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_mux_44_nl;
  wire[0:0] FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_23_nl;
  wire[0:0] inp_lookup_if_mux_600_nl;
  wire[0:0] nor_1802_nl;
  wire[0:0] FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_4_nl;
  wire[0:0] inp_lookup_or_nl;
  wire[0:0] inp_lookup_and_82_nl;
  wire[2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_3_nl;
  wire[2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_nl;
  wire[2:0] inp_lookup_1_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl;
  wire[3:0] nl_inp_lookup_1_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl;
  wire[0:0] IsZero_6U_23U_aelse_IsZero_6U_23U_or_3_nl;
  wire[0:0] inp_lookup_if_mux_601_nl;
  wire[0:0] nor_1803_nl;
  wire[0:0] FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_9_nl;
  wire[0:0] inp_lookup_or_1_nl;
  wire[0:0] inp_lookup_and_86_nl;
  wire[2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_8_nl;
  wire[2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_5_nl;
  wire[2:0] inp_lookup_2_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl;
  wire[3:0] nl_inp_lookup_2_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl;
  wire[0:0] IsZero_6U_23U_aelse_IsZero_6U_23U_or_2_nl;
  wire[0:0] inp_lookup_if_mux_602_nl;
  wire[0:0] nor_1804_nl;
  wire[0:0] FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_14_nl;
  wire[0:0] inp_lookup_or_2_nl;
  wire[0:0] inp_lookup_and_90_nl;
  wire[2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_13_nl;
  wire[2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_10_nl;
  wire[2:0] inp_lookup_3_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl;
  wire[3:0] nl_inp_lookup_3_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl;
  wire[0:0] IsZero_6U_23U_aelse_IsZero_6U_23U_or_1_nl;
  wire[0:0] inp_lookup_if_mux_603_nl;
  wire[0:0] nor_1805_nl;
  wire[0:0] FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_19_nl;
  wire[0:0] inp_lookup_or_3_nl;
  wire[0:0] inp_lookup_and_94_nl;
  wire[2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_18_nl;
  wire[2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_15_nl;
  wire[2:0] inp_lookup_4_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl;
  wire[3:0] nl_inp_lookup_4_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl;
  wire[0:0] IsZero_6U_23U_aelse_IsZero_6U_23U_or_nl;
  wire[0:0] mux_78_nl;
  wire[0:0] mux_80_nl;
  wire[0:0] nor_1721_nl;
  wire[0:0] nor_1722_nl;
  wire[0:0] inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_nl;
  wire[0:0] IsZero_6U_10U_7_IsZero_6U_10U_7_and_nl;
  wire[9:0] FpFractionToFloat_35U_6U_10U_1_if_else_else_FpFractionToFloat_35U_6U_10U_1_if_else_else_and_nl;
  wire[0:0] FpFractionToFloat_35U_6U_10U_1_o_mant_and_nl;
  wire[0:0] FpFractionToFloat_35U_6U_10U_1_o_mant_and_10_nl;
  wire[0:0] mux_86_nl;
  wire[0:0] nor_1717_nl;
  wire[0:0] nor_1718_nl;
  wire[0:0] inp_lookup_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_nl;
  wire[0:0] IsZero_6U_10U_7_IsZero_6U_10U_7_and_1_nl;
  wire[0:0] mux_92_nl;
  wire[0:0] nand_nl;
  wire[9:0] FpFractionToFloat_35U_6U_10U_1_if_else_else_FpFractionToFloat_35U_6U_10U_1_if_else_else_and_1_nl;
  wire[0:0] FpFractionToFloat_35U_6U_10U_1_o_mant_and_8_nl;
  wire[0:0] FpFractionToFloat_35U_6U_10U_1_o_mant_and_9_nl;
  wire[0:0] mux_94_nl;
  wire[0:0] nor_1715_nl;
  wire[0:0] nor_1716_nl;
  wire[0:0] inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_nl;
  wire[0:0] IsZero_6U_10U_7_IsZero_6U_10U_7_and_2_nl;
  wire[9:0] FpFractionToFloat_35U_6U_10U_1_if_else_else_FpFractionToFloat_35U_6U_10U_1_if_else_else_and_2_nl;
  wire[0:0] FpFractionToFloat_35U_6U_10U_1_o_mant_and_6_nl;
  wire[0:0] FpFractionToFloat_35U_6U_10U_1_o_mant_and_7_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_FpAdd_8U_23U_is_a_greater_or_3_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_nl;
  wire[8:0] FpAdd_8U_23U_is_a_greater_acc_3_nl;
  wire[10:0] nl_FpAdd_8U_23U_is_a_greater_acc_3_nl;
  wire[0:0] mux_99_nl;
  wire[0:0] nor_1760_nl;
  wire[0:0] nor_1761_nl;
  wire[0:0] inp_lookup_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_nl;
  wire[0:0] IsZero_6U_10U_7_IsZero_6U_10U_7_and_3_nl;
  wire[0:0] mux_105_nl;
  wire[0:0] mux_104_nl;
  wire[0:0] nand_2_nl;
  wire[9:0] FpFractionToFloat_35U_6U_10U_1_if_else_else_FpFractionToFloat_35U_6U_10U_1_if_else_else_and_3_nl;
  wire[0:0] FpFractionToFloat_35U_6U_10U_1_o_mant_and_4_nl;
  wire[0:0] FpFractionToFloat_35U_6U_10U_1_o_mant_and_5_nl;
  wire[0:0] mux_108_nl;
  wire[0:0] mux_110_nl;
  wire[9:0] FpFractionToFloat_35U_6U_10U_if_else_else_FpFractionToFloat_35U_6U_10U_if_else_else_and_nl;
  wire[0:0] mux_111_nl;
  wire[0:0] nor_1707_nl;
  wire[0:0] nor_1708_nl;
  wire[0:0] mux_114_nl;
  wire[0:0] nor_1703_nl;
  wire[0:0] mux_112_nl;
  wire[0:0] or_156_nl;
  wire[0:0] mux_113_nl;
  wire[0:0] nor_1704_nl;
  wire[0:0] mux_116_nl;
  wire[0:0] mux_119_nl;
  wire[0:0] and_3369_nl;
  wire[0:0] nor_1700_nl;
  wire[7:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_asn_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_conc_40_cgspt_7_mux_nl;
  wire[0:0] mux_1866_nl;
  wire[0:0] mux_2045_nl;
  wire[0:0] mux_2043_nl;
  wire[0:0] nor_1893_nl;
  wire[0:0] mux_2044_nl;
  wire[0:0] nor_1894_nl;
  wire[0:0] mux_2047_nl;
  wire[0:0] mux_2046_nl;
  wire[0:0] and_4147_nl;
  wire[0:0] and_4148_nl;
  wire[4:0] FpFractionToFloat_35U_6U_10U_nor_nl;
  wire[4:0] FpFractionToFloat_35U_6U_10U_if_else_mux_nl;
  wire[4:0] inp_lookup_1_FpFractionToFloat_35U_6U_10U_if_else_else_else_acc_nl;
  wire[5:0] nl_inp_lookup_1_FpFractionToFloat_35U_6U_10U_if_else_else_else_acc_nl;
  wire[0:0] mux_127_nl;
  wire[0:0] mux_126_nl;
  wire[0:0] or_205_nl;
  wire[0:0] or_208_nl;
  wire[0:0] mux_129_nl;
  wire[0:0] mux_133_nl;
  wire[9:0] FpFractionToFloat_35U_6U_10U_if_else_else_FpFractionToFloat_35U_6U_10U_if_else_else_and_1_nl;
  wire[0:0] mux_134_nl;
  wire[0:0] nor_1690_nl;
  wire[0:0] nor_1691_nl;
  wire[0:0] mux_137_nl;
  wire[0:0] nor_1686_nl;
  wire[0:0] mux_135_nl;
  wire[0:0] or_226_nl;
  wire[0:0] mux_136_nl;
  wire[0:0] nor_1687_nl;
  wire[0:0] mux_139_nl;
  wire[0:0] mux_142_nl;
  wire[0:0] nor_1682_nl;
  wire[0:0] mux_141_nl;
  wire[0:0] nor_1683_nl;
  wire[0:0] nor_1684_nl;
  wire[7:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_asn_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_conc_41_cgspt_7_mux_nl;
  wire[0:0] mux_1867_nl;
  wire[0:0] mux_2050_nl;
  wire[0:0] mux_2049_nl;
  wire[0:0] mux_2048_nl;
  wire[0:0] nor_1889_nl;
  wire[0:0] nor_1890_nl;
  wire[0:0] and_4146_nl;
  wire[0:0] mux_2051_nl;
  wire[0:0] and_3610_nl;
  wire[4:0] FpFractionToFloat_35U_6U_10U_nor_1_nl;
  wire[4:0] FpFractionToFloat_35U_6U_10U_if_else_mux_16_nl;
  wire[4:0] inp_lookup_2_FpFractionToFloat_35U_6U_10U_if_else_else_else_acc_nl;
  wire[5:0] nl_inp_lookup_2_FpFractionToFloat_35U_6U_10U_if_else_else_else_acc_nl;
  wire[0:0] mux_149_nl;
  wire[0:0] mux_148_nl;
  wire[0:0] or_269_nl;
  wire[0:0] or_272_nl;
  wire[0:0] mux_151_nl;
  wire[0:0] mux_155_nl;
  wire[9:0] FpFractionToFloat_35U_6U_10U_if_else_else_FpFractionToFloat_35U_6U_10U_if_else_else_and_2_nl;
  wire[0:0] mux_156_nl;
  wire[0:0] nor_1671_nl;
  wire[0:0] nor_1672_nl;
  wire[0:0] mux_159_nl;
  wire[0:0] mux_157_nl;
  wire[0:0] nor_1665_nl;
  wire[0:0] mux_158_nl;
  wire[0:0] nor_1668_nl;
  wire[0:0] mux_161_nl;
  wire[0:0] mux_164_nl;
  wire[0:0] and_3364_nl;
  wire[0:0] nor_1662_nl;
  wire[0:0] mux_165_nl;
  wire[0:0] nor_1661_nl;
  wire[0:0] and_3363_nl;
  wire[4:0] FpFractionToFloat_35U_6U_10U_nor_2_nl;
  wire[4:0] FpFractionToFloat_35U_6U_10U_if_else_mux_17_nl;
  wire[4:0] inp_lookup_3_FpFractionToFloat_35U_6U_10U_if_else_else_else_acc_nl;
  wire[5:0] nl_inp_lookup_3_FpFractionToFloat_35U_6U_10U_if_else_else_else_acc_nl;
  wire[0:0] mux_169_nl;
  wire[0:0] mux_168_nl;
  wire[0:0] or_339_nl;
  wire[0:0] or_342_nl;
  wire[0:0] mux_170_nl;
  wire[0:0] mux_174_nl;
  wire[9:0] FpFractionToFloat_35U_6U_10U_if_else_else_FpFractionToFloat_35U_6U_10U_if_else_else_and_3_nl;
  wire[0:0] mux_175_nl;
  wire[0:0] nor_1656_nl;
  wire[0:0] nor_1658_nl;
  wire[0:0] mux_177_nl;
  wire[0:0] nor_1654_nl;
  wire[0:0] mux_176_nl;
  wire[0:0] or_360_nl;
  wire[0:0] nor_1655_nl;
  wire[0:0] mux_179_nl;
  wire[0:0] mux_182_nl;
  wire[0:0] mux_181_nl;
  wire[0:0] nor_1650_nl;
  wire[0:0] and_3388_nl;
  wire[0:0] nor_1652_nl;
  wire[7:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_asn_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_conc_42_cgspt_7_mux_nl;
  wire[0:0] mux_1868_nl;
  wire[0:0] mux_2053_nl;
  wire[0:0] mux_2052_nl;
  wire[0:0] and_4143_nl;
  wire[0:0] and_4144_nl;
  wire[0:0] mux_2054_nl;
  wire[0:0] and_3622_nl;
  wire[4:0] FpFractionToFloat_35U_6U_10U_nor_3_nl;
  wire[4:0] FpFractionToFloat_35U_6U_10U_if_else_mux_18_nl;
  wire[4:0] inp_lookup_4_FpFractionToFloat_35U_6U_10U_if_else_else_else_acc_nl;
  wire[5:0] nl_inp_lookup_4_FpFractionToFloat_35U_6U_10U_if_else_else_else_acc_nl;
  wire[0:0] mux_187_nl;
  wire[0:0] nor_1644_nl;
  wire[0:0] nor_1645_nl;
  wire[0:0] mux_189_nl;
  wire[0:0] nor_1641_nl;
  wire[0:0] mux_188_nl;
  wire[0:0] nor_1642_nl;
  wire[0:0] nor_1643_nl;
  wire[0:0] mux_190_nl;
  wire[0:0] mux_1870_nl;
  wire[22:0] and_3421_nl;
  wire[0:0] FpAdd_8U_23U_o_mant_not_nl;
  wire[0:0] and_894_nl;
  wire[0:0] mux_2225_nl;
  wire[0:0] mux_2223_nl;
  wire[0:0] mux_2218_nl;
  wire[0:0] mux_2213_nl;
  wire[0:0] mux_2210_nl;
  wire[0:0] mux_2212_nl;
  wire[0:0] mux_2211_nl;
  wire[0:0] nor_1977_nl;
  wire[0:0] and_4228_nl;
  wire[0:0] mux_2217_nl;
  wire[0:0] mux_2214_nl;
  wire[0:0] mux_2216_nl;
  wire[0:0] mux_2215_nl;
  wire[0:0] and_4237_nl;
  wire[0:0] mux_2222_nl;
  wire[0:0] and_4229_nl;
  wire[0:0] mux_2221_nl;
  wire[0:0] mux_2219_nl;
  wire[0:0] or_6247_nl;
  wire[0:0] mux_2220_nl;
  wire[0:0] or_6249_nl;
  wire[0:0] mux_2224_nl;
  wire[0:0] or_6250_nl;
  wire[0:0] mux_196_nl;
  wire[0:0] nand_684_nl;
  wire[7:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_nl;
  wire[7:0] inp_lookup_1_FpNormalize_8U_49U_else_acc_nl;
  wire[9:0] nl_inp_lookup_1_FpNormalize_8U_49U_else_acc_nl;
  wire[0:0] FpNormalize_8U_49U_oelse_not_4_nl;
  wire[7:0] inp_lookup_1_FpAdd_8U_23U_if_3_if_acc_nl;
  wire[8:0] nl_inp_lookup_1_FpAdd_8U_23U_if_3_if_acc_nl;
  wire[0:0] mux_200_nl;
  wire[0:0] or_433_nl;
  wire[0:0] mux_191_nl;
  wire[0:0] or_5922_nl;
  wire[0:0] or_436_nl;
  wire[0:0] mux_2057_nl;
  wire[0:0] or_5925_nl;
  wire[0:0] mux_201_nl;
  wire[0:0] and_3359_nl;
  wire[0:0] and_3360_nl;
  wire[0:0] mux_202_nl;
  wire[29:0] inp_lookup_1_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_nl;
  wire[0:0] inp_lookup_1_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_nl;
  wire[0:0] mux_208_nl;
  wire[0:0] mux_207_nl;
  wire[0:0] mux_206_nl;
  wire[0:0] mux_213_nl;
  wire[0:0] mux_212_nl;
  wire[0:0] or_456_nl;
  wire[0:0] mux_224_nl;
  wire[0:0] mux_219_nl;
  wire[0:0] mux_218_nl;
  wire[0:0] mux_217_nl;
  wire[0:0] mux_216_nl;
  wire[0:0] nor_1639_nl;
  wire[0:0] and_3356_nl;
  wire[0:0] mux_223_nl;
  wire[0:0] mux_221_nl;
  wire[0:0] mux_220_nl;
  wire[0:0] or_468_nl;
  wire[0:0] mux_222_nl;
  wire[0:0] nand_15_nl;
  wire[0:0] mux_226_nl;
  wire[0:0] mux_225_nl;
  wire[0:0] or_474_nl;
  wire[0:0] or_476_nl;
  wire[0:0] mux_228_nl;
  wire[0:0] or_478_nl;
  wire[0:0] mux_227_nl;
  wire[0:0] or_481_nl;
  wire[0:0] mux_230_nl;
  wire[0:0] or_483_nl;
  wire[0:0] mux_229_nl;
  wire[0:0] or_485_nl;
  wire[0:0] or_482_nl;
  wire[0:0] mux_1874_nl;
  wire[0:0] or_4352_nl;
  wire[22:0] and_3422_nl;
  wire[0:0] FpAdd_8U_23U_o_mant_not_1_nl;
  wire[0:0] and_931_nl;
  wire[0:0] mux_2241_nl;
  wire[0:0] mux_2239_nl;
  wire[0:0] mux_2235_nl;
  wire[0:0] mux_2230_nl;
  wire[0:0] mux_2227_nl;
  wire[0:0] mux_2229_nl;
  wire[0:0] mux_2228_nl;
  wire[0:0] nor_1976_nl;
  wire[0:0] and_4231_nl;
  wire[0:0] mux_2234_nl;
  wire[0:0] mux_2231_nl;
  wire[0:0] mux_2233_nl;
  wire[0:0] mux_2232_nl;
  wire[0:0] and_4239_nl;
  wire[0:0] mux_2238_nl;
  wire[0:0] and_4232_nl;
  wire[0:0] mux_2237_nl;
  wire[0:0] and_4240_nl;
  wire[0:0] mux_2236_nl;
  wire[0:0] or_6265_nl;
  wire[0:0] mux_2240_nl;
  wire[0:0] or_6266_nl;
  wire[0:0] mux_236_nl;
  wire[0:0] nand_599_nl;
  wire[7:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_2_nl;
  wire[7:0] inp_lookup_2_FpNormalize_8U_49U_else_acc_nl;
  wire[9:0] nl_inp_lookup_2_FpNormalize_8U_49U_else_acc_nl;
  wire[0:0] FpNormalize_8U_49U_oelse_not_5_nl;
  wire[7:0] inp_lookup_2_FpAdd_8U_23U_if_3_if_acc_nl;
  wire[8:0] nl_inp_lookup_2_FpAdd_8U_23U_if_3_if_acc_nl;
  wire[0:0] mux_238_nl;
  wire[0:0] or_498_nl;
  wire[0:0] mux_231_nl;
  wire[0:0] or_5933_nl;
  wire[0:0] or_499_nl;
  wire[0:0] mux_2062_nl;
  wire[0:0] mux_239_nl;
  wire[29:0] inp_lookup_2_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_nl;
  wire[0:0] inp_lookup_2_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_nl;
  wire[0:0] mux_246_nl;
  wire[0:0] mux_245_nl;
  wire[0:0] mux_244_nl;
  wire[0:0] mux_251_nl;
  wire[0:0] mux_250_nl;
  wire[0:0] or_518_nl;
  wire[0:0] mux_263_nl;
  wire[0:0] mux_257_nl;
  wire[0:0] mux_256_nl;
  wire[0:0] mux_255_nl;
  wire[0:0] mux_254_nl;
  wire[0:0] nor_1637_nl;
  wire[0:0] and_3352_nl;
  wire[0:0] mux_262_nl;
  wire[0:0] mux_259_nl;
  wire[0:0] mux_258_nl;
  wire[0:0] or_530_nl;
  wire[0:0] mux_261_nl;
  wire[0:0] mux_260_nl;
  wire[0:0] nor_1638_nl;
  wire[0:0] or_531_nl;
  wire[0:0] mux_264_nl;
  wire[0:0] or_535_nl;
  wire[0:0] mux_265_nl;
  wire[0:0] nor_1959_nl;
  wire[0:0] nor_1960_nl;
  wire[0:0] mux_267_nl;
  wire[0:0] or_539_nl;
  wire[0:0] mux_266_nl;
  wire[0:0] or_541_nl;
  wire[0:0] or_538_nl;
  wire[0:0] mux_1880_nl;
  wire[0:0] or_4363_nl;
  wire[22:0] and_3423_nl;
  wire[0:0] FpAdd_8U_23U_o_mant_not_2_nl;
  wire[0:0] and_969_nl;
  wire[0:0] mux_2258_nl;
  wire[0:0] mux_2256_nl;
  wire[0:0] mux_2251_nl;
  wire[0:0] mux_2246_nl;
  wire[0:0] mux_2243_nl;
  wire[0:0] mux_2245_nl;
  wire[0:0] mux_2244_nl;
  wire[0:0] nor_1974_nl;
  wire[0:0] and_4234_nl;
  wire[0:0] mux_2250_nl;
  wire[0:0] mux_2247_nl;
  wire[0:0] mux_2249_nl;
  wire[0:0] mux_2248_nl;
  wire[0:0] and_4242_nl;
  wire[0:0] mux_2255_nl;
  wire[0:0] and_4235_nl;
  wire[0:0] mux_2254_nl;
  wire[0:0] mux_2252_nl;
  wire[0:0] or_6278_nl;
  wire[0:0] mux_2253_nl;
  wire[0:0] or_6280_nl;
  wire[0:0] mux_2257_nl;
  wire[0:0] or_6281_nl;
  wire[0:0] mux_273_nl;
  wire[0:0] nand_597_nl;
  wire[7:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_4_nl;
  wire[7:0] inp_lookup_3_FpNormalize_8U_49U_else_acc_nl;
  wire[9:0] nl_inp_lookup_3_FpNormalize_8U_49U_else_acc_nl;
  wire[0:0] FpNormalize_8U_49U_oelse_not_6_nl;
  wire[7:0] inp_lookup_3_FpAdd_8U_23U_if_3_if_acc_nl;
  wire[8:0] nl_inp_lookup_3_FpAdd_8U_23U_if_3_if_acc_nl;
  wire[0:0] mux_276_nl;
  wire[0:0] or_557_nl;
  wire[0:0] mux_275_nl;
  wire[0:0] or_560_nl;
  wire[0:0] or_563_nl;
  wire[0:0] mux_277_nl;
  wire[29:0] inp_lookup_3_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_nl;
  wire[0:0] inp_lookup_3_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_nl;
  wire[0:0] mux_284_nl;
  wire[0:0] mux_283_nl;
  wire[0:0] mux_282_nl;
  wire[0:0] mux_289_nl;
  wire[0:0] mux_288_nl;
  wire[0:0] or_579_nl;
  wire[0:0] mux_296_nl;
  wire[0:0] mux_291_nl;
  wire[0:0] mux_290_nl;
  wire[0:0] or_582_nl;
  wire[0:0] mux_295_nl;
  wire[0:0] mux_293_nl;
  wire[0:0] mux_292_nl;
  wire[0:0] nor_1634_nl;
  wire[0:0] mux_294_nl;
  wire[0:0] nor_1635_nl;
  wire[0:0] mux_308_nl;
  wire[0:0] mux_302_nl;
  wire[0:0] mux_301_nl;
  wire[0:0] mux_300_nl;
  wire[0:0] mux_299_nl;
  wire[0:0] nor_1632_nl;
  wire[0:0] and_3347_nl;
  wire[0:0] mux_307_nl;
  wire[0:0] mux_304_nl;
  wire[0:0] mux_303_nl;
  wire[0:0] mux_306_nl;
  wire[0:0] mux_305_nl;
  wire[0:0] nor_1633_nl;
  wire[0:0] or_605_nl;
  wire[0:0] mux_310_nl;
  wire[0:0] mux_309_nl;
  wire[0:0] or_609_nl;
  wire[0:0] or_610_nl;
  wire[0:0] mux_312_nl;
  wire[0:0] or_611_nl;
  wire[0:0] mux_311_nl;
  wire[0:0] or_613_nl;
  wire[0:0] mux_313_nl;
  wire[0:0] nor_1630_nl;
  wire[0:0] nor_1631_nl;
  wire[22:0] and_3424_nl;
  wire[22:0] mux_74_nl;
  wire[0:0] FpAdd_8U_23U_o_mant_not_3_nl;
  wire[0:0] and_1004_nl;
  wire[0:0] mux_314_nl;
  wire[7:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_6_nl;
  wire[7:0] inp_lookup_4_FpNormalize_8U_49U_else_acc_nl;
  wire[9:0] nl_inp_lookup_4_FpNormalize_8U_49U_else_acc_nl;
  wire[0:0] FpNormalize_8U_49U_oelse_not_7_nl;
  wire[7:0] inp_lookup_4_FpAdd_8U_23U_if_3_if_acc_nl;
  wire[8:0] nl_inp_lookup_4_FpAdd_8U_23U_if_3_if_acc_nl;
  wire[0:0] mux_319_nl;
  wire[0:0] or_625_nl;
  wire[0:0] mux_317_nl;
  wire[0:0] mux_316_nl;
  wire[0:0] or_624_nl;
  wire[0:0] or_628_nl;
  wire[0:0] mux_318_nl;
  wire[0:0] or_627_nl;
  wire[0:0] mux_320_nl;
  wire[29:0] inp_lookup_4_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_nl;
  wire[0:0] inp_lookup_4_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_nl;
  wire[0:0] mux_335_nl;
  wire[0:0] mux_334_nl;
  wire[0:0] mux_333_nl;
  wire[0:0] mux_331_nl;
  wire[0:0] mux_1992_nl;
  wire[0:0] mux_332_nl;
  wire[0:0] mux_330_nl;
  wire[0:0] or_637_nl;
  wire[0:0] mux_343_nl;
  wire[0:0] mux_342_nl;
  wire[0:0] mux_341_nl;
  wire[0:0] and_3344_nl;
  wire[0:0] mux_347_nl;
  wire[0:0] nor_1626_nl;
  wire[0:0] nor_1628_nl;
  wire[0:0] mux_348_nl;
  wire[0:0] or_663_nl;
  wire[0:0] mux_349_nl;
  wire[0:0] nor_1957_nl;
  wire[0:0] nor_1958_nl;
  wire[0:0] mux_351_nl;
  wire[0:0] and_3342_nl;
  wire[0:0] mux_350_nl;
  wire[0:0] or_667_nl;
  wire[0:0] and_3343_nl;
  wire[0:0] mux_355_nl;
  wire[0:0] and_3340_nl;
  wire[0:0] mux_352_nl;
  wire[0:0] or_671_nl;
  wire[0:0] and_3341_nl;
  wire[0:0] mux_354_nl;
  wire[0:0] or_672_nl;
  wire[0:0] mux_353_nl;
  wire[0:0] or_674_nl;
  wire[0:0] FpMul_6U_10U_1_FpMul_6U_10U_1_and_nl;
  wire[0:0] mux_367_nl;
  wire[0:0] nor_1622_nl;
  wire[0:0] nor_1623_nl;
  wire[0:0] mux_370_nl;
  wire[0:0] mux_368_nl;
  wire[0:0] or_697_nl;
  wire[0:0] mux_358_nl;
  wire[0:0] mux_357_nl;
  wire[0:0] mux_369_nl;
  wire[0:0] or_699_nl;
  wire[0:0] mux_361_nl;
  wire[0:0] or_687_nl;
  wire[0:0] mux_360_nl;
  wire[0:0] mux_380_nl;
  wire[0:0] mux_373_nl;
  wire[0:0] mux_372_nl;
  wire[0:0] mux_371_nl;
  wire[0:0] nor_1619_nl;
  wire[0:0] or_704_nl;
  wire[0:0] or_700_nl;
  wire[0:0] mux_379_nl;
  wire[0:0] mux_375_nl;
  wire[0:0] mux_374_nl;
  wire[0:0] mux_378_nl;
  wire[0:0] mux_376_nl;
  wire[0:0] mux_377_nl;
  wire[0:0] nor_1620_nl;
  wire[0:0] mux_382_nl;
  wire[0:0] and_3337_nl;
  wire[0:0] and_3338_nl;
  wire[0:0] mux_386_nl;
  wire[0:0] and_3335_nl;
  wire[0:0] mux_383_nl;
  wire[0:0] or_720_nl;
  wire[0:0] and_3336_nl;
  wire[0:0] mux_385_nl;
  wire[0:0] or_721_nl;
  wire[0:0] mux_384_nl;
  wire[0:0] or_723_nl;
  wire[0:0] FpMul_6U_10U_1_FpMul_6U_10U_1_and_16_nl;
  wire[0:0] mux_407_nl;
  wire[0:0] nor_1615_nl;
  wire[0:0] nor_1616_nl;
  wire[0:0] mux_410_nl;
  wire[0:0] mux_408_nl;
  wire[0:0] or_749_nl;
  wire[0:0] mux_401_nl;
  wire[0:0] mux_409_nl;
  wire[0:0] or_751_nl;
  wire[0:0] mux_404_nl;
  wire[0:0] or_737_nl;
  wire[0:0] mux_403_nl;
  wire[0:0] mux_420_nl;
  wire[0:0] mux_413_nl;
  wire[0:0] mux_412_nl;
  wire[0:0] mux_411_nl;
  wire[0:0] nor_1612_nl;
  wire[0:0] or_756_nl;
  wire[0:0] or_752_nl;
  wire[0:0] mux_419_nl;
  wire[0:0] mux_415_nl;
  wire[0:0] mux_414_nl;
  wire[0:0] mux_418_nl;
  wire[0:0] mux_416_nl;
  wire[0:0] mux_417_nl;
  wire[0:0] nor_1613_nl;
  wire[0:0] mux_422_nl;
  wire[0:0] and_3332_nl;
  wire[0:0] and_3333_nl;
  wire[0:0] mux_425_nl;
  wire[0:0] and_3330_nl;
  wire[0:0] mux_423_nl;
  wire[0:0] or_772_nl;
  wire[0:0] and_3331_nl;
  wire[0:0] mux_424_nl;
  wire[0:0] or_774_nl;
  wire[0:0] FpMul_6U_10U_1_FpMul_6U_10U_1_and_17_nl;
  wire[0:0] mux_439_nl;
  wire[0:0] nor_1608_nl;
  wire[0:0] nor_1609_nl;
  wire[0:0] mux_449_nl;
  wire[0:0] mux_442_nl;
  wire[0:0] mux_441_nl;
  wire[0:0] mux_440_nl;
  wire[0:0] mux_448_nl;
  wire[0:0] mux_444_nl;
  wire[0:0] mux_443_nl;
  wire[0:0] mux_447_nl;
  wire[0:0] mux_445_nl;
  wire[0:0] mux_446_nl;
  wire[0:0] nor_1606_nl;
  wire[0:0] mux_459_nl;
  wire[0:0] mux_452_nl;
  wire[0:0] mux_451_nl;
  wire[0:0] mux_450_nl;
  wire[0:0] nor_1603_nl;
  wire[0:0] or_811_nl;
  wire[0:0] mux_458_nl;
  wire[0:0] mux_454_nl;
  wire[0:0] mux_453_nl;
  wire[0:0] mux_457_nl;
  wire[0:0] mux_455_nl;
  wire[0:0] mux_456_nl;
  wire[0:0] nor_1604_nl;
  wire[0:0] mux_464_nl;
  wire[0:0] mux_462_nl;
  wire[0:0] mux_463_nl;
  wire[0:0] mux_466_nl;
  wire[0:0] and_3327_nl;
  wire[0:0] and_3328_nl;
  wire[0:0] mux_465_nl;
  wire[0:0] or_833_nl;
  wire[0:0] FpMul_6U_10U_1_FpMul_6U_10U_1_and_18_nl;
  wire[0:0] mux_469_nl;
  wire[0:0] mux_467_nl;
  wire[0:0] or_654_nl;
  wire[0:0] mux_468_nl;
  wire[0:0] mux_470_nl;
  wire[0:0] nor_1596_nl;
  wire[0:0] nor_1597_nl;
  wire[0:0] mux_471_nl;
  wire[0:0] and_3325_nl;
  wire[0:0] nor_1595_nl;
  wire[49:0] inp_lookup_1_FpAdd_8U_23U_1_if_2_acc_nl;
  wire[50:0] nl_inp_lookup_1_FpAdd_8U_23U_1_if_2_acc_nl;
  wire[49:0] inp_lookup_1_FpAdd_8U_23U_1_else_2_acc_nl;
  wire[51:0] nl_inp_lookup_1_FpAdd_8U_23U_1_else_2_acc_nl;
  wire[0:0] mux_474_nl;
  wire[0:0] nand_585_nl;
  wire[0:0] mux_475_nl;
  wire[7:0] FpMul_6U_10U_2_o_mant_asn_FpMul_6U_10U_2_o_mant_conc_80_cgspt_7_mux_nl;
  wire[0:0] and_1127_nl;
  wire[0:0] mux_1897_nl;
  wire[0:0] mux_2073_nl;
  wire[0:0] mux_2072_nl;
  wire[0:0] mux_2071_nl;
  wire[0:0] mux_2070_nl;
  wire[0:0] and_4166_nl;
  wire[0:0] mux_2078_nl;
  wire[0:0] mux_2077_nl;
  wire[0:0] mux_2076_nl;
  wire[0:0] mux_2075_nl;
  wire[0:0] mux_2074_nl;
  wire[0:0] and_4138_nl;
  wire[0:0] mux_481_nl;
  wire[0:0] and_3323_nl;
  wire[0:0] nor_1589_nl;
  wire[49:0] inp_lookup_2_FpAdd_8U_23U_1_if_2_acc_nl;
  wire[50:0] nl_inp_lookup_2_FpAdd_8U_23U_1_if_2_acc_nl;
  wire[49:0] inp_lookup_2_FpAdd_8U_23U_1_else_2_acc_nl;
  wire[51:0] nl_inp_lookup_2_FpAdd_8U_23U_1_else_2_acc_nl;
  wire[0:0] mux_484_nl;
  wire[0:0] nand_582_nl;
  wire[7:0] FpMul_6U_10U_2_o_mant_asn_FpMul_6U_10U_2_o_mant_conc_81_cgspt_7_mux_nl;
  wire[0:0] and_1135_nl;
  wire[0:0] mux_1898_nl;
  wire[0:0] mux_2082_nl;
  wire[0:0] mux_2081_nl;
  wire[0:0] mux_2080_nl;
  wire[0:0] mux_2079_nl;
  wire[0:0] and_4161_nl;
  wire[0:0] mux_2087_nl;
  wire[0:0] mux_2086_nl;
  wire[0:0] mux_2085_nl;
  wire[0:0] mux_2084_nl;
  wire[0:0] mux_2083_nl;
  wire[0:0] and_4133_nl;
  wire[0:0] mux_492_nl;
  wire[0:0] mux_490_nl;
  wire[0:0] mux_491_nl;
  wire[49:0] inp_lookup_3_FpAdd_8U_23U_1_if_2_acc_nl;
  wire[50:0] nl_inp_lookup_3_FpAdd_8U_23U_1_if_2_acc_nl;
  wire[49:0] inp_lookup_3_FpAdd_8U_23U_1_else_2_acc_nl;
  wire[51:0] nl_inp_lookup_3_FpAdd_8U_23U_1_else_2_acc_nl;
  wire[0:0] mux_499_nl;
  wire[0:0] nand_581_nl;
  wire[0:0] mux_2089_nl;
  wire[0:0] and_4130_nl;
  wire[0:0] mux_2088_nl;
  wire[0:0] and_4131_nl;
  wire[0:0] nor_1876_nl;
  wire[0:0] mux_2094_nl;
  wire[0:0] nor_1875_nl;
  wire[0:0] mux_2093_nl;
  wire[0:0] mux_2092_nl;
  wire[0:0] or_5992_nl;
  wire[0:0] mux_2091_nl;
  wire[0:0] or_5993_nl;
  wire[0:0] or_5994_nl;
  wire[7:0] FpMul_6U_10U_2_o_mant_asn_FpMul_6U_10U_2_o_mant_conc_82_cgspt_7_mux_nl;
  wire[0:0] and_1143_nl;
  wire[0:0] mux_2098_nl;
  wire[0:0] mux_2097_nl;
  wire[0:0] mux_2096_nl;
  wire[0:0] mux_2095_nl;
  wire[0:0] and_4156_nl;
  wire[0:0] mux_2103_nl;
  wire[0:0] mux_2102_nl;
  wire[0:0] mux_2101_nl;
  wire[0:0] mux_2100_nl;
  wire[0:0] mux_2099_nl;
  wire[0:0] and_4123_nl;
  wire[0:0] mux_510_nl;
  wire[0:0] and_3319_nl;
  wire[0:0] nor_1578_nl;
  wire[49:0] inp_lookup_4_FpAdd_8U_23U_1_if_2_acc_nl;
  wire[50:0] nl_inp_lookup_4_FpAdd_8U_23U_1_if_2_acc_nl;
  wire[49:0] inp_lookup_4_FpAdd_8U_23U_1_else_2_acc_nl;
  wire[51:0] nl_inp_lookup_4_FpAdd_8U_23U_1_else_2_acc_nl;
  wire[0:0] mux_513_nl;
  wire[7:0] mux_2004_nl;
  wire[0:0] and_1151_nl;
  wire[0:0] mux_1900_nl;
  wire[0:0] mux_515_nl;
  wire[0:0] nor_1572_nl;
  wire[0:0] mux_514_nl;
  wire[0:0] nor_1574_nl;
  wire[0:0] nor_1575_nl;
  wire[0:0] and_1166_nl;
  wire[0:0] and_3443_nl;
  wire[0:0] or_6170_nl;
  wire[0:0] and_1172_nl;
  wire[0:0] mux_517_nl;
  wire[0:0] mux_518_nl;
  wire[0:0] mux_521_nl;
  wire[0:0] nor_1568_nl;
  wire[0:0] mux_520_nl;
  wire[0:0] nor_1569_nl;
  wire[0:0] nor_1570_nl;
  wire[0:0] mux_526_nl;
  wire[0:0] mux_525_nl;
  wire[0:0] mux_523_nl;
  wire[0:0] mux_524_nl;
  wire[0:0] mux_529_nl;
  wire[0:0] mux_527_nl;
  wire[0:0] nor_1562_nl;
  wire[0:0] nor_1564_nl;
  wire[0:0] nor_1566_nl;
  wire[0:0] mux_528_nl;
  wire[0:0] nor_1567_nl;
  wire[0:0] and_1177_nl;
  wire[0:0] and_3444_nl;
  wire[0:0] or_6171_nl;
  wire[0:0] and_1183_nl;
  wire[0:0] mux_531_nl;
  wire[0:0] mux_534_nl;
  wire[0:0] nor_1559_nl;
  wire[0:0] mux_533_nl;
  wire[0:0] nor_1560_nl;
  wire[0:0] nor_1561_nl;
  wire[0:0] mux_539_nl;
  wire[0:0] mux_538_nl;
  wire[0:0] mux_536_nl;
  wire[0:0] mux_537_nl;
  wire[0:0] and_1188_nl;
  wire[0:0] nor_1910_nl;
  wire[0:0] and_4169_nl;
  wire[0:0] mux_541_nl;
  wire[0:0] mux_544_nl;
  wire[0:0] nor_1557_nl;
  wire[0:0] nor_1558_nl;
  wire[0:0] mux_547_nl;
  wire[0:0] mux_546_nl;
  wire[0:0] mux_550_nl;
  wire[0:0] mux_548_nl;
  wire[0:0] nor_1552_nl;
  wire[0:0] nor_1553_nl;
  wire[0:0] mux_549_nl;
  wire[0:0] nor_1554_nl;
  wire[0:0] nor_1555_nl;
  wire[0:0] and_1195_nl;
  wire[0:0] and_3446_nl;
  wire[0:0] or_6172_nl;
  wire[0:0] and_1201_nl;
  wire[0:0] mux_552_nl;
  wire[0:0] mux_555_nl;
  wire[0:0] nor_1549_nl;
  wire[0:0] mux_554_nl;
  wire[0:0] nor_1550_nl;
  wire[0:0] nor_1551_nl;
  wire[0:0] mux_558_nl;
  wire[0:0] mux_557_nl;
  wire[0:0] or_1054_nl;
  wire[0:0] or_1057_nl;
  wire[0:0] and_4221_nl;
  wire[0:0] mux_562_nl;
  wire[0:0] and_3314_nl;
  wire[0:0] mux_561_nl;
  wire[0:0] mux_560_nl;
  wire[0:0] nor_1545_nl;
  wire[0:0] and_3315_nl;
  wire[0:0] mux_563_nl;
  wire[0:0] nor_1543_nl;
  wire[0:0] nor_1544_nl;
  wire[0:0] mux_565_nl;
  wire[0:0] nor_1540_nl;
  wire[0:0] mux_567_nl;
  wire[0:0] mux_569_nl;
  wire[0:0] nor_1535_nl;
  wire[0:0] mux_568_nl;
  wire[0:0] nor_1536_nl;
  wire[0:0] nor_1537_nl;
  wire[0:0] mux_570_nl;
  wire[0:0] or_1102_nl;
  wire[0:0] FpNormalize_6U_23U_1_if_or_nl;
  wire[0:0] mux_572_nl;
  wire[0:0] mux_571_nl;
  wire[0:0] FpAdd_6U_10U_1_mux_2_nl;
  wire[0:0] or_1106_nl;
  wire[0:0] and_4220_nl;
  wire[0:0] mux_575_nl;
  wire[0:0] nor_1530_nl;
  wire[0:0] mux_574_nl;
  wire[0:0] and_3387_nl;
  wire[0:0] and_3309_nl;
  wire[0:0] mux_576_nl;
  wire[0:0] nor_1528_nl;
  wire[0:0] nor_1529_nl;
  wire[0:0] mux_578_nl;
  wire[0:0] nor_1524_nl;
  wire[0:0] nor_1525_nl;
  wire[0:0] mux_581_nl;
  wire[0:0] nor_1518_nl;
  wire[0:0] mux_580_nl;
  wire[0:0] nor_1519_nl;
  wire[0:0] nor_1520_nl;
  wire[0:0] mux_582_nl;
  wire[0:0] or_1147_nl;
  wire[0:0] FpNormalize_6U_23U_1_if_or_1_nl;
  wire[0:0] mux_585_nl;
  wire[0:0] mux_583_nl;
  wire[0:0] FpAdd_6U_10U_1_mux_18_nl;
  wire[0:0] mux_584_nl;
  wire[0:0] mux_590_nl;
  wire[0:0] nor_1514_nl;
  wire[0:0] mux_589_nl;
  wire[0:0] and_3307_nl;
  wire[0:0] mux_588_nl;
  wire[0:0] nor_1516_nl;
  wire[0:0] mux_592_nl;
  wire[0:0] nor_1512_nl;
  wire[0:0] mux_595_nl;
  wire[0:0] or_1179_nl;
  wire[0:0] mux_594_nl;
  wire[0:0] or_1182_nl;
  wire[0:0] mux_596_nl;
  wire[0:0] or_1189_nl;
  wire[0:0] FpNormalize_6U_23U_1_if_or_2_nl;
  wire[0:0] mux_597_nl;
  wire[0:0] nor_1507_nl;
  wire[0:0] FpAdd_6U_10U_1_mux_34_nl;
  wire[0:0] nor_1509_nl;
  wire[0:0] and_4219_nl;
  wire[0:0] mux_601_nl;
  wire[0:0] nor_1504_nl;
  wire[0:0] mux_600_nl;
  wire[0:0] and_3386_nl;
  wire[0:0] and_3300_nl;
  wire[0:0] mux_602_nl;
  wire[0:0] nor_1502_nl;
  wire[0:0] nor_1503_nl;
  wire[0:0] mux_604_nl;
  wire[0:0] nor_1500_nl;
  wire[0:0] nor_1501_nl;
  wire[0:0] mux_609_nl;
  wire[0:0] or_1232_nl;
  wire[0:0] mux_608_nl;
  wire[0:0] mux_607_nl;
  wire[0:0] mux_606_nl;
  wire[0:0] or_1236_nl;
  wire[0:0] nor_158_nl;
  wire[0:0] mux_610_nl;
  wire[0:0] FpNormalize_6U_23U_1_if_or_3_nl;
  wire[0:0] mux_611_nl;
  wire[0:0] nor_1496_nl;
  wire[0:0] FpAdd_6U_10U_1_mux_50_nl;
  wire[0:0] nor_1498_nl;
  wire[0:0] nand_62_nl;
  wire[0:0] mux_614_nl;
  wire[0:0] mux_619_nl;
  wire[0:0] nor_1491_nl;
  wire[0:0] mux_616_nl;
  wire[0:0] and_3293_nl;
  wire[0:0] mux_618_nl;
  wire[0:0] mux_617_nl;
  wire[0:0] nor_1492_nl;
  wire[0:0] inp_lookup_1_IsInf_6U_23U_1_IsInf_6U_23U_1_and_nl;
  wire[0:0] mux_620_nl;
  wire[0:0] nor_1489_nl;
  wire[0:0] mux_621_nl;
  wire[0:0] mux_622_nl;
  wire[0:0] inp_lookup_1_FpMul_6U_10U_xor_1_nl;
  wire[0:0] mux_625_nl;
  wire[0:0] nor_1486_nl;
  wire[0:0] mux_624_nl;
  wire[0:0] or_1284_nl;
  wire[0:0] mux_629_nl;
  wire[0:0] nor_1482_nl;
  wire[0:0] mux_626_nl;
  wire[0:0] and_3291_nl;
  wire[0:0] mux_628_nl;
  wire[0:0] mux_627_nl;
  wire[0:0] nor_1483_nl;
  wire[0:0] inp_lookup_2_IsInf_6U_23U_1_IsInf_6U_23U_1_and_nl;
  wire[0:0] mux_630_nl;
  wire[0:0] nor_1480_nl;
  wire[0:0] nor_1481_nl;
  wire[0:0] mux_631_nl;
  wire[0:0] inp_lookup_2_FpMul_6U_10U_xor_1_nl;
  wire[0:0] nand_561_nl;
  wire[0:0] mux_634_nl;
  wire[0:0] inp_lookup_3_IsInf_6U_23U_1_IsInf_6U_23U_1_and_nl;
  wire[0:0] mux_640_nl;
  wire[0:0] nor_1474_nl;
  wire[0:0] nor_1475_nl;
  wire[0:0] mux_641_nl;
  wire[0:0] inp_lookup_3_FpMul_6U_10U_xor_1_nl;
  wire[0:0] nand_560_nl;
  wire[0:0] mux_644_nl;
  wire[0:0] mux_649_nl;
  wire[0:0] nor_1470_nl;
  wire[0:0] mux_646_nl;
  wire[0:0] and_3287_nl;
  wire[0:0] mux_648_nl;
  wire[0:0] mux_647_nl;
  wire[0:0] nor_1471_nl;
  wire[0:0] inp_lookup_4_IsInf_6U_23U_1_IsInf_6U_23U_1_and_nl;
  wire[0:0] mux_650_nl;
  wire[0:0] nor_1468_nl;
  wire[0:0] mux_651_nl;
  wire[0:0] inp_lookup_4_FpMul_6U_10U_xor_1_nl;
  wire[5:0] FpMul_6U_10U_else_2_else_acc_nl;
  wire[6:0] nl_FpMul_6U_10U_else_2_else_acc_nl;
  wire[0:0] mux_654_nl;
  wire[0:0] nor_1464_nl;
  wire[0:0] nor_1465_nl;
  wire[0:0] mux_656_nl;
  wire[0:0] nor_1912_nl;
  wire[0:0] nor_1463_nl;
  wire[0:0] mux_660_nl;
  wire[5:0] FpMul_6U_10U_else_2_else_acc_2_nl;
  wire[6:0] nl_FpMul_6U_10U_else_2_else_acc_2_nl;
  wire[0:0] mux_662_nl;
  wire[0:0] nor_1454_nl;
  wire[0:0] nor_1455_nl;
  wire[0:0] mux_664_nl;
  wire[0:0] nor_1452_nl;
  wire[0:0] nor_1453_nl;
  wire[0:0] mux_667_nl;
  wire[5:0] FpMul_6U_10U_else_2_else_acc_3_nl;
  wire[6:0] nl_FpMul_6U_10U_else_2_else_acc_3_nl;
  wire[0:0] mux_669_nl;
  wire[0:0] nor_1446_nl;
  wire[0:0] nor_1447_nl;
  wire[0:0] mux_671_nl;
  wire[0:0] and_3284_nl;
  wire[0:0] nor_1445_nl;
  wire[0:0] mux_674_nl;
  wire[5:0] FpMul_6U_10U_else_2_else_acc_4_nl;
  wire[6:0] nl_FpMul_6U_10U_else_2_else_acc_4_nl;
  wire[0:0] mux_676_nl;
  wire[0:0] nor_1441_nl;
  wire[0:0] nor_1442_nl;
  wire[0:0] mux_678_nl;
  wire[0:0] and_3282_nl;
  wire[0:0] nor_1440_nl;
  wire[0:0] mux_681_nl;
  wire[0:0] mux_682_nl;
  wire[0:0] mux_685_nl;
  wire[0:0] and_4207_nl;
  wire[0:0] mux_690_nl;
  wire[0:0] nor_1435_nl;
  wire[0:0] mux_698_nl;
  wire[0:0] nand_776_nl;
  wire[0:0] mux_699_nl;
  wire[0:0] mux_700_nl;
  wire[0:0] mux_703_nl;
  wire[0:0] and_4206_nl;
  wire[0:0] mux_708_nl;
  wire[0:0] nor_1430_nl;
  wire[0:0] mux_716_nl;
  wire[0:0] nand_775_nl;
  wire[0:0] mux_717_nl;
  wire[0:0] mux_718_nl;
  wire[0:0] mux_721_nl;
  wire[0:0] and_4205_nl;
  wire[0:0] mux_726_nl;
  wire[0:0] nor_1425_nl;
  wire[0:0] mux_734_nl;
  wire[0:0] mux_736_nl;
  wire[0:0] mux_739_nl;
  wire[0:0] and_4204_nl;
  wire[0:0] mux_744_nl;
  wire[0:0] nor_1420_nl;
  wire[0:0] mux_752_nl;
  wire[0:0] mux_754_nl;
  wire[0:0] mux_755_nl;
  wire[0:0] mux_756_nl;
  wire[0:0] mux_760_nl;
  wire[0:0] mux_761_nl;
  wire[0:0] mux_765_nl;
  wire[0:0] mux_766_nl;
  wire[0:0] mux_770_nl;
  wire[0:0] mux_771_nl;
  wire[0:0] mux_775_nl;
  wire[0:0] mux_780_nl;
  wire[0:0] mux_777_nl;
  wire[0:0] nand_491_nl;
  wire[0:0] mux_779_nl;
  wire[0:0] or_5699_nl;
  wire[0:0] mux_778_nl;
  wire[0:0] mux_781_nl;
  wire[0:0] nor_1418_nl;
  wire[0:0] and_3276_nl;
  wire[0:0] mux_784_nl;
  wire[0:0] or_1676_nl;
  wire[0:0] mux_783_nl;
  wire[0:0] or_1679_nl;
  wire[0:0] mux_785_nl;
  wire[0:0] nor_1415_nl;
  wire[0:0] nor_1416_nl;
  wire[0:0] mux_788_nl;
  wire[0:0] mux_787_nl;
  wire[0:0] nand_87_nl;
  wire[0:0] mux_790_nl;
  wire[0:0] mux_789_nl;
  wire[0:0] mux_791_nl;
  wire[0:0] and_3275_nl;
  wire[0:0] mux_797_nl;
  wire[0:0] or_1697_nl;
  wire[0:0] mux_796_nl;
  wire[0:0] mux_794_nl;
  wire[0:0] mux_792_nl;
  wire[0:0] mux_795_nl;
  wire[0:0] or_1705_nl;
  wire[0:0] mux_798_nl;
  wire[0:0] or_1708_nl;
  wire[0:0] mux_800_nl;
  wire[0:0] or_1712_nl;
  wire[0:0] mux_801_nl;
  wire[0:0] nor_1410_nl;
  wire[0:0] nor_1411_nl;
  wire[0:0] mux_802_nl;
  wire[0:0] nor_1408_nl;
  wire[0:0] mux_804_nl;
  wire[0:0] mux_803_nl;
  wire[0:0] or_1732_nl;
  wire[0:0] mux_805_nl;
  wire[0:0] and_3274_nl;
  wire[0:0] mux_814_nl;
  wire[0:0] mux_807_nl;
  wire[0:0] mux_806_nl;
  wire[0:0] nand_88_nl;
  wire[0:0] or_1740_nl;
  wire[0:0] mux_813_nl;
  wire[0:0] mux_812_nl;
  wire[0:0] mux_808_nl;
  wire[0:0] mux_810_nl;
  wire[0:0] or_1745_nl;
  wire[0:0] mux_815_nl;
  wire[0:0] nor_1404_nl;
  wire[0:0] nor_1405_nl;
  wire[0:0] mux_818_nl;
  wire[0:0] nor_1400_nl;
  wire[0:0] mux_817_nl;
  wire[0:0] nor_1402_nl;
  wire[0:0] nor_1403_nl;
  wire[0:0] mux_819_nl;
  wire[0:0] or_1763_nl;
  wire[0:0] mux_820_nl;
  wire[0:0] nor_1398_nl;
  wire[0:0] mux_822_nl;
  wire[0:0] mux_821_nl;
  wire[0:0] or_1778_nl;
  wire[0:0] mux_823_nl;
  wire[0:0] and_3273_nl;
  wire[0:0] mux_827_nl;
  wire[0:0] or_1782_nl;
  wire[0:0] mux_826_nl;
  wire[0:0] mux_824_nl;
  wire[0:0] nand_667_nl;
  wire[0:0] mux_825_nl;
  wire[0:0] mux_828_nl;
  wire[0:0] nor_1394_nl;
  wire[0:0] and_3384_nl;
  wire[0:0] mux_830_nl;
  wire[0:0] or_1797_nl;
  wire[0:0] mux_831_nl;
  wire[0:0] nor_1392_nl;
  wire[0:0] nor_1393_nl;
  wire[0:0] mux_833_nl;
  wire[0:0] nand_665_nl;
  wire[0:0] mux_834_nl;
  wire[0:0] nand_664_nl;
  wire[0:0] mux_835_nl;
  wire[0:0] and_3272_nl;
  wire[0:0] mux_836_nl;
  wire[0:0] mux_837_nl;
  wire[0:0] or_1821_nl;
  wire[0:0] mux_839_nl;
  wire[0:0] mux_838_nl;
  wire[0:0] nor_1387_nl;
  wire[0:0] mux_841_nl;
  wire[0:0] or_1826_nl;
  wire[0:0] mux_840_nl;
  wire[0:0] or_1830_nl;
  wire[0:0] mux_844_nl;
  wire[0:0] mux_843_nl;
  wire[0:0] nor_1386_nl;
  wire[0:0] mux_846_nl;
  wire[0:0] or_1837_nl;
  wire[0:0] mux_845_nl;
  wire[0:0] or_1840_nl;
  wire[0:0] mux_842_nl;
  wire[0:0] or_1832_nl;
  wire[0:0] mux_847_nl;
  wire[0:0] or_1843_nl;
  wire[0:0] mux_848_nl;
  wire[0:0] and_3266_nl;
  wire[0:0] mux_849_nl;
  wire[0:0] or_1849_nl;
  wire[0:0] mux_852_nl;
  wire[0:0] mux_851_nl;
  wire[0:0] nor_1385_nl;
  wire[0:0] mux_853_nl;
  wire[0:0] or_1860_nl;
  wire[0:0] mux_850_nl;
  wire[0:0] or_1852_nl;
  wire[0:0] FpMul_6U_10U_2_o_mant_or_nl;
  wire[0:0] mux_1919_nl;
  wire[0:0] mux_1872_nl;
  wire[0:0] nor_732_nl;
  wire[0:0] or_4349_nl;
  wire[0:0] or_4671_nl;
  wire[0:0] mux_865_nl;
  wire[0:0] mux_861_nl;
  wire[0:0] mux_858_nl;
  wire[0:0] mux_856_nl;
  wire[0:0] nand_89_nl;
  wire[0:0] mux_855_nl;
  wire[0:0] nor_1375_nl;
  wire[0:0] nor_1377_nl;
  wire[0:0] mux_864_nl;
  wire[0:0] mux_862_nl;
  wire[0:0] nor_1378_nl;
  wire[0:0] nor_1379_nl;
  wire[0:0] mux_863_nl;
  wire[0:0] mux_871_nl;
  wire[0:0] mux_867_nl;
  wire[0:0] mux_866_nl;
  wire[0:0] or_1889_nl;
  wire[0:0] mux_870_nl;
  wire[0:0] mux_868_nl;
  wire[0:0] nor_1372_nl;
  wire[0:0] mux_869_nl;
  wire[0:0] nor_1373_nl;
  wire[0:0] mux_888_nl;
  wire[0:0] mux_884_nl;
  wire[0:0] mux_883_nl;
  wire[0:0] or_1927_nl;
  wire[0:0] mux_887_nl;
  wire[0:0] mux_885_nl;
  wire[0:0] nor_1359_nl;
  wire[0:0] mux_886_nl;
  wire[0:0] nor_1360_nl;
  wire[0:0] mux_899_nl;
  wire[0:0] mux_895_nl;
  wire[0:0] mux_892_nl;
  wire[0:0] mux_890_nl;
  wire[0:0] nand_97_nl;
  wire[0:0] mux_889_nl;
  wire[0:0] nor_1349_nl;
  wire[0:0] nor_1351_nl;
  wire[0:0] mux_898_nl;
  wire[0:0] mux_896_nl;
  wire[0:0] nor_1352_nl;
  wire[0:0] nor_1353_nl;
  wire[0:0] mux_897_nl;
  wire[0:0] mux_905_nl;
  wire[0:0] mux_901_nl;
  wire[0:0] mux_900_nl;
  wire[0:0] or_1965_nl;
  wire[0:0] nor_279_nl;
  wire[0:0] mux_904_nl;
  wire[0:0] mux_902_nl;
  wire[0:0] nor_1346_nl;
  wire[0:0] mux_903_nl;
  wire[0:0] nor_1347_nl;
  wire[7:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_asn_FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_conc_10_cgspt_7_mux_nl;
  wire[0:0] mux_918_nl;
  wire[0:0] inp_lookup_2_IsZero_6U_10U_1_IsZero_6U_10U_1_nor_nl;
  wire[0:0] mux_919_nl;
  wire[0:0] mux_920_nl;
  wire[0:0] inp_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_nl;
  wire[0:0] IsZero_6U_10U_5_IsZero_6U_10U_5_and_1_nl;
  wire[0:0] inp_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_nl;
  wire[0:0] IsZero_6U_10U_5_IsZero_6U_10U_5_and_3_nl;
  wire[0:0] mux_921_nl;
  wire[0:0] mux_922_nl;
  wire[0:0] mux_923_nl;
  wire[0:0] mux_924_nl;
  wire[0:0] and_1693_nl;
  wire[0:0] and_1695_nl;
  wire[0:0] mux_1924_nl;
  wire[0:0] mux_2106_nl;
  wire[0:0] mux_2105_nl;
  wire[0:0] mux_2109_nl;
  wire[0:0] and_4209_nl;
  wire[0:0] mux_1925_nl;
  wire[0:0] mux_2113_nl;
  wire[0:0] mux_2112_nl;
  wire[0:0] and_1711_nl;
  wire[0:0] and_1714_nl;
  wire[0:0] mux_1926_nl;
  wire[0:0] mux_2116_nl;
  wire[0:0] mux_2115_nl;
  wire[0:0] mux_939_nl;
  wire[0:0] and_227_nl;
  wire[0:0] mux_118_nl;
  wire[0:0] mux_117_nl;
  wire[0:0] or_171_nl;
  wire[0:0] or_174_nl;
  wire[0:0] mux_940_nl;
  wire[0:0] nor_1310_nl;
  wire[0:0] and_3251_nl;
  wire[0:0] mux_123_nl;
  wire[0:0] mux_121_nl;
  wire[0:0] mux_120_nl;
  wire[0:0] nor_1695_nl;
  wire[0:0] and_3392_nl;
  wire[0:0] mux_122_nl;
  wire[0:0] nor_1698_nl;
  wire[0:0] or_192_nl;
  wire[0:0] mux_941_nl;
  wire[0:0] and_231_nl;
  wire[0:0] mux_140_nl;
  wire[0:0] or_239_nl;
  wire[0:0] mux_942_nl;
  wire[0:0] nor_1309_nl;
  wire[0:0] and_3250_nl;
  wire[0:0] mux_146_nl;
  wire[0:0] mux_144_nl;
  wire[0:0] mux_143_nl;
  wire[0:0] nor_1677_nl;
  wire[0:0] and_3390_nl;
  wire[0:0] mux_145_nl;
  wire[0:0] nor_1680_nl;
  wire[0:0] or_258_nl;
  wire[0:0] mux_943_nl;
  wire[0:0] and_235_nl;
  wire[0:0] mux_163_nl;
  wire[0:0] mux_162_nl;
  wire[0:0] or_311_nl;
  wire[0:0] or_314_nl;
  wire[0:0] mux_946_nl;
  wire[0:0] nor_1305_nl;
  wire[0:0] mux_944_nl;
  wire[0:0] nand_458_nl;
  wire[0:0] mux_945_nl;
  wire[0:0] nor_1307_nl;
  wire[0:0] or_2090_nl;
  wire[0:0] mux_947_nl;
  wire[0:0] and_237_nl;
  wire[0:0] mux_180_nl;
  wire[0:0] or_374_nl;
  wire[0:0] mux_948_nl;
  wire[0:0] nor_1304_nl;
  wire[0:0] and_3248_nl;
  wire[0:0] mux_951_nl;
  wire[0:0] mux_949_nl;
  wire[0:0] nor_1300_nl;
  wire[0:0] nor_1301_nl;
  wire[0:0] mux_950_nl;
  wire[0:0] nor_1302_nl;
  wire[0:0] nor_1303_nl;
  wire[0:0] mux_954_nl;
  wire[0:0] mux_952_nl;
  wire[0:0] nor_1296_nl;
  wire[0:0] nor_1297_nl;
  wire[0:0] mux_953_nl;
  wire[0:0] nor_1298_nl;
  wire[0:0] nor_1299_nl;
  wire[0:0] mux_957_nl;
  wire[0:0] mux_955_nl;
  wire[0:0] nor_1292_nl;
  wire[0:0] nor_1293_nl;
  wire[0:0] mux_956_nl;
  wire[0:0] nor_1294_nl;
  wire[0:0] nor_1295_nl;
  wire[0:0] mux_960_nl;
  wire[0:0] mux_958_nl;
  wire[0:0] nor_1288_nl;
  wire[0:0] nor_1289_nl;
  wire[0:0] mux_959_nl;
  wire[0:0] nor_1290_nl;
  wire[0:0] nor_1291_nl;
  wire[0:0] mux_962_nl;
  wire[0:0] mux_961_nl;
  wire[0:0] nor_1284_nl;
  wire[0:0] nor_1285_nl;
  wire[0:0] mux_964_nl;
  wire[0:0] mux_963_nl;
  wire[0:0] nor_1279_nl;
  wire[0:0] nor_1280_nl;
  wire[0:0] mux_966_nl;
  wire[0:0] mux_965_nl;
  wire[0:0] nor_1275_nl;
  wire[0:0] nor_1276_nl;
  wire[0:0] mux_210_nl;
  wire[0:0] mux_214_nl;
  wire[0:0] or_460_nl;
  wire[0:0] or_458_nl;
  wire[0:0] FpMul_6U_10U_2_else_2_else_and_nl;
  wire[0:0] mux_970_nl;
  wire[0:0] mux_969_nl;
  wire[0:0] mux_968_nl;
  wire[0:0] mux_967_nl;
  wire[0:0] or_2179_nl;
  wire[0:0] or_2174_nl;
  wire[0:0] or_2171_nl;
  wire[0:0] or_2185_nl;
  wire[0:0] mux_971_nl;
  wire[0:0] nor_1267_nl;
  wire[0:0] nor_1268_nl;
  wire[0:0] mux_972_nl;
  wire[0:0] nor_1265_nl;
  wire[0:0] nor_1266_nl;
  wire[0:0] mux_975_nl;
  wire[0:0] and_3230_nl;
  wire[0:0] mux_973_nl;
  wire[0:0] or_2197_nl;
  wire[0:0] and_3231_nl;
  wire[0:0] mux_974_nl;
  wire[0:0] or_2198_nl;
  wire[0:0] FpMul_6U_10U_2_FpMul_6U_10U_2_and_nl;
  wire[0:0] mux_248_nl;
  wire[0:0] or_520_nl;
  wire[0:0] mux_252_nl;
  wire[0:0] or_522_nl;
  wire[0:0] mux_976_nl;
  wire[0:0] nor_1261_nl;
  wire[0:0] nor_1263_nl;
  wire[0:0] FpMul_6U_10U_2_else_2_else_and_1_nl;
  wire[0:0] mux_980_nl;
  wire[0:0] mux_979_nl;
  wire[0:0] mux_978_nl;
  wire[0:0] mux_977_nl;
  wire[0:0] or_2216_nl;
  wire[0:0] or_2211_nl;
  wire[0:0] or_2223_nl;
  wire[0:0] mux_981_nl;
  wire[0:0] nor_1254_nl;
  wire[0:0] nor_1255_nl;
  wire[0:0] mux_982_nl;
  wire[0:0] nor_1252_nl;
  wire[0:0] nor_1253_nl;
  wire[0:0] mux_985_nl;
  wire[0:0] and_3228_nl;
  wire[0:0] mux_983_nl;
  wire[0:0] or_2232_nl;
  wire[0:0] and_3229_nl;
  wire[0:0] mux_984_nl;
  wire[0:0] or_2233_nl;
  wire[0:0] FpMul_6U_10U_2_FpMul_6U_10U_2_and_16_nl;
  wire[0:0] mux_286_nl;
  wire[0:0] mux_297_nl;
  wire[0:0] or_596_nl;
  wire[0:0] or_594_nl;
  wire[0:0] mux_986_nl;
  wire[0:0] nor_1248_nl;
  wire[0:0] nor_1250_nl;
  wire[0:0] FpMul_6U_10U_2_else_2_else_and_2_nl;
  wire[0:0] mux_990_nl;
  wire[0:0] mux_989_nl;
  wire[0:0] mux_988_nl;
  wire[0:0] mux_987_nl;
  wire[0:0] or_2254_nl;
  wire[0:0] or_2246_nl;
  wire[0:0] or_2260_nl;
  wire[0:0] mux_991_nl;
  wire[0:0] nor_1241_nl;
  wire[0:0] nor_1242_nl;
  wire[0:0] mux_992_nl;
  wire[0:0] nor_1239_nl;
  wire[0:0] nor_1240_nl;
  wire[0:0] mux_995_nl;
  wire[0:0] mux_993_nl;
  wire[0:0] or_2269_nl;
  wire[0:0] nand_116_nl;
  wire[0:0] mux_994_nl;
  wire[0:0] or_2270_nl;
  wire[0:0] FpMul_6U_10U_2_FpMul_6U_10U_2_and_17_nl;
  wire[0:0] mux_336_nl;
  wire[0:0] or_640_nl;
  wire[0:0] or_642_nl;
  wire[0:0] FpMul_6U_10U_2_else_2_else_and_3_nl;
  wire[0:0] mux_1001_nl;
  wire[0:0] mux_998_nl;
  wire[0:0] mux_997_nl;
  wire[0:0] mux_996_nl;
  wire[0:0] or_2277_nl;
  wire[0:0] or_2274_nl;
  wire[0:0] or_2272_nl;
  wire[0:0] mux_1000_nl;
  wire[0:0] mux_999_nl;
  wire[0:0] or_2287_nl;
  wire[0:0] or_2278_nl;
  wire[0:0] mux_1002_nl;
  wire[0:0] nor_1233_nl;
  wire[0:0] nor_1234_nl;
  wire[0:0] mux_1003_nl;
  wire[0:0] nor_1231_nl;
  wire[0:0] nor_1232_nl;
  wire[0:0] mux_1005_nl;
  wire[0:0] and_3226_nl;
  wire[0:0] mux_1004_nl;
  wire[0:0] or_2296_nl;
  wire[0:0] and_3227_nl;
  wire[0:0] FpMul_6U_10U_2_FpMul_6U_10U_2_and_18_nl;
  wire[0:0] mux_1006_nl;
  wire[0:0] nor_1226_nl;
  wire[0:0] nor_1227_nl;
  wire[0:0] mux_1927_nl;
  wire[0:0] FpMul_6U_10U_1_else_2_else_and_nl;
  wire[0:0] mux_1011_nl;
  wire[0:0] mux_1008_nl;
  wire[0:0] and_3222_nl;
  wire[0:0] mux_1007_nl;
  wire[0:0] nor_1218_nl;
  wire[0:0] or_2308_nl;
  wire[0:0] or_2306_nl;
  wire[0:0] mux_1010_nl;
  wire[0:0] and_3397_nl;
  wire[0:0] mux_1009_nl;
  wire[0:0] nor_1222_nl;
  wire[0:0] or_2313_nl;
  wire[0:0] mux_1014_nl;
  wire[0:0] nor_1215_nl;
  wire[0:0] and_3220_nl;
  wire[0:0] mux_1013_nl;
  wire[0:0] and_3221_nl;
  wire[0:0] nor_1216_nl;
  wire[0:0] and_4218_nl;
  wire[0:0] mux_1017_nl;
  wire[0:0] nor_1213_nl;
  wire[0:0] nor_1214_nl;
  wire[0:0] mux_1016_nl;
  wire[0:0] mux_1022_nl;
  wire[0:0] nor_1209_nl;
  wire[0:0] mux_1019_nl;
  wire[0:0] nor_1211_nl;
  wire[0:0] mux_1021_nl;
  wire[0:0] mux_1020_nl;
  wire[0:0] nor_1212_nl;
  wire[0:0] mux_1928_nl;
  wire[0:0] FpMul_6U_10U_1_else_2_else_and_1_nl;
  wire[0:0] mux_1027_nl;
  wire[0:0] mux_1024_nl;
  wire[0:0] and_3218_nl;
  wire[0:0] mux_1023_nl;
  wire[0:0] nor_1201_nl;
  wire[0:0] or_2345_nl;
  wire[0:0] or_2343_nl;
  wire[0:0] mux_1026_nl;
  wire[0:0] and_3396_nl;
  wire[0:0] mux_1025_nl;
  wire[0:0] nor_1205_nl;
  wire[0:0] or_2350_nl;
  wire[0:0] mux_1030_nl;
  wire[0:0] and_3216_nl;
  wire[0:0] and_3217_nl;
  wire[0:0] mux_1029_nl;
  wire[0:0] nor_1198_nl;
  wire[0:0] nor_1199_nl;
  wire[0:0] and_4217_nl;
  wire[0:0] mux_1033_nl;
  wire[0:0] nor_1196_nl;
  wire[0:0] nor_1197_nl;
  wire[0:0] mux_1032_nl;
  wire[0:0] mux_1038_nl;
  wire[0:0] nor_1192_nl;
  wire[0:0] mux_1035_nl;
  wire[0:0] nor_1194_nl;
  wire[0:0] mux_1037_nl;
  wire[0:0] mux_1036_nl;
  wire[0:0] nor_1195_nl;
  wire[0:0] mux_1929_nl;
  wire[0:0] FpMul_6U_10U_1_else_2_else_and_2_nl;
  wire[0:0] mux_1043_nl;
  wire[0:0] mux_1040_nl;
  wire[0:0] and_3214_nl;
  wire[0:0] mux_1039_nl;
  wire[0:0] nor_1184_nl;
  wire[0:0] or_2382_nl;
  wire[0:0] or_2380_nl;
  wire[0:0] mux_1042_nl;
  wire[0:0] and_3395_nl;
  wire[0:0] mux_1041_nl;
  wire[0:0] nor_1188_nl;
  wire[0:0] or_2387_nl;
  wire[0:0] mux_1046_nl;
  wire[0:0] and_3212_nl;
  wire[0:0] and_3213_nl;
  wire[0:0] and_4216_nl;
  wire[0:0] mux_1049_nl;
  wire[0:0] nor_1181_nl;
  wire[0:0] mux_1047_nl;
  wire[0:0] nor_1182_nl;
  wire[0:0] mux_1048_nl;
  wire[0:0] mux_1052_nl;
  wire[0:0] and_3210_nl;
  wire[0:0] mux_1050_nl;
  wire[0:0] or_2410_nl;
  wire[0:0] and_3211_nl;
  wire[0:0] mux_1051_nl;
  wire[0:0] or_2411_nl;
  wire[0:0] mux_1930_nl;
  wire[0:0] FpMul_6U_10U_1_else_2_else_and_3_nl;
  wire[0:0] mux_1056_nl;
  wire[0:0] mux_1054_nl;
  wire[0:0] or_2418_nl;
  wire[0:0] mux_1053_nl;
  wire[0:0] nand_433_nl;
  wire[0:0] or_2415_nl;
  wire[0:0] or_2427_nl;
  wire[0:0] mux_1055_nl;
  wire[0:0] nor_1178_nl;
  wire[0:0] nor_1179_nl;
  wire[0:0] mux_1060_nl;
  wire[0:0] mux_1058_nl;
  wire[0:0] nand_432_nl;
  wire[0:0] mux_1059_nl;
  wire[0:0] or_2433_nl;
  wire[0:0] and_4117_nl;
  wire[0:0] mux_1063_nl;
  wire[0:0] nor_1173_nl;
  wire[0:0] nor_1174_nl;
  wire[0:0] mux_1062_nl;
  wire[0:0] mux_1065_nl;
  wire[0:0] nor_1171_nl;
  wire[0:0] mux_1064_nl;
  wire[0:0] nor_1172_nl;
  wire[0:0] mux_1068_nl;
  wire[0:0] nor_1169_nl;
  wire[0:0] nor_1170_nl;
  wire[0:0] mux_1070_nl;
  wire[0:0] nor_1167_nl;
  wire[0:0] nor_1168_nl;
  wire[0:0] mux_1931_nl;
  wire[0:0] mux_1932_nl;
  wire[0:0] mux_1933_nl;
  wire[0:0] mux_1934_nl;
  wire[0:0] mux_1081_nl;
  wire[0:0] or_2486_nl;
  wire[0:0] mux_1082_nl;
  wire[0:0] or_2490_nl;
  wire[0:0] mux_1083_nl;
  wire[0:0] or_2494_nl;
  wire[0:0] mux_1084_nl;
  wire[0:0] or_2498_nl;
  wire[0:0] mux_1091_nl;
  wire[0:0] nor_1151_nl;
  wire[0:0] nor_1153_nl;
  wire[0:0] mux_1090_nl;
  wire[0:0] or_2520_nl;
  wire[0:0] nand_136_nl;
  wire[0:0] mux_1098_nl;
  wire[0:0] or_2525_nl;
  wire[0:0] mux_1092_nl;
  wire[0:0] mux_1097_nl;
  wire[0:0] mux_1096_nl;
  wire[0:0] mux_1095_nl;
  wire[0:0] mux_1094_nl;
  wire[0:0] or_2531_nl;
  wire[0:0] or_860_nl;
  wire[0:0] mux_1101_nl;
  wire[0:0] mux_1108_nl;
  wire[0:0] nor_1143_nl;
  wire[0:0] nor_1145_nl;
  wire[0:0] mux_1107_nl;
  wire[0:0] or_2557_nl;
  wire[0:0] nand_140_nl;
  wire[0:0] mux_1115_nl;
  wire[0:0] or_2562_nl;
  wire[0:0] mux_1109_nl;
  wire[0:0] mux_1114_nl;
  wire[0:0] mux_1113_nl;
  wire[0:0] mux_1112_nl;
  wire[0:0] mux_1111_nl;
  wire[0:0] or_2568_nl;
  wire[0:0] or_889_nl;
  wire[0:0] mux_1118_nl;
  wire[0:0] mux_1125_nl;
  wire[0:0] nor_1135_nl;
  wire[0:0] nor_1137_nl;
  wire[0:0] mux_1124_nl;
  wire[0:0] or_2594_nl;
  wire[0:0] nand_144_nl;
  wire[0:0] mux_1132_nl;
  wire[0:0] or_2599_nl;
  wire[0:0] mux_1126_nl;
  wire[0:0] mux_1131_nl;
  wire[0:0] mux_1130_nl;
  wire[0:0] mux_1129_nl;
  wire[0:0] mux_1128_nl;
  wire[0:0] or_2605_nl;
  wire[0:0] or_926_nl;
  wire[0:0] mux_1135_nl;
  wire[0:0] mux_1143_nl;
  wire[0:0] nor_1127_nl;
  wire[0:0] nor_1129_nl;
  wire[0:0] mux_1142_nl;
  wire[0:0] or_2632_nl;
  wire[0:0] mux_1150_nl;
  wire[0:0] or_2637_nl;
  wire[0:0] mux_1144_nl;
  wire[0:0] mux_1149_nl;
  wire[0:0] mux_1148_nl;
  wire[0:0] mux_1147_nl;
  wire[0:0] mux_1146_nl;
  wire[0:0] or_2643_nl;
  wire[0:0] or_2638_nl;
  wire[0:0] mux_1153_nl;
  wire[0:0] mux_1156_nl;
  wire[0:0] mux_1154_nl;
  wire[0:0] nor_1123_nl;
  wire[0:0] or_2650_nl;
  wire[0:0] mux_1155_nl;
  wire[0:0] nor_1125_nl;
  wire[0:0] nor_1126_nl;
  wire[0:0] or_2656_nl;
  wire[0:0] mux_1157_nl;
  wire[0:0] mux_1160_nl;
  wire[0:0] mux_1158_nl;
  wire[0:0] nor_1119_nl;
  wire[0:0] nor_1120_nl;
  wire[0:0] mux_1159_nl;
  wire[0:0] nor_1121_nl;
  wire[0:0] nor_1122_nl;
  wire[0:0] or_2669_nl;
  wire[0:0] mux_1161_nl;
  wire[0:0] mux_1164_nl;
  wire[0:0] nor_1116_nl;
  wire[0:0] mux_1162_nl;
  wire[0:0] and_3198_nl;
  wire[0:0] mux_1163_nl;
  wire[0:0] nor_1117_nl;
  wire[0:0] nor_1118_nl;
  wire[0:0] or_2678_nl;
  wire[0:0] mux_1165_nl;
  wire[0:0] mux_1168_nl;
  wire[0:0] mux_1166_nl;
  wire[0:0] nor_1112_nl;
  wire[0:0] or_2685_nl;
  wire[0:0] mux_1167_nl;
  wire[0:0] nor_1114_nl;
  wire[0:0] nor_1115_nl;
  wire[0:0] or_2691_nl;
  wire[0:0] mux_1169_nl;
  wire[0:0] mux_2118_nl;
  wire[0:0] mux_2117_nl;
  wire[0:0] or_6073_nl;
  wire[4:0] inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_nl;
  wire[5:0] nl_inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_nl;
  wire[0:0] mux_1184_nl;
  wire[0:0] and_3191_nl;
  wire[0:0] mux_1183_nl;
  wire[0:0] and_3192_nl;
  wire[0:0] and_3193_nl;
  wire[0:0] mux_1941_nl;
  wire[0:0] mux_2120_nl;
  wire[0:0] mux_2119_nl;
  wire[0:0] or_6080_nl;
  wire[0:0] mux_1190_nl;
  wire[0:0] mux_1188_nl;
  wire[0:0] nor_1101_nl;
  wire[0:0] and_3380_nl;
  wire[0:0] mux_1189_nl;
  wire[0:0] nor_1103_nl;
  wire[0:0] nor_1104_nl;
  wire[0:0] mux_1942_nl;
  wire[0:0] mux_2122_nl;
  wire[0:0] mux_2121_nl;
  wire[0:0] or_6087_nl;
  wire[0:0] mux_1196_nl;
  wire[0:0] mux_1194_nl;
  wire[0:0] nor_1094_nl;
  wire[0:0] and_3378_nl;
  wire[0:0] mux_1195_nl;
  wire[0:0] nor_1096_nl;
  wire[0:0] nor_1097_nl;
  wire[0:0] mux_1198_nl;
  wire[0:0] mux_1197_nl;
  wire[0:0] or_2773_nl;
  wire[0:0] or_2771_nl;
  wire[0:0] mux_1201_nl;
  wire[0:0] mux_1199_nl;
  wire[0:0] nor_1090_nl;
  wire[0:0] and_3377_nl;
  wire[0:0] mux_1200_nl;
  wire[0:0] nor_1092_nl;
  wire[0:0] nor_1093_nl;
  wire[0:0] mux_1943_nl;
  wire[0:0] mux_2126_nl;
  wire[0:0] mux_2125_nl;
  wire[0:0] nor_1866_nl;
  wire[0:0] or_6101_nl;
  wire[0:0] mux_1208_nl;
  wire[0:0] and_3184_nl;
  wire[0:0] mux_1207_nl;
  wire[0:0] and_3375_nl;
  wire[0:0] mux_1211_nl;
  wire[0:0] or_2805_nl;
  wire[0:0] mux_1210_nl;
  wire[0:0] mux_1213_nl;
  wire[0:0] nor_1082_nl;
  wire[0:0] mux_1212_nl;
  wire[0:0] mux_1219_nl;
  wire[0:0] and_3182_nl;
  wire[0:0] mux_1218_nl;
  wire[0:0] and_3373_nl;
  wire[0:0] mux_1220_nl;
  wire[0:0] nor_1078_nl;
  wire[0:0] and_3181_nl;
  wire[0:0] mux_1221_nl;
  wire[0:0] nor_1076_nl;
  wire[0:0] nor_1077_nl;
  wire[0:0] mux_1222_nl;
  wire[0:0] nand_676_nl;
  wire[0:0] mux_1223_nl;
  wire[0:0] nor_1074_nl;
  wire[0:0] nor_1075_nl;
  wire[0:0] mux_1224_nl;
  wire[0:0] nor_1072_nl;
  wire[0:0] and_3180_nl;
  wire[0:0] mux_1225_nl;
  wire[0:0] nor_1070_nl;
  wire[0:0] nor_1071_nl;
  wire[0:0] mux_1226_nl;
  wire[0:0] nand_674_nl;
  wire[0:0] mux_1227_nl;
  wire[0:0] nor_1068_nl;
  wire[0:0] nor_1069_nl;
  wire[0:0] mux_1228_nl;
  wire[0:0] and_3178_nl;
  wire[0:0] and_3179_nl;
  wire[0:0] mux_1229_nl;
  wire[0:0] nor_1065_nl;
  wire[0:0] nor_1066_nl;
  wire[0:0] mux_1230_nl;
  wire[0:0] nand_672_nl;
  wire[0:0] mux_1231_nl;
  wire[0:0] nor_1063_nl;
  wire[0:0] nor_1064_nl;
  wire[0:0] mux_1232_nl;
  wire[0:0] and_3176_nl;
  wire[0:0] and_3177_nl;
  wire[0:0] mux_1233_nl;
  wire[0:0] nor_1061_nl;
  wire[0:0] nor_1062_nl;
  wire[0:0] mux_1234_nl;
  wire[0:0] nand_390_nl;
  wire[0:0] mux_1235_nl;
  wire[0:0] nor_1059_nl;
  wire[0:0] nor_1060_nl;
  wire[0:0] mux_1237_nl;
  wire[0:0] mux_1239_nl;
  wire[0:0] mux_1241_nl;
  wire[0:0] mux_1243_nl;
  wire[0:0] mux_1245_nl;
  wire[0:0] or_2923_nl;
  wire[0:0] mux_1244_nl;
  wire[0:0] mux_1246_nl;
  wire[0:0] or_2930_nl;
  wire[0:0] mux_1247_nl;
  wire[0:0] or_2934_nl;
  wire[0:0] mux_1248_nl;
  wire[0:0] mux_1249_nl;
  wire[0:0] nor_1049_nl;
  wire[0:0] mux_1251_nl;
  wire[0:0] mux_1250_nl;
  wire[0:0] or_2949_nl;
  wire[0:0] or_2952_nl;
  wire[0:0] mux_1252_nl;
  wire[0:0] mux_1253_nl;
  wire[0:0] nor_1046_nl;
  wire[0:0] mux_1255_nl;
  wire[0:0] mux_1254_nl;
  wire[0:0] or_2967_nl;
  wire[0:0] or_2970_nl;
  wire[0:0] mux_1257_nl;
  wire[0:0] or_2973_nl;
  wire[0:0] mux_1256_nl;
  wire[0:0] mux_1259_nl;
  wire[0:0] nand_166_nl;
  wire[0:0] mux_1258_nl;
  wire[0:0] nor_1042_nl;
  wire[0:0] nor_1043_nl;
  wire[0:0] mux_1260_nl;
  wire[0:0] or_2983_nl;
  wire[0:0] mux_1263_nl;
  wire[0:0] mux_1262_nl;
  wire[0:0] and_284_nl;
  wire[0:0] mux_1267_nl;
  wire[0:0] mux_1266_nl;
  wire[0:0] and_286_nl;
  wire[0:0] mux_1271_nl;
  wire[0:0] mux_1275_nl;
  wire[0:0] mux_1274_nl;
  wire[0:0] and_290_nl;
  wire[0:0] mux_1264_nl;
  wire[0:0] mux_1268_nl;
  wire[0:0] mux_1272_nl;
  wire[0:0] mux_1276_nl;
  wire[0:0] mux_1281_nl;
  wire[0:0] and_3173_nl;
  wire[0:0] mux_2192_nl;
  wire[0:0] nor_1040_nl;
  wire[0:0] and_3174_nl;
  wire[0:0] mux_2197_nl;
  wire[0:0] nor_1041_nl;
  wire[0:0] mux_1286_nl;
  wire[0:0] and_3171_nl;
  wire[0:0] mux_1282_nl;
  wire[0:0] nor_1038_nl;
  wire[0:0] and_3172_nl;
  wire[0:0] mux_1284_nl;
  wire[0:0] nor_1039_nl;
  wire[0:0] mux_1288_nl;
  wire[0:0] mux_1293_nl;
  wire[0:0] and_3167_nl;
  wire[0:0] mux_2191_nl;
  wire[0:0] nor_1036_nl;
  wire[0:0] and_3168_nl;
  wire[0:0] mux_2196_nl;
  wire[0:0] nor_1037_nl;
  wire[0:0] mux_1298_nl;
  wire[0:0] and_3165_nl;
  wire[0:0] mux_1294_nl;
  wire[0:0] nor_1034_nl;
  wire[0:0] and_3166_nl;
  wire[0:0] mux_1296_nl;
  wire[0:0] nor_1035_nl;
  wire[0:0] mux_1300_nl;
  wire[0:0] mux_1305_nl;
  wire[0:0] and_3161_nl;
  wire[0:0] mux_2190_nl;
  wire[0:0] nor_1032_nl;
  wire[0:0] and_3162_nl;
  wire[0:0] mux_2195_nl;
  wire[0:0] nor_1033_nl;
  wire[0:0] mux_1310_nl;
  wire[0:0] and_3159_nl;
  wire[0:0] mux_1306_nl;
  wire[0:0] nor_1030_nl;
  wire[0:0] and_3160_nl;
  wire[0:0] mux_1308_nl;
  wire[0:0] nor_1031_nl;
  wire[0:0] mux_1312_nl;
  wire[0:0] mux_1317_nl;
  wire[0:0] and_3155_nl;
  wire[0:0] mux_2189_nl;
  wire[0:0] nor_1028_nl;
  wire[0:0] and_3156_nl;
  wire[0:0] mux_2194_nl;
  wire[0:0] nor_1029_nl;
  wire[0:0] mux_1322_nl;
  wire[0:0] and_3153_nl;
  wire[0:0] mux_1318_nl;
  wire[0:0] nor_1026_nl;
  wire[0:0] and_3154_nl;
  wire[0:0] mux_1320_nl;
  wire[0:0] nor_1027_nl;
  wire[0:0] mux_1324_nl;
  wire[0:0] mux_882_nl;
  wire[0:0] mux_878_nl;
  wire[0:0] mux_875_nl;
  wire[0:0] mux_873_nl;
  wire[0:0] nand_93_nl;
  wire[0:0] mux_872_nl;
  wire[0:0] nor_1362_nl;
  wire[0:0] nor_1364_nl;
  wire[0:0] mux_881_nl;
  wire[0:0] mux_879_nl;
  wire[0:0] nor_1365_nl;
  wire[0:0] nor_1366_nl;
  wire[0:0] mux_880_nl;
  wire[0:0] nor_1367_nl;
  wire[0:0] mux_1325_nl;
  wire[0:0] and_3150_nl;
  wire[0:0] nor_1025_nl;
  wire[0:0] mux_1327_nl;
  wire[0:0] nor_1021_nl;
  wire[0:0] mux_1326_nl;
  wire[0:0] nand_378_nl;
  wire[0:0] nor_1022_nl;
  wire[0:0] mux_1329_nl;
  wire[0:0] nor_1018_nl;
  wire[0:0] mux_1328_nl;
  wire[0:0] nand_376_nl;
  wire[0:0] nor_1019_nl;
  wire[0:0] mux_1331_nl;
  wire[0:0] mux_1330_nl;
  wire[0:0] nor_1014_nl;
  wire[0:0] nor_1015_nl;
  wire[0:0] mux_1333_nl;
  wire[0:0] mux_1332_nl;
  wire[0:0] and_3371_nl;
  wire[0:0] nor_1010_nl;
  wire[0:0] nor_1011_nl;
  wire[0:0] and_2058_nl;
  wire[0:0] and_2060_nl;
  wire[0:0] or_5554_nl;
  wire[0:0] mux_1948_nl;
  wire[0:0] or_5132_nl;
  wire[0:0] mux_1949_nl;
  wire[0:0] or_5136_nl;
  wire[0:0] mux_2001_nl;
  wire[0:0] nor_1801_nl;
  wire[0:0] or_5835_nl;
  wire[0:0] mux_1342_nl;
  wire[0:0] mux_1337_nl;
  wire[0:0] or_3121_nl;
  wire[0:0] mux_1335_nl;
  wire[0:0] mux_1334_nl;
  wire[0:0] or_3116_nl;
  wire[0:0] or_3118_nl;
  wire[0:0] mux_1336_nl;
  wire[0:0] mux_1341_nl;
  wire[0:0] mux_1340_nl;
  wire[0:0] mux_1339_nl;
  wire[0:0] or_3130_nl;
  wire[0:0] mux_1952_nl;
  wire[0:0] mux_1884_nl;
  wire[0:0] mux_1883_nl;
  wire[0:0] and_994_nl;
  wire[0:0] nor_682_nl;
  wire[0:0] or_4372_nl;
  wire[0:0] or_5142_nl;
  wire[0:0] and_2082_nl;
  wire[0:0] and_2085_nl;
  wire[0:0] or_5558_nl;
  wire[0:0] mux_1953_nl;
  wire[0:0] nor_nl;
  wire[0:0] nor_1787_nl;
  wire[0:0] mux_2002_nl;
  wire[0:0] or_5834_nl;
  wire[0:0] mux_2003_nl;
  wire[0:0] or_nl;
  wire[0:0] inp_lookup_1_FpAdd_6U_10U_1_IsZero_6U_10U_8_or_nl;
  wire[0:0] inp_lookup_2_FpAdd_6U_10U_1_IsZero_6U_10U_8_or_nl;
  wire[0:0] inp_lookup_3_FpAdd_6U_10U_1_IsZero_6U_10U_8_or_nl;
  wire[0:0] inp_lookup_4_FpAdd_6U_10U_1_IsZero_6U_10U_8_or_nl;
  wire[0:0] mux_1345_nl;
  wire[0:0] mux_1343_nl;
  wire[0:0] nor_1005_nl;
  wire[0:0] nor_1006_nl;
  wire[0:0] nor_1007_nl;
  wire[0:0] mux_1344_nl;
  wire[0:0] mux_1346_nl;
  wire[0:0] nor_1003_nl;
  wire[0:0] nor_1004_nl;
  wire[0:0] mux_1350_nl;
  wire[0:0] mux_1348_nl;
  wire[0:0] mux_1349_nl;
  wire[0:0] mux_1351_nl;
  wire[0:0] mux_1352_nl;
  wire[0:0] FpMul_6U_10U_1_o_mant_or_nl;
  wire[0:0] FpMul_6U_10U_1_o_mant_and_8_nl;
  wire[0:0] mux_2129_nl;
  wire[0:0] nor_1864_nl;
  wire[0:0] mux_2128_nl;
  wire[0:0] or_6120_nl;
  wire[0:0] mux_2127_nl;
  wire[0:0] nor_1865_nl;
  wire[0:0] mux_1359_nl;
  wire[0:0] mux_1357_nl;
  wire[0:0] and_3370_nl;
  wire[0:0] and_3140_nl;
  wire[0:0] nor_996_nl;
  wire[0:0] mux_1358_nl;
  wire[0:0] mux_1361_nl;
  wire[0:0] nor_992_nl;
  wire[0:0] and_3139_nl;
  wire[0:0] mux_1360_nl;
  wire[0:0] nor_993_nl;
  wire[0:0] nor_994_nl;
  wire[0:0] mux_1365_nl;
  wire[0:0] mux_1363_nl;
  wire[0:0] nor_988_nl;
  wire[0:0] nor_989_nl;
  wire[0:0] nor_990_nl;
  wire[0:0] mux_1364_nl;
  wire[0:0] mux_1366_nl;
  wire[0:0] nor_986_nl;
  wire[0:0] nor_987_nl;
  wire[0:0] IsNaN_6U_23U_2_IsNaN_6U_23U_2_nand_nl;
  wire[0:0] IsNaN_6U_23U_2_IsNaN_6U_23U_2_nand_1_nl;
  wire[0:0] IsNaN_6U_23U_2_IsNaN_6U_23U_2_nand_2_nl;
  wire[0:0] IsNaN_6U_23U_2_IsNaN_6U_23U_2_nand_3_nl;
  wire[0:0] mux_1368_nl;
  wire[0:0] mux_1369_nl;
  wire[0:0] mux_1370_nl;
  wire[0:0] mux_1371_nl;
  wire[0:0] mux_1372_nl;
  wire[0:0] mux_1373_nl;
  wire[0:0] mux_1374_nl;
  wire[0:0] mux_1375_nl;
  wire[0:0] mux_1384_nl;
  wire[0:0] and_3137_nl;
  wire[0:0] mux_1379_nl;
  wire[0:0] or_3241_nl;
  wire[0:0] and_3138_nl;
  wire[0:0] mux_1383_nl;
  wire[0:0] or_3246_nl;
  wire[0:0] mux_1393_nl;
  wire[0:0] and_3135_nl;
  wire[0:0] mux_1388_nl;
  wire[0:0] or_3252_nl;
  wire[0:0] and_3136_nl;
  wire[0:0] mux_1392_nl;
  wire[0:0] or_3257_nl;
  wire[0:0] mux_1402_nl;
  wire[0:0] and_3133_nl;
  wire[0:0] mux_1397_nl;
  wire[0:0] or_3263_nl;
  wire[0:0] and_3134_nl;
  wire[0:0] mux_1401_nl;
  wire[0:0] or_3268_nl;
  wire[0:0] mux_1411_nl;
  wire[0:0] and_3131_nl;
  wire[0:0] mux_1406_nl;
  wire[0:0] or_3274_nl;
  wire[0:0] and_3132_nl;
  wire[0:0] mux_1410_nl;
  wire[0:0] or_3279_nl;
  wire[0:0] mux_1376_nl;
  wire[0:0] mux_1385_nl;
  wire[0:0] mux_1394_nl;
  wire[0:0] mux_1403_nl;
  wire[0:0] mux_1419_nl;
  wire[0:0] mux_1414_nl;
  wire[0:0] mux_1412_nl;
  wire[0:0] or_3282_nl;
  wire[0:0] nand_198_nl;
  wire[0:0] mux_1413_nl;
  wire[0:0] nor_975_nl;
  wire[0:0] nor_976_nl;
  wire[0:0] nand_199_nl;
  wire[0:0] mux_1418_nl;
  wire[0:0] or_3292_nl;
  wire[0:0] mux_1420_nl;
  wire[0:0] and_3129_nl;
  wire[0:0] mux_1428_nl;
  wire[0:0] mux_1423_nl;
  wire[0:0] mux_1421_nl;
  wire[0:0] or_3298_nl;
  wire[0:0] nand_200_nl;
  wire[0:0] mux_1422_nl;
  wire[0:0] nor_973_nl;
  wire[0:0] nor_974_nl;
  wire[0:0] nand_201_nl;
  wire[0:0] mux_1427_nl;
  wire[0:0] or_3308_nl;
  wire[0:0] mux_1436_nl;
  wire[0:0] mux_1431_nl;
  wire[0:0] mux_1429_nl;
  wire[0:0] or_3311_nl;
  wire[0:0] nand_202_nl;
  wire[0:0] mux_1430_nl;
  wire[0:0] nor_971_nl;
  wire[0:0] nor_972_nl;
  wire[0:0] nand_203_nl;
  wire[0:0] mux_1435_nl;
  wire[0:0] or_3321_nl;
  wire[0:0] mux_1444_nl;
  wire[0:0] mux_1439_nl;
  wire[0:0] mux_1437_nl;
  wire[0:0] or_3324_nl;
  wire[0:0] nand_204_nl;
  wire[0:0] mux_1438_nl;
  wire[0:0] nor_969_nl;
  wire[0:0] nor_970_nl;
  wire[0:0] nand_205_nl;
  wire[0:0] mux_1443_nl;
  wire[0:0] or_3334_nl;
  wire[0:0] mux_1446_nl;
  wire[0:0] nand_206_nl;
  wire[0:0] mux_1448_nl;
  wire[0:0] or_3342_nl;
  wire[0:0] mux_1450_nl;
  wire[0:0] or_3345_nl;
  wire[0:0] mux_1452_nl;
  wire[0:0] or_3348_nl;
  wire[0:0] mux_1451_nl;
  wire[0:0] mux_1455_nl;
  wire[0:0] and_3127_nl;
  wire[0:0] mux_1453_nl;
  wire[0:0] and_3128_nl;
  wire[0:0] mux_1454_nl;
  wire[0:0] or_3350_nl;
  wire[0:0] mux_1458_nl;
  wire[0:0] and_3125_nl;
  wire[0:0] mux_1456_nl;
  wire[0:0] or_3353_nl;
  wire[0:0] and_3126_nl;
  wire[0:0] mux_1457_nl;
  wire[0:0] mux_1461_nl;
  wire[0:0] mux_1459_nl;
  wire[0:0] or_3356_nl;
  wire[0:0] nand_211_nl;
  wire[0:0] mux_1460_nl;
  wire[0:0] mux_1464_nl;
  wire[0:0] nor_967_nl;
  wire[0:0] mux_1462_nl;
  wire[0:0] nor_968_nl;
  wire[0:0] inp_lookup_1_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_nl;
  wire[0:0] mux_1467_nl;
  wire[0:0] nand_214_nl;
  wire[0:0] mux_1466_nl;
  wire[0:0] or_3363_nl;
  wire[0:0] mux_1465_nl;
  wire[0:0] inp_lookup_2_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_nl;
  wire[0:0] mux_1470_nl;
  wire[0:0] nand_215_nl;
  wire[0:0] mux_1469_nl;
  wire[0:0] or_3366_nl;
  wire[0:0] mux_1468_nl;
  wire[0:0] inp_lookup_3_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_nl;
  wire[0:0] mux_1473_nl;
  wire[0:0] nand_216_nl;
  wire[0:0] mux_1472_nl;
  wire[0:0] or_3369_nl;
  wire[0:0] mux_1471_nl;
  wire[0:0] inp_lookup_4_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_nl;
  wire[0:0] mux_1475_nl;
  wire[0:0] nand_217_nl;
  wire[0:0] mux_1474_nl;
  wire[0:0] nor_963_nl;
  wire[0:0] nor_965_nl;
  wire[0:0] mux_2206_nl;
  wire[0:0] mux_1482_nl;
  wire[0:0] mux_1478_nl;
  wire[0:0] mux_1481_nl;
  wire[0:0] mux_1488_nl;
  wire[0:0] mux_1484_nl;
  wire[0:0] mux_1487_nl;
  wire[0:0] mux_2207_nl;
  wire[0:0] mux_1495_nl;
  wire[0:0] mux_1491_nl;
  wire[0:0] mux_1494_nl;
  wire[0:0] mux_1501_nl;
  wire[0:0] mux_1497_nl;
  wire[0:0] mux_1500_nl;
  wire[0:0] or_3417_nl;
  wire[0:0] mux_2208_nl;
  wire[0:0] mux_1508_nl;
  wire[0:0] mux_1504_nl;
  wire[0:0] mux_1507_nl;
  wire[0:0] mux_1514_nl;
  wire[0:0] mux_1510_nl;
  wire[0:0] mux_1513_nl;
  wire[0:0] mux_1479_nl;
  wire[0:0] mux_1521_nl;
  wire[0:0] mux_1517_nl;
  wire[0:0] mux_1520_nl;
  wire[0:0] mux_1527_nl;
  wire[0:0] mux_1523_nl;
  wire[0:0] mux_1526_nl;
  wire[0:0] mux_1529_nl;
  wire[0:0] mux_1531_nl;
  wire[0:0] mux_1535_nl;
  wire[0:0] mux_1534_nl;
  wire[0:0] mux_1539_nl;
  wire[0:0] mux_1538_nl;
  wire[0:0] mux_1540_nl;
  wire[0:0] or_3482_nl;
  wire[0:0] and_3550_nl;
  wire[0:0] nor_1756_nl;
  wire[0:0] mux_1547_nl;
  wire[0:0] and_4212_nl;
  wire[0:0] and_4214_nl;
  wire[0:0] mux_2198_nl;
  wire[0:0] nor_1758_nl;
  wire[0:0] mux_1548_nl;
  wire[0:0] or_3495_nl;
  wire[0:0] and_3552_nl;
  wire[0:0] mux_1555_nl;
  wire[0:0] and_4213_nl;
  wire[0:0] and_4215_nl;
  wire[0:0] mux_2199_nl;
  wire[0:0] nor_1754_nl;
  wire[0:0] mux_1556_nl;
  wire[0:0] or_3508_nl;
  wire[0:0] and_3554_nl;
  wire[0:0] mux_1557_nl;
  wire[0:0] or_3510_nl;
  wire[0:0] and_3556_nl;
  wire[3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_mux_44_nl;
  wire[2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_15_nl;
  wire[2:0] inp_lookup_4_FpExpoWidthInc_6U_8U_23U_0U_1U_1_else_acc_nl;
  wire[3:0] nl_inp_lookup_4_FpExpoWidthInc_6U_8U_23U_0U_1U_1_else_acc_nl;
  wire[0:0] IsZero_6U_23U_1_aelse_IsZero_6U_23U_1_or_3_nl;
  wire[0:0] IsInf_6U_23U_1_aelse_mux_7_nl;
  wire[0:0] or_5264_nl;
  wire[3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_mux_31_nl;
  wire[2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_10_nl;
  wire[2:0] inp_lookup_3_FpExpoWidthInc_6U_8U_23U_0U_1U_1_else_acc_nl;
  wire[3:0] nl_inp_lookup_3_FpExpoWidthInc_6U_8U_23U_0U_1U_1_else_acc_nl;
  wire[0:0] IsZero_6U_23U_1_aelse_IsZero_6U_23U_1_or_2_nl;
  wire[0:0] IsInf_6U_23U_1_aelse_mux_5_nl;
  wire[0:0] or_5260_nl;
  wire[3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_mux_18_nl;
  wire[2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_5_nl;
  wire[2:0] inp_lookup_2_FpExpoWidthInc_6U_8U_23U_0U_1U_1_else_acc_nl;
  wire[3:0] nl_inp_lookup_2_FpExpoWidthInc_6U_8U_23U_0U_1U_1_else_acc_nl;
  wire[0:0] IsZero_6U_23U_1_aelse_IsZero_6U_23U_1_or_1_nl;
  wire[0:0] IsInf_6U_23U_1_aelse_mux_3_nl;
  wire[0:0] or_5256_nl;
  wire[3:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_mux_48_nl;
  wire[2:0] FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_nl;
  wire[2:0] inp_lookup_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_else_acc_nl;
  wire[3:0] nl_inp_lookup_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_else_acc_nl;
  wire[0:0] IsZero_6U_23U_1_aelse_IsZero_6U_23U_1_or_nl;
  wire[0:0] IsInf_6U_23U_1_aelse_mux_1_nl;
  wire[0:0] or_5251_nl;
  wire[0:0] mux_1564_nl;
  wire[0:0] mux_1567_nl;
  wire[0:0] mux_1570_nl;
  wire[0:0] mux_1573_nl;
  wire[0:0] mux_1574_nl;
  wire[0:0] mux_1579_nl;
  wire[0:0] or_3533_nl;
  wire[0:0] mux_1580_nl;
  wire[0:0] or_3537_nl;
  wire[0:0] mux_1581_nl;
  wire[0:0] or_3541_nl;
  wire[0:0] mux_1582_nl;
  wire[0:0] or_3545_nl;
  wire[0:0] mux_1583_nl;
  wire[0:0] mux_1584_nl;
  wire[0:0] mux_1585_nl;
  wire[0:0] mux_1588_nl;
  wire[0:0] mux_1590_nl;
  wire[0:0] mux_1592_nl;
  wire[0:0] mux_1595_nl;
  wire[0:0] mux_1597_nl;
  wire[0:0] mux_1598_nl;
  wire[0:0] mux_1599_nl;
  wire[0:0] mux_1600_nl;
  wire[0:0] mux_1601_nl;
  wire[0:0] mux_1602_nl;
  wire[0:0] IsZero_6U_10U_1_IsZero_6U_10U_1_and_1_nl;
  wire[0:0] IsZero_6U_10U_1_IsZero_6U_10U_1_and_3_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_46_nl;
  wire[0:0] mux_1605_nl;
  wire[0:0] nor_921_nl;
  wire[0:0] nor_923_nl;
  wire[0:0] mux_1604_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_45_nl;
  wire[0:0] mux_1608_nl;
  wire[0:0] nor_917_nl;
  wire[0:0] nor_919_nl;
  wire[0:0] mux_1607_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_44_nl;
  wire[0:0] mux_1612_nl;
  wire[0:0] nor_911_nl;
  wire[0:0] mux_1611_nl;
  wire[0:0] nor_913_nl;
  wire[0:0] mux_1610_nl;
  wire[0:0] and_3394_nl;
  wire[0:0] nor_915_nl;
  wire[0:0] or_3596_nl;
  wire[0:0] mux_1613_nl;
  wire[0:0] mux_1614_nl;
  wire[0:0] mux_1615_nl;
  wire[0:0] mux_1616_nl;
  wire[0:0] mux_1617_nl;
  wire[0:0] mux_1618_nl;
  wire[0:0] mux_1619_nl;
  wire[0:0] mux_1620_nl;
  wire[0:0] mux_1622_nl;
  wire[0:0] mux_1624_nl;
  wire[0:0] mux_1629_nl;
  wire[0:0] mux_1632_nl;
  wire[0:0] mux_1633_nl;
  wire[0:0] mux_1634_nl;
  wire[0:0] mux_1635_nl;
  wire[0:0] mux_1636_nl;
  wire[0:0] mux_1637_nl;
  wire[0:0] IsZero_6U_10U_5_IsZero_6U_10U_5_and_nl;
  wire[0:0] IsZero_6U_10U_1_IsZero_6U_10U_1_and_nl;
  wire[0:0] IsZero_6U_10U_5_IsZero_6U_10U_5_and_2_nl;
  wire[0:0] IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_nl;
  wire[0:0] mux_1640_nl;
  wire[0:0] nor_902_nl;
  wire[0:0] mux_1638_nl;
  wire[0:0] mux_1639_nl;
  wire[0:0] nor_907_nl;
  wire[0:0] or_3645_nl;
  wire[0:0] mux_1643_nl;
  wire[0:0] nor_895_nl;
  wire[0:0] mux_1641_nl;
  wire[0:0] mux_1642_nl;
  wire[0:0] nor_900_nl;
  wire[0:0] or_3660_nl;
  wire[0:0] mux_1646_nl;
  wire[0:0] nor_889_nl;
  wire[0:0] mux_1644_nl;
  wire[0:0] mux_1645_nl;
  wire[0:0] nor_893_nl;
  wire[0:0] or_3674_nl;
  wire[0:0] mux_1647_nl;
  wire[0:0] mux_1648_nl;
  wire[0:0] mux_1649_nl;
  wire[0:0] mux_1650_nl;
  wire[0:0] mux_1652_nl;
  wire[0:0] mux_1654_nl;
  wire[0:0] mux_1656_nl;
  wire[0:0] mux_1658_nl;
  wire[0:0] mux_1660_nl;
  wire[0:0] mux_1662_nl;
  wire[0:0] mux_1664_nl;
  wire[0:0] mux_1666_nl;
  wire[0:0] mux_1667_nl;
  wire[0:0] and_3089_nl;
  wire[0:0] mux_1668_nl;
  wire[0:0] mux_1669_nl;
  wire[0:0] mux_1670_nl;
  wire[0:0] mux_1671_nl;
  wire[0:0] mux_1673_nl;
  wire[0:0] mux_1675_nl;
  wire[0:0] mux_1677_nl;
  wire[0:0] mux_1679_nl;
  wire[0:0] IsNaN_6U_10U_6_IsNaN_6U_10U_6_nor_nl;
  wire[0:0] IsNaN_6U_10U_6_IsNaN_6U_10U_6_nor_1_nl;
  wire[0:0] IsNaN_6U_10U_6_IsNaN_6U_10U_6_nor_2_nl;
  wire[0:0] IsNaN_6U_10U_6_IsNaN_6U_10U_6_nor_3_nl;
  wire[0:0] mux_1682_nl;
  wire[0:0] nor_881_nl;
  wire[0:0] mux_1680_nl;
  wire[0:0] nand_320_nl;
  wire[0:0] mux_1681_nl;
  wire[0:0] nor_883_nl;
  wire[0:0] or_3742_nl;
  wire[0:0] mux_1685_nl;
  wire[0:0] nor_876_nl;
  wire[0:0] mux_1683_nl;
  wire[0:0] nand_318_nl;
  wire[0:0] mux_1684_nl;
  wire[0:0] nor_879_nl;
  wire[0:0] or_3753_nl;
  wire[0:0] mux_1688_nl;
  wire[0:0] nor_871_nl;
  wire[0:0] mux_1686_nl;
  wire[0:0] nand_317_nl;
  wire[0:0] mux_1687_nl;
  wire[0:0] nor_874_nl;
  wire[0:0] or_3764_nl;
  wire[0:0] mux_1689_nl;
  wire[0:0] and_336_nl;
  wire[0:0] mux_1691_nl;
  wire[0:0] and_337_nl;
  wire[0:0] mux_1692_nl;
  wire[0:0] and_338_nl;
  wire[0:0] mux_1693_nl;
  wire[0:0] and_339_nl;
  wire[0:0] mux_1697_nl;
  wire[0:0] mux_1695_nl;
  wire[0:0] mux_1696_nl;
  wire[0:0] mux_1703_nl;
  wire[0:0] and_3084_nl;
  wire[0:0] mux_1701_nl;
  wire[0:0] nor_860_nl;
  wire[0:0] mux_1700_nl;
  wire[0:0] or_5649_nl;
  wire[0:0] nor_862_nl;
  wire[0:0] mux_1699_nl;
  wire[0:0] or_3788_nl;
  wire[0:0] or_3789_nl;
  wire[0:0] and_3085_nl;
  wire[0:0] mux_1702_nl;
  wire[0:0] nor_864_nl;
  wire[0:0] nor_865_nl;
  wire[0:0] mux_1711_nl;
  wire[0:0] mux_1709_nl;
  wire[0:0] mux_1705_nl;
  wire[0:0] mux_1708_nl;
  wire[0:0] mux_1706_nl;
  wire[0:0] or_3798_nl;
  wire[0:0] mux_1707_nl;
  wire[0:0] or_3809_nl;
  wire[0:0] nand_226_nl;
  wire[0:0] mux_1710_nl;
  wire[0:0] nor_853_nl;
  wire[0:0] nor_854_nl;
  wire[0:0] mux_1719_nl;
  wire[0:0] mux_1717_nl;
  wire[0:0] or_3817_nl;
  wire[0:0] mux_1716_nl;
  wire[0:0] mux_1714_nl;
  wire[0:0] mux_1713_nl;
  wire[0:0] or_3828_nl;
  wire[0:0] mux_1715_nl;
  wire[0:0] or_3825_nl;
  wire[0:0] or_3827_nl;
  wire[0:0] nor_600_nl;
  wire[0:0] nand_227_nl;
  wire[0:0] mux_1718_nl;
  wire[0:0] nor_845_nl;
  wire[0:0] nor_846_nl;
  wire[0:0] mux_1729_nl;
  wire[0:0] nor_836_nl;
  wire[0:0] mux_1725_nl;
  wire[0:0] mux_1721_nl;
  wire[0:0] mux_1720_nl;
  wire[0:0] or_3836_nl;
  wire[0:0] mux_1724_nl;
  wire[0:0] mux_1722_nl;
  wire[0:0] or_3840_nl;
  wire[0:0] or_3839_nl;
  wire[0:0] mux_1723_nl;
  wire[0:0] or_3843_nl;
  wire[0:0] mux_1728_nl;
  wire[0:0] mux_1726_nl;
  wire[0:0] nor_839_nl;
  wire[0:0] nor_840_nl;
  wire[0:0] nor_841_nl;
  wire[0:0] mux_1727_nl;
  wire[0:0] or_3853_nl;
  wire[0:0] mux_1731_nl;
  wire[0:0] mux_1733_nl;
  wire[0:0] mux_1735_nl;
  wire[0:0] mux_1737_nl;
  wire[0:0] mux_1744_nl;
  wire[0:0] nor_833_nl;
  wire[0:0] nor_1944_nl;
  wire[0:0] mux_1742_nl;
  wire[0:0] or_3867_nl;
  wire[0:0] or_3870_nl;
  wire[0:0] mux_1752_nl;
  wire[0:0] mux_1746_nl;
  wire[0:0] mux_1745_nl;
  wire[0:0] nor_825_nl;
  wire[0:0] nor_826_nl;
  wire[0:0] and_3081_nl;
  wire[0:0] nor_828_nl;
  wire[0:0] nor_1953_nl;
  wire[0:0] mux_1750_nl;
  wire[0:0] mux_1749_nl;
  wire[0:0] mux_1748_nl;
  wire[0:0] mux_1747_nl;
  wire[0:0] nand_779_nl;
  wire[0:0] mux_1759_nl;
  wire[0:0] nor_822_nl;
  wire[0:0] nor_1939_nl;
  wire[0:0] mux_1757_nl;
  wire[0:0] or_3895_nl;
  wire[0:0] or_3898_nl;
  wire[0:0] mux_1767_nl;
  wire[0:0] mux_1761_nl;
  wire[0:0] mux_1760_nl;
  wire[0:0] nor_814_nl;
  wire[0:0] nor_815_nl;
  wire[0:0] and_3079_nl;
  wire[0:0] nor_817_nl;
  wire[0:0] nor_1952_nl;
  wire[0:0] mux_1765_nl;
  wire[0:0] mux_1764_nl;
  wire[0:0] mux_1763_nl;
  wire[0:0] mux_1762_nl;
  wire[0:0] nand_778_nl;
  wire[0:0] mux_1774_nl;
  wire[0:0] nor_811_nl;
  wire[0:0] nor_1935_nl;
  wire[0:0] mux_1772_nl;
  wire[0:0] or_3923_nl;
  wire[0:0] or_3926_nl;
  wire[0:0] mux_1782_nl;
  wire[0:0] mux_1776_nl;
  wire[0:0] mux_1775_nl;
  wire[0:0] nor_803_nl;
  wire[0:0] nor_804_nl;
  wire[0:0] and_3077_nl;
  wire[0:0] nor_806_nl;
  wire[0:0] nor_1951_nl;
  wire[0:0] mux_1780_nl;
  wire[0:0] mux_1779_nl;
  wire[0:0] mux_1778_nl;
  wire[0:0] mux_1777_nl;
  wire[0:0] nand_777_nl;
  wire[0:0] mux_1789_nl;
  wire[0:0] nor_800_nl;
  wire[0:0] nor_1931_nl;
  wire[0:0] mux_1787_nl;
  wire[0:0] or_3951_nl;
  wire[0:0] or_3954_nl;
  wire[0:0] mux_1797_nl;
  wire[0:0] mux_1791_nl;
  wire[0:0] mux_1790_nl;
  wire[0:0] nor_792_nl;
  wire[0:0] nor_793_nl;
  wire[0:0] and_3075_nl;
  wire[0:0] nor_795_nl;
  wire[0:0] nor_1954_nl;
  wire[0:0] mux_1795_nl;
  wire[0:0] mux_1794_nl;
  wire[0:0] mux_1793_nl;
  wire[0:0] mux_1792_nl;
  wire[0:0] nand_780_nl;
  wire[0:0] mux_1802_nl;
  wire[0:0] or_5648_nl;
  wire[0:0] mux_1798_nl;
  wire[0:0] nor_791_nl;
  wire[0:0] mux_1801_nl;
  wire[0:0] or_3978_nl;
  wire[0:0] mux_1799_nl;
  wire[0:0] mux_1800_nl;
  wire[0:0] mux_1805_nl;
  wire[0:0] mux_1808_nl;
  wire[0:0] mux_1810_nl;
  wire[0:0] mux_1812_nl;
  wire[0:0] mux_1814_nl;
  wire[0:0] mux_1816_nl;
  wire[0:0] mux_1818_nl;
  wire[0:0] mux_1820_nl;
  wire[0:0] mux_1824_nl;
  wire[0:0] mux_1822_nl;
  wire[0:0] mux_1823_nl;
  wire[0:0] mux_1828_nl;
  wire[0:0] mux_1826_nl;
  wire[0:0] mux_1827_nl;
  wire[0:0] mux_1831_nl;
  wire[0:0] mux_1829_nl;
  wire[0:0] or_4004_nl;
  wire[0:0] mux_1830_nl;
  wire[0:0] or_4005_nl;
  wire[0:0] inp_lookup_4_IntShiftRight_69U_6U_32U_obits_fixed_and_nl;
  wire[0:0] mux_1833_nl;
  wire[0:0] nand_236_nl;
  wire[0:0] inp_lookup_3_IntShiftRight_69U_6U_32U_obits_fixed_and_nl;
  wire[0:0] mux_1835_nl;
  wire[0:0] or_4013_nl;
  wire[0:0] inp_lookup_2_IntShiftRight_69U_6U_32U_obits_fixed_and_nl;
  wire[0:0] mux_1837_nl;
  wire[0:0] nand_237_nl;
  wire[0:0] inp_lookup_1_IntShiftRight_69U_6U_32U_obits_fixed_and_nl;
  wire[0:0] mux_1840_nl;
  wire[0:0] nand_238_nl;
  wire[0:0] inp_lookup_4_IsZero_6U_10U_1_IsZero_6U_10U_1_nor_nl;
  wire[0:0] inp_lookup_1_IntShiftRight_69U_6U_32U_obits_fixed_or_nl;
  wire[0:0] inp_lookup_1_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_nl;
  wire[0:0] mux_1845_nl;
  wire[0:0] mux_1842_nl;
  wire[0:0] mux_1841_nl;
  wire[0:0] nor_782_nl;
  wire[0:0] mux_1844_nl;
  wire[0:0] mux_1843_nl;
  wire[0:0] nor_783_nl;
  wire[0:0] inp_lookup_2_IntShiftRight_69U_6U_32U_obits_fixed_or_nl;
  wire[0:0] inp_lookup_2_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_nl;
  wire[0:0] mux_1850_nl;
  wire[0:0] mux_1847_nl;
  wire[0:0] mux_1846_nl;
  wire[0:0] nor_776_nl;
  wire[0:0] mux_1849_nl;
  wire[0:0] mux_1848_nl;
  wire[0:0] nor_777_nl;
  wire[0:0] inp_lookup_3_IntShiftRight_69U_6U_32U_obits_fixed_or_nl;
  wire[0:0] inp_lookup_3_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_nl;
  wire[0:0] mux_1855_nl;
  wire[0:0] mux_1852_nl;
  wire[0:0] mux_1851_nl;
  wire[0:0] nor_770_nl;
  wire[0:0] mux_1854_nl;
  wire[0:0] mux_1853_nl;
  wire[0:0] nor_771_nl;
  wire[0:0] inp_lookup_4_IntShiftRight_69U_6U_32U_obits_fixed_or_nl;
  wire[0:0] inp_lookup_4_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_nl;
  wire[0:0] mux_1860_nl;
  wire[0:0] mux_1857_nl;
  wire[0:0] mux_1856_nl;
  wire[0:0] nor_764_nl;
  wire[0:0] mux_1859_nl;
  wire[0:0] mux_1858_nl;
  wire[0:0] nor_765_nl;
  wire[35:0] inp_lookup_1_else_else_a0_acc_nl;
  wire[36:0] nl_inp_lookup_1_else_else_a0_acc_nl;
  wire[33:0] inp_lookup_1_if_else_a_acc_nl;
  wire[34:0] nl_inp_lookup_1_if_else_a_acc_nl;
  wire[31:0] inp_lookup_if_else_ob_acc_8_nl;
  wire[32:0] nl_inp_lookup_if_else_ob_acc_8_nl;
  wire[32:0] inp_lookup_if_else_ob_acc_nl;
  wire[33:0] nl_inp_lookup_if_else_ob_acc_nl;
  wire[0:0] and_2521_nl;
  wire[0:0] mux_1972_nl;
  wire[0:0] mux_1973_nl;
  wire[0:0] mux_1861_nl;
  wire[0:0] nor_761_nl;
  wire[0:0] nor_762_nl;
  wire[35:0] inp_lookup_2_else_else_a0_acc_nl;
  wire[36:0] nl_inp_lookup_2_else_else_a0_acc_nl;
  wire[33:0] inp_lookup_2_if_else_a_acc_nl;
  wire[34:0] nl_inp_lookup_2_if_else_a_acc_nl;
  wire[31:0] inp_lookup_if_else_ob_acc_9_nl;
  wire[32:0] nl_inp_lookup_if_else_ob_acc_9_nl;
  wire[32:0] inp_lookup_if_else_ob_acc_2_nl;
  wire[33:0] nl_inp_lookup_if_else_ob_acc_2_nl;
  wire[0:0] and_2524_nl;
  wire[0:0] mux_1974_nl;
  wire[0:0] mux_1975_nl;
  wire[0:0] mux_1862_nl;
  wire[0:0] nor_759_nl;
  wire[0:0] nor_760_nl;
  wire[35:0] inp_lookup_3_else_else_a0_acc_nl;
  wire[36:0] nl_inp_lookup_3_else_else_a0_acc_nl;
  wire[33:0] inp_lookup_3_if_else_a_acc_nl;
  wire[34:0] nl_inp_lookup_3_if_else_a_acc_nl;
  wire[31:0] inp_lookup_if_else_ob_acc_10_nl;
  wire[32:0] nl_inp_lookup_if_else_ob_acc_10_nl;
  wire[32:0] inp_lookup_if_else_ob_acc_4_nl;
  wire[33:0] nl_inp_lookup_if_else_ob_acc_4_nl;
  wire[0:0] and_2527_nl;
  wire[0:0] mux_1976_nl;
  wire[0:0] mux_1977_nl;
  wire[0:0] mux_1863_nl;
  wire[0:0] nor_757_nl;
  wire[0:0] and_3058_nl;
  wire[35:0] inp_lookup_4_else_else_a0_acc_nl;
  wire[36:0] nl_inp_lookup_4_else_else_a0_acc_nl;
  wire[33:0] inp_lookup_4_if_else_a_acc_nl;
  wire[34:0] nl_inp_lookup_4_if_else_a_acc_nl;
  wire[31:0] inp_lookup_if_else_ob_acc_11_nl;
  wire[32:0] nl_inp_lookup_if_else_ob_acc_11_nl;
  wire[32:0] inp_lookup_if_else_ob_acc_6_nl;
  wire[33:0] nl_inp_lookup_if_else_ob_acc_6_nl;
  wire[0:0] and_2530_nl;
  wire[0:0] mux_1978_nl;
  wire[0:0] mux_1979_nl;
  wire[0:0] mux_1864_nl;
  wire[0:0] nor_755_nl;
  wire[0:0] and_nl;
  wire[0:0] and_518_nl;
  wire[0:0] and_522_nl;
  wire[0:0] and_524_nl;
  wire[0:0] and_528_nl;
  wire[0:0] and_530_nl;
  wire[0:0] and_534_nl;
  wire[0:0] and_536_nl;
  wire[0:0] and_540_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_nl;
  wire[8:0] FpAdd_8U_23U_is_a_greater_acc_nl;
  wire[10:0] nl_FpAdd_8U_23U_is_a_greater_acc_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_mux_2_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_mux1h_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_and_2_nl;
  wire[0:0] IsZero_5U_10U_3_aelse_not_27_nl;
  wire[5:0] inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_nl;
  wire[6:0] nl_inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_nl;
  wire[8:0] FpAdd_8U_23U_is_a_greater_acc_1_nl;
  wire[10:0] nl_FpAdd_8U_23U_is_a_greater_acc_1_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_mux_7_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_1_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_mux1h_1_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_and_5_nl;
  wire[0:0] IsZero_5U_10U_3_aelse_not_26_nl;
  wire[5:0] inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_nl;
  wire[6:0] nl_inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_nl;
  wire[23:0] FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_nl;
  wire[25:0] nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_nl;
  wire[8:0] FpAdd_8U_23U_is_a_greater_acc_2_nl;
  wire[10:0] nl_FpAdd_8U_23U_is_a_greater_acc_2_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_mux_12_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_2_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_mux1h_2_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_and_8_nl;
  wire[0:0] IsZero_5U_10U_3_aelse_not_25_nl;
  wire[5:0] inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_nl;
  wire[6:0] nl_inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_mux_17_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_3_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_mux1h_3_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_and_11_nl;
  wire[0:0] IsZero_5U_10U_3_aelse_not_24_nl;
  wire[5:0] inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_nl;
  wire[6:0] nl_inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_nl;
  wire[0:0] mux_75_nl;
  wire[6:0] inp_lookup_1_FpMul_6U_10U_2_else_2_if_acc_nl;
  wire[7:0] nl_inp_lookup_1_FpMul_6U_10U_2_else_2_if_acc_nl;
  wire[6:0] inp_lookup_1_FpMul_6U_10U_2_else_2_acc_1_nl;
  wire[7:0] nl_inp_lookup_1_FpMul_6U_10U_2_else_2_acc_1_nl;
  wire[7:0] inp_lookup_1_FpMul_6U_10U_2_oelse_1_acc_nl;
  wire[8:0] nl_inp_lookup_1_FpMul_6U_10U_2_oelse_1_acc_nl;
  wire[6:0] FpMul_6U_10U_2_oelse_1_acc_nl;
  wire[7:0] nl_FpMul_6U_10U_2_oelse_1_acc_nl;
  wire[0:0] mux_76_nl;
  wire[6:0] inp_lookup_2_FpMul_6U_10U_2_else_2_if_acc_nl;
  wire[7:0] nl_inp_lookup_2_FpMul_6U_10U_2_else_2_if_acc_nl;
  wire[6:0] inp_lookup_2_FpMul_6U_10U_2_else_2_acc_1_nl;
  wire[7:0] nl_inp_lookup_2_FpMul_6U_10U_2_else_2_acc_1_nl;
  wire[7:0] inp_lookup_2_FpMul_6U_10U_2_oelse_1_acc_nl;
  wire[8:0] nl_inp_lookup_2_FpMul_6U_10U_2_oelse_1_acc_nl;
  wire[6:0] FpMul_6U_10U_2_oelse_1_acc_1_nl;
  wire[7:0] nl_FpMul_6U_10U_2_oelse_1_acc_1_nl;
  wire[0:0] mux_77_nl;
  wire[6:0] inp_lookup_3_FpMul_6U_10U_2_else_2_if_acc_nl;
  wire[7:0] nl_inp_lookup_3_FpMul_6U_10U_2_else_2_if_acc_nl;
  wire[6:0] inp_lookup_3_FpMul_6U_10U_2_else_2_acc_1_nl;
  wire[7:0] nl_inp_lookup_3_FpMul_6U_10U_2_else_2_acc_1_nl;
  wire[7:0] inp_lookup_3_FpMul_6U_10U_2_oelse_1_acc_nl;
  wire[8:0] nl_inp_lookup_3_FpMul_6U_10U_2_oelse_1_acc_nl;
  wire[6:0] FpMul_6U_10U_2_oelse_1_acc_2_nl;
  wire[7:0] nl_FpMul_6U_10U_2_oelse_1_acc_2_nl;
  wire[0:0] mux_69_nl;
  wire[6:0] inp_lookup_4_FpMul_6U_10U_2_else_2_if_acc_nl;
  wire[7:0] nl_inp_lookup_4_FpMul_6U_10U_2_else_2_if_acc_nl;
  wire[6:0] inp_lookup_4_FpMul_6U_10U_2_else_2_acc_1_nl;
  wire[7:0] nl_inp_lookup_4_FpMul_6U_10U_2_else_2_acc_1_nl;
  wire[7:0] inp_lookup_4_FpMul_6U_10U_2_oelse_1_acc_nl;
  wire[8:0] nl_inp_lookup_4_FpMul_6U_10U_2_oelse_1_acc_nl;
  wire[6:0] FpMul_6U_10U_2_oelse_1_acc_3_nl;
  wire[7:0] nl_FpMul_6U_10U_2_oelse_1_acc_3_nl;
  wire[7:0] inp_lookup_1_FpAdd_8U_23U_if_3_if_acc_1_nl;
  wire[8:0] nl_inp_lookup_1_FpAdd_8U_23U_if_3_if_acc_1_nl;
  wire[7:0] inp_lookup_1_FpAdd_8U_23U_if_4_if_acc_nl;
  wire[8:0] nl_inp_lookup_1_FpAdd_8U_23U_if_4_if_acc_nl;
  wire[0:0] FpAdd_8U_23U_and_nl;
  wire[0:0] FpAdd_8U_23U_and_6_nl;
  wire[0:0] FpAdd_8U_23U_and_28_nl;
  wire[6:0] inp_lookup_1_FpMul_6U_10U_1_else_2_if_acc_nl;
  wire[7:0] nl_inp_lookup_1_FpMul_6U_10U_1_else_2_if_acc_nl;
  wire[6:0] inp_lookup_1_FpMul_6U_10U_1_else_2_acc_1_nl;
  wire[7:0] nl_inp_lookup_1_FpMul_6U_10U_1_else_2_acc_1_nl;
  wire[5:0] inp_lookup_1_FpMul_6U_10U_2_else_2_else_if_if_acc_1_nl;
  wire[6:0] nl_inp_lookup_1_FpMul_6U_10U_2_else_2_else_if_if_acc_1_nl;
  wire[0:0] FpMul_6U_10U_2_FpMul_6U_10U_2_and_20_nl;
  wire[7:0] inp_lookup_2_FpAdd_8U_23U_if_3_if_acc_1_nl;
  wire[8:0] nl_inp_lookup_2_FpAdd_8U_23U_if_3_if_acc_1_nl;
  wire[7:0] inp_lookup_2_FpAdd_8U_23U_if_4_if_acc_nl;
  wire[8:0] nl_inp_lookup_2_FpAdd_8U_23U_if_4_if_acc_nl;
  wire[0:0] FpAdd_8U_23U_and_29_nl;
  wire[0:0] FpAdd_8U_23U_and_13_nl;
  wire[0:0] FpAdd_8U_23U_and_30_nl;
  wire[6:0] inp_lookup_2_FpMul_6U_10U_1_else_2_if_acc_nl;
  wire[7:0] nl_inp_lookup_2_FpMul_6U_10U_1_else_2_if_acc_nl;
  wire[6:0] inp_lookup_2_FpMul_6U_10U_1_else_2_acc_1_nl;
  wire[7:0] nl_inp_lookup_2_FpMul_6U_10U_1_else_2_acc_1_nl;
  wire[5:0] inp_lookup_2_FpMul_6U_10U_2_else_2_else_if_if_acc_1_nl;
  wire[6:0] nl_inp_lookup_2_FpMul_6U_10U_2_else_2_else_if_if_acc_1_nl;
  wire[0:0] FpMul_6U_10U_2_FpMul_6U_10U_2_and_22_nl;
  wire[7:0] inp_lookup_3_FpAdd_8U_23U_if_3_if_acc_1_nl;
  wire[8:0] nl_inp_lookup_3_FpAdd_8U_23U_if_3_if_acc_1_nl;
  wire[7:0] inp_lookup_3_FpAdd_8U_23U_if_4_if_acc_nl;
  wire[8:0] nl_inp_lookup_3_FpAdd_8U_23U_if_4_if_acc_nl;
  wire[0:0] FpAdd_8U_23U_and_31_nl;
  wire[0:0] FpAdd_8U_23U_and_19_nl;
  wire[0:0] FpAdd_8U_23U_and_32_nl;
  wire[9:0] FpMul_6U_10U_2_FpMul_6U_10U_2_FpMul_6U_10U_2_nor_6_nl;
  wire[9:0] FpMul_6U_10U_2_nor_5_nl;
  wire[9:0] mux_2023_nl;
  wire[9:0] inp_lookup_3_FpMantRNE_22U_11U_2_else_acc_nl;
  wire[10:0] nl_inp_lookup_3_FpMantRNE_22U_11U_2_else_acc_nl;
  wire[0:0] or_5848_nl;
  wire[6:0] inp_lookup_3_FpMul_6U_10U_1_else_2_if_acc_nl;
  wire[7:0] nl_inp_lookup_3_FpMul_6U_10U_1_else_2_if_acc_nl;
  wire[6:0] inp_lookup_3_FpMul_6U_10U_1_else_2_acc_1_nl;
  wire[7:0] nl_inp_lookup_3_FpMul_6U_10U_1_else_2_acc_1_nl;
  wire[5:0] inp_lookup_3_FpMul_6U_10U_2_else_2_else_if_if_acc_1_nl;
  wire[6:0] nl_inp_lookup_3_FpMul_6U_10U_2_else_2_else_if_if_acc_1_nl;
  wire[0:0] FpMul_6U_10U_2_FpMul_6U_10U_2_and_24_nl;
  wire[7:0] inp_lookup_4_FpAdd_8U_23U_if_3_if_acc_1_nl;
  wire[8:0] nl_inp_lookup_4_FpAdd_8U_23U_if_3_if_acc_1_nl;
  wire[7:0] inp_lookup_4_FpAdd_8U_23U_if_4_if_acc_nl;
  wire[8:0] nl_inp_lookup_4_FpAdd_8U_23U_if_4_if_acc_nl;
  wire[0:0] FpAdd_8U_23U_and_33_nl;
  wire[0:0] FpAdd_8U_23U_and_25_nl;
  wire[0:0] FpAdd_8U_23U_and_34_nl;
  wire[6:0] inp_lookup_4_FpMul_6U_10U_1_else_2_if_acc_nl;
  wire[7:0] nl_inp_lookup_4_FpMul_6U_10U_1_else_2_if_acc_nl;
  wire[6:0] inp_lookup_4_FpMul_6U_10U_1_else_2_acc_1_nl;
  wire[7:0] nl_inp_lookup_4_FpMul_6U_10U_1_else_2_acc_1_nl;
  wire[5:0] inp_lookup_4_FpMul_6U_10U_2_else_2_else_if_if_acc_1_nl;
  wire[6:0] nl_inp_lookup_4_FpMul_6U_10U_2_else_2_else_if_if_acc_1_nl;
  wire[5:0] FpMul_6U_10U_1_else_2_else_acc_nl;
  wire[6:0] nl_FpMul_6U_10U_1_else_2_else_acc_nl;
  wire[5:0] inp_lookup_1_FpMul_6U_10U_1_else_2_else_if_if_acc_1_nl;
  wire[6:0] nl_inp_lookup_1_FpMul_6U_10U_1_else_2_else_if_if_acc_1_nl;
  wire[0:0] FpMul_6U_10U_1_FpMul_6U_10U_1_and_20_nl;
  wire[0:0] FpMul_6U_10U_2_FpMul_6U_10U_2_and_1_nl;
  wire[3:0] FpMul_6U_10U_2_FpMul_6U_10U_2_and_19_nl;
  wire[0:0] FpMul_6U_10U_2_oelse_2_not_27_nl;
  wire[0:0] FpMul_6U_10U_1_FpMul_6U_10U_1_and_1_nl;
  wire[3:0] FpMul_6U_10U_1_FpMul_6U_10U_1_and_19_nl;
  wire[0:0] FpMul_6U_10U_1_oelse_2_not_27_nl;
  wire[5:0] FpMul_6U_10U_1_else_2_else_acc_2_nl;
  wire[6:0] nl_FpMul_6U_10U_1_else_2_else_acc_2_nl;
  wire[5:0] inp_lookup_2_FpMul_6U_10U_1_else_2_else_if_if_acc_1_nl;
  wire[6:0] nl_inp_lookup_2_FpMul_6U_10U_1_else_2_else_if_if_acc_1_nl;
  wire[0:0] FpMul_6U_10U_1_FpMul_6U_10U_1_and_22_nl;
  wire[0:0] FpMul_6U_10U_2_FpMul_6U_10U_2_and_5_nl;
  wire[3:0] FpMul_6U_10U_2_FpMul_6U_10U_2_and_21_nl;
  wire[0:0] FpMul_6U_10U_2_oelse_2_not_26_nl;
  wire[0:0] FpMul_6U_10U_1_FpMul_6U_10U_1_and_5_nl;
  wire[3:0] FpMul_6U_10U_1_FpMul_6U_10U_1_and_21_nl;
  wire[0:0] FpMul_6U_10U_1_oelse_2_not_26_nl;
  wire[5:0] FpMul_6U_10U_1_else_2_else_acc_3_nl;
  wire[6:0] nl_FpMul_6U_10U_1_else_2_else_acc_3_nl;
  wire[5:0] inp_lookup_3_FpMul_6U_10U_1_else_2_else_if_if_acc_1_nl;
  wire[6:0] nl_inp_lookup_3_FpMul_6U_10U_1_else_2_else_if_if_acc_1_nl;
  wire[0:0] FpMul_6U_10U_1_FpMul_6U_10U_1_and_24_nl;
  wire[0:0] FpMul_6U_10U_2_FpMul_6U_10U_2_and_9_nl;
  wire[3:0] FpMul_6U_10U_2_FpMul_6U_10U_2_and_23_nl;
  wire[0:0] FpMul_6U_10U_2_oelse_2_not_25_nl;
  wire[9:0] FpMul_6U_10U_1_FpMul_6U_10U_1_FpMul_6U_10U_1_nor_6_nl;
  wire[9:0] FpMul_6U_10U_1_nor_5_nl;
  wire[9:0] mux_2024_nl;
  wire[9:0] inp_lookup_3_FpMantRNE_22U_11U_1_else_acc_nl;
  wire[10:0] nl_inp_lookup_3_FpMantRNE_22U_11U_1_else_acc_nl;
  wire[0:0] or_5849_nl;
  wire[0:0] FpMul_6U_10U_1_or_9_nl;
  wire[0:0] FpMul_6U_10U_1_FpMul_6U_10U_1_and_9_nl;
  wire[3:0] FpMul_6U_10U_1_FpMul_6U_10U_1_and_23_nl;
  wire[0:0] FpMul_6U_10U_1_oelse_2_not_25_nl;
  wire[5:0] FpMul_6U_10U_1_else_2_else_acc_4_nl;
  wire[6:0] nl_FpMul_6U_10U_1_else_2_else_acc_4_nl;
  wire[5:0] inp_lookup_4_FpMul_6U_10U_1_else_2_else_if_if_acc_1_nl;
  wire[6:0] nl_inp_lookup_4_FpMul_6U_10U_1_else_2_else_if_if_acc_1_nl;
  wire[0:0] FpMul_6U_10U_1_FpMul_6U_10U_1_and_26_nl;
  wire[0:0] FpMul_6U_10U_2_FpMul_6U_10U_2_and_26_nl;
  wire[0:0] FpMul_6U_10U_2_FpMul_6U_10U_2_and_13_nl;
  wire[3:0] FpMul_6U_10U_2_FpMul_6U_10U_2_and_25_nl;
  wire[0:0] FpMul_6U_10U_2_oelse_2_not_24_nl;
  wire[0:0] FpMul_6U_10U_1_FpMul_6U_10U_1_and_13_nl;
  wire[3:0] FpMul_6U_10U_1_FpMul_6U_10U_1_and_25_nl;
  wire[0:0] FpMul_6U_10U_1_oelse_2_not_24_nl;
  wire[7:0] FpNormalize_8U_49U_1_FpNormalize_8U_49U_1_and_nl;
  wire[7:0] inp_lookup_1_FpNormalize_8U_49U_1_else_acc_nl;
  wire[9:0] nl_inp_lookup_1_FpNormalize_8U_49U_1_else_acc_nl;
  wire[7:0] inp_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_nl;
  wire[8:0] nl_inp_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_nl;
  wire[0:0] FpAdd_8U_23U_1_and_4_nl;
  wire[0:0] FpAdd_8U_23U_1_and_5_nl;
  wire[7:0] FpNormalize_8U_49U_1_FpNormalize_8U_49U_1_and_2_nl;
  wire[7:0] inp_lookup_2_FpNormalize_8U_49U_1_else_acc_nl;
  wire[9:0] nl_inp_lookup_2_FpNormalize_8U_49U_1_else_acc_nl;
  wire[7:0] inp_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_nl;
  wire[8:0] nl_inp_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_nl;
  wire[0:0] FpAdd_8U_23U_1_and_10_nl;
  wire[0:0] FpAdd_8U_23U_1_and_11_nl;
  wire[7:0] FpNormalize_8U_49U_1_FpNormalize_8U_49U_1_and_4_nl;
  wire[7:0] inp_lookup_3_FpNormalize_8U_49U_1_else_acc_nl;
  wire[9:0] nl_inp_lookup_3_FpNormalize_8U_49U_1_else_acc_nl;
  wire[7:0] inp_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_nl;
  wire[8:0] nl_inp_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_nl;
  wire[0:0] FpAdd_8U_23U_1_and_16_nl;
  wire[0:0] FpAdd_8U_23U_1_and_17_nl;
  wire[7:0] FpNormalize_8U_49U_1_FpNormalize_8U_49U_1_and_6_nl;
  wire[7:0] inp_lookup_4_FpNormalize_8U_49U_1_else_acc_nl;
  wire[9:0] nl_inp_lookup_4_FpNormalize_8U_49U_1_else_acc_nl;
  wire[7:0] inp_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_nl;
  wire[8:0] nl_inp_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_nl;
  wire[0:0] FpAdd_8U_23U_1_and_22_nl;
  wire[0:0] FpAdd_8U_23U_1_and_23_nl;
  wire[8:0] inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_nl;
  wire[9:0] nl_inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_nl;
  wire[22:0] inp_lookup_1_FpMantRNE_49U_24U_1_else_acc_nl;
  wire[23:0] nl_inp_lookup_1_FpMantRNE_49U_24U_1_else_acc_nl;
  wire[7:0] inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_nl;
  wire[8:0] nl_inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_nl;
  wire[8:0] inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_nl;
  wire[9:0] nl_inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_nl;
  wire[22:0] inp_lookup_2_FpMantRNE_49U_24U_1_else_acc_nl;
  wire[23:0] nl_inp_lookup_2_FpMantRNE_49U_24U_1_else_acc_nl;
  wire[8:0] inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_nl;
  wire[9:0] nl_inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_nl;
  wire[7:0] inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_nl;
  wire[8:0] nl_inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_nl;
  wire[8:0] inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_nl;
  wire[9:0] nl_inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_nl;
  wire[22:0] FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_6_nl;
  wire[22:0] inp_lookup_3_FpMantRNE_49U_24U_1_else_acc_nl;
  wire[23:0] nl_inp_lookup_3_FpMantRNE_49U_24U_1_else_acc_nl;
  wire[8:0] inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_nl;
  wire[9:0] nl_inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_nl;
  wire[7:0] inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_nl;
  wire[8:0] nl_inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_nl;
  wire[8:0] inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_nl;
  wire[9:0] nl_inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_nl;
  wire[22:0] inp_lookup_4_FpMantRNE_49U_24U_1_else_acc_nl;
  wire[23:0] nl_inp_lookup_4_FpMantRNE_49U_24U_1_else_acc_nl;
  wire[8:0] inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_nl;
  wire[9:0] nl_inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_nl;
  wire[7:0] inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_nl;
  wire[8:0] nl_inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_nl;
  wire[8:0] inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_nl;
  wire[9:0] nl_inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_nl;
  wire[0:0] FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_else_mux_8_nl;
  wire[4:0] FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_and_nl;
  wire[4:0] FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_mux1h_nl;
  wire[0:0] FpWidthDec_8U_23U_6U_10U_0U_1U_and_11_nl;
  wire[0:0] FpWidthDec_8U_23U_6U_10U_0U_1U_and_12_nl;
  wire[0:0] FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_not_8_nl;
  wire[0:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_14_nl;
  wire[0:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_2_nl;
  wire[9:0] inp_lookup_1_FpMantRNE_23U_11U_1_else_acc_nl;
  wire[10:0] nl_inp_lookup_1_FpMantRNE_23U_11U_1_else_acc_nl;
  wire[0:0] FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_else_mux_9_nl;
  wire[4:0] FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_and_2_nl;
  wire[4:0] FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_mux1h_1_nl;
  wire[0:0] FpWidthDec_8U_23U_6U_10U_0U_1U_and_13_nl;
  wire[0:0] FpWidthDec_8U_23U_6U_10U_0U_1U_and_14_nl;
  wire[0:0] FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_not_9_nl;
  wire[0:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_17_nl;
  wire[0:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_5_nl;
  wire[9:0] inp_lookup_2_FpMantRNE_23U_11U_1_else_acc_nl;
  wire[10:0] nl_inp_lookup_2_FpMantRNE_23U_11U_1_else_acc_nl;
  wire[0:0] FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_else_mux_10_nl;
  wire[4:0] FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_and_4_nl;
  wire[4:0] FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_mux1h_2_nl;
  wire[0:0] FpWidthDec_8U_23U_6U_10U_0U_1U_and_15_nl;
  wire[0:0] FpWidthDec_8U_23U_6U_10U_0U_1U_and_16_nl;
  wire[0:0] FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_not_10_nl;
  wire[0:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_20_nl;
  wire[0:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_8_nl;
  wire[9:0] inp_lookup_3_FpMantRNE_23U_11U_1_else_acc_nl;
  wire[10:0] nl_inp_lookup_3_FpMantRNE_23U_11U_1_else_acc_nl;
  wire[0:0] FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_else_mux_11_nl;
  wire[4:0] FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_and_6_nl;
  wire[4:0] FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_mux1h_3_nl;
  wire[0:0] FpWidthDec_8U_23U_6U_10U_0U_1U_and_17_nl;
  wire[0:0] FpWidthDec_8U_23U_6U_10U_0U_1U_and_18_nl;
  wire[0:0] FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_not_11_nl;
  wire[0:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_23_nl;
  wire[0:0] FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_11_nl;
  wire[9:0] inp_lookup_4_FpMantRNE_23U_11U_1_else_acc_nl;
  wire[10:0] nl_inp_lookup_4_FpMantRNE_23U_11U_1_else_acc_nl;
  wire[6:0] inp_lookup_1_FpMul_6U_10U_else_2_if_acc_nl;
  wire[7:0] nl_inp_lookup_1_FpMul_6U_10U_else_2_if_acc_nl;
  wire[6:0] inp_lookup_1_FpMul_6U_10U_else_2_acc_1_nl;
  wire[7:0] nl_inp_lookup_1_FpMul_6U_10U_else_2_acc_1_nl;
  wire[6:0] inp_lookup_2_FpMul_6U_10U_else_2_if_acc_nl;
  wire[7:0] nl_inp_lookup_2_FpMul_6U_10U_else_2_if_acc_nl;
  wire[6:0] inp_lookup_2_FpMul_6U_10U_else_2_acc_1_nl;
  wire[7:0] nl_inp_lookup_2_FpMul_6U_10U_else_2_acc_1_nl;
  wire[6:0] inp_lookup_3_FpMul_6U_10U_else_2_if_acc_nl;
  wire[7:0] nl_inp_lookup_3_FpMul_6U_10U_else_2_if_acc_nl;
  wire[6:0] inp_lookup_3_FpMul_6U_10U_else_2_acc_1_nl;
  wire[7:0] nl_inp_lookup_3_FpMul_6U_10U_else_2_acc_1_nl;
  wire[6:0] inp_lookup_4_FpMul_6U_10U_else_2_if_acc_nl;
  wire[7:0] nl_inp_lookup_4_FpMul_6U_10U_else_2_if_acc_nl;
  wire[6:0] inp_lookup_4_FpMul_6U_10U_else_2_acc_1_nl;
  wire[7:0] nl_inp_lookup_4_FpMul_6U_10U_else_2_acc_1_nl;
  wire[9:0] FpMul_6U_10U_FpMul_6U_10U_FpMul_6U_10U_nor_4_nl;
  wire[9:0] FpMul_6U_10U_nor_nl;
  wire[9:0] mux_2025_nl;
  wire[9:0] inp_lookup_1_FpMantRNE_22U_11U_else_acc_nl;
  wire[10:0] nl_inp_lookup_1_FpMantRNE_22U_11U_else_acc_nl;
  wire[0:0] or_5850_nl;
  wire[0:0] FpMul_6U_10U_or_8_nl;
  wire[3:0] FpMul_6U_10U_FpMul_6U_10U_and_15_nl;
  wire[0:0] FpMul_6U_10U_oelse_2_not_27_nl;
  wire[6:0] FpAdd_6U_10U_is_a_greater_acc_nl;
  wire[8:0] nl_FpAdd_6U_10U_is_a_greater_acc_nl;
  wire[9:0] FpMul_6U_10U_FpMul_6U_10U_FpMul_6U_10U_nor_5_nl;
  wire[9:0] FpMul_6U_10U_nor_4_nl;
  wire[9:0] mux_2026_nl;
  wire[9:0] inp_lookup_2_FpMantRNE_22U_11U_else_acc_nl;
  wire[10:0] nl_inp_lookup_2_FpMantRNE_22U_11U_else_acc_nl;
  wire[0:0] or_5851_nl;
  wire[0:0] FpMul_6U_10U_or_9_nl;
  wire[3:0] FpMul_6U_10U_FpMul_6U_10U_and_17_nl;
  wire[0:0] FpMul_6U_10U_oelse_2_not_26_nl;
  wire[6:0] FpAdd_6U_10U_is_a_greater_acc_1_nl;
  wire[8:0] nl_FpAdd_6U_10U_is_a_greater_acc_1_nl;
  wire[9:0] FpMul_6U_10U_FpMul_6U_10U_FpMul_6U_10U_nor_6_nl;
  wire[9:0] FpMul_6U_10U_nor_5_nl;
  wire[9:0] mux_2027_nl;
  wire[9:0] inp_lookup_3_FpMantRNE_22U_11U_else_acc_nl;
  wire[10:0] nl_inp_lookup_3_FpMantRNE_22U_11U_else_acc_nl;
  wire[0:0] or_5852_nl;
  wire[0:0] FpMul_6U_10U_or_10_nl;
  wire[3:0] FpMul_6U_10U_FpMul_6U_10U_and_19_nl;
  wire[0:0] FpMul_6U_10U_oelse_2_not_25_nl;
  wire[6:0] FpAdd_6U_10U_is_a_greater_acc_2_nl;
  wire[8:0] nl_FpAdd_6U_10U_is_a_greater_acc_2_nl;
  wire[9:0] FpMul_6U_10U_FpMul_6U_10U_FpMul_6U_10U_nor_7_nl;
  wire[9:0] FpMul_6U_10U_nor_6_nl;
  wire[9:0] mux_2028_nl;
  wire[9:0] inp_lookup_4_FpMantRNE_22U_11U_else_acc_nl;
  wire[10:0] nl_inp_lookup_4_FpMantRNE_22U_11U_else_acc_nl;
  wire[0:0] or_5853_nl;
  wire[0:0] FpMul_6U_10U_or_11_nl;
  wire[3:0] FpMul_6U_10U_FpMul_6U_10U_and_21_nl;
  wire[0:0] FpMul_6U_10U_oelse_2_not_24_nl;
  wire[6:0] FpAdd_6U_10U_is_a_greater_acc_3_nl;
  wire[8:0] nl_FpAdd_6U_10U_is_a_greater_acc_3_nl;
  wire[1:0] FpAdd_6U_10U_FpAdd_6U_10U_mux1h_13_nl;
  wire[5:0] inp_lookup_1_FpAdd_6U_10U_if_3_if_acc_1_nl;
  wire[6:0] nl_inp_lookup_1_FpAdd_6U_10U_if_3_if_acc_1_nl;
  wire[6:0] inp_lookup_1_FpNormalize_6U_23U_acc_nl;
  wire[8:0] nl_inp_lookup_1_FpNormalize_6U_23U_acc_nl;
  wire[1:0] FpAdd_6U_10U_FpAdd_6U_10U_mux1h_15_nl;
  wire[5:0] inp_lookup_2_FpAdd_6U_10U_if_3_if_acc_1_nl;
  wire[6:0] nl_inp_lookup_2_FpAdd_6U_10U_if_3_if_acc_1_nl;
  wire[6:0] inp_lookup_2_FpNormalize_6U_23U_acc_nl;
  wire[8:0] nl_inp_lookup_2_FpNormalize_6U_23U_acc_nl;
  wire[1:0] FpAdd_6U_10U_FpAdd_6U_10U_mux1h_17_nl;
  wire[5:0] inp_lookup_3_FpAdd_6U_10U_if_3_if_acc_1_nl;
  wire[6:0] nl_inp_lookup_3_FpAdd_6U_10U_if_3_if_acc_1_nl;
  wire[6:0] inp_lookup_3_FpNormalize_6U_23U_acc_nl;
  wire[8:0] nl_inp_lookup_3_FpNormalize_6U_23U_acc_nl;
  wire[1:0] FpAdd_6U_10U_FpAdd_6U_10U_mux1h_19_nl;
  wire[5:0] inp_lookup_4_FpAdd_6U_10U_if_3_if_acc_1_nl;
  wire[6:0] nl_inp_lookup_4_FpAdd_6U_10U_if_3_if_acc_1_nl;
  wire[6:0] inp_lookup_4_FpNormalize_6U_23U_acc_nl;
  wire[8:0] nl_inp_lookup_4_FpNormalize_6U_23U_acc_nl;
  wire[7:0] inp_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_nl;
  wire[8:0] nl_inp_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_nl;
  wire[0:0] FpAdd_8U_23U_1_or_nl;
  wire[0:0] FpAdd_8U_23U_1_and_6_nl;
  wire[0:0] FpAdd_8U_23U_1_and_28_nl;
  wire[0:0] or_6234_nl;
  wire[0:0] or_6233_nl;
  wire[0:0] or_6232_nl;
  wire[9:0] FpMul_6U_10U_2_FpMul_6U_10U_2_FpMul_6U_10U_2_nor_4_nl;
  wire[9:0] FpMul_6U_10U_2_nor_nl;
  wire[9:0] mux_2029_nl;
  wire[9:0] inp_lookup_1_FpMantRNE_22U_11U_2_else_acc_nl;
  wire[10:0] nl_inp_lookup_1_FpMantRNE_22U_11U_2_else_acc_nl;
  wire[0:0] or_5854_nl;
  wire[9:0] FpMul_6U_10U_2_nor_4_nl;
  wire[9:0] mux_2030_nl;
  wire[9:0] inp_lookup_2_FpMantRNE_22U_11U_2_else_acc_nl;
  wire[10:0] nl_inp_lookup_2_FpMantRNE_22U_11U_2_else_acc_nl;
  wire[0:0] or_5855_nl;
  wire[9:0] FpMul_6U_10U_2_FpMul_6U_10U_2_FpMul_6U_10U_2_nor_7_nl;
  wire[9:0] FpMul_6U_10U_2_nor_6_nl;
  wire[9:0] mux_2031_nl;
  wire[9:0] inp_lookup_4_FpMantRNE_22U_11U_2_else_acc_nl;
  wire[10:0] nl_inp_lookup_4_FpMantRNE_22U_11U_2_else_acc_nl;
  wire[0:0] or_5856_nl;
  wire[0:0] inp_lookup_else_if_not_nl;
  wire[0:0] inp_lookup_else_if_not_1_nl;
  wire[0:0] inp_lookup_else_if_not_2_nl;
  wire[0:0] inp_lookup_else_if_not_3_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_mux_4_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_and_nl;
  wire[0:0] IsZero_5U_10U_3_aelse_not_23_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_mux_36_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_and_3_nl;
  wire[0:0] IsZero_5U_10U_3_aelse_not_22_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_mux_37_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_and_6_nl;
  wire[0:0] IsZero_5U_10U_3_aelse_not_21_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_mux_38_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_and_9_nl;
  wire[0:0] IsZero_5U_10U_3_aelse_not_20_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_18_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_4_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux1h_4_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_16_nl;
  wire[0:0] IsZero_5U_10U_1_aelse_not_27_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_20_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_6_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux1h_6_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_18_nl;
  wire[0:0] IsZero_5U_10U_1_aelse_not_26_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_22_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_8_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux1h_8_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_20_nl;
  wire[0:0] IsZero_5U_10U_1_aelse_not_25_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_24_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_10_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux1h_10_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_22_nl;
  wire[0:0] IsZero_5U_10U_1_aelse_not_24_nl;
  wire[4:0] inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_else_else_else_acc_nl;
  wire[5:0] nl_inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_else_else_else_acc_nl;
  wire[0:0] FpFractionToFloat_35U_6U_10U_1_and_nl;
  wire[4:0] FpFractionToFloat_35U_6U_10U_1_nor_4_nl;
  wire[4:0] inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_else_else_else_acc_nl;
  wire[5:0] nl_inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_else_else_else_acc_nl;
  wire[4:0] FpFractionToFloat_35U_6U_10U_1_nor_nl;
  wire[4:0] inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_else_else_else_acc_nl;
  wire[5:0] nl_inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_else_else_else_acc_nl;
  wire[4:0] FpFractionToFloat_35U_6U_10U_1_nor_5_nl;
  wire[4:0] inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_else_else_else_acc_nl;
  wire[5:0] nl_inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_else_else_else_acc_nl;
  wire[0:0] FpFractionToFloat_35U_6U_10U_1_and_3_nl;
  wire[4:0] FpFractionToFloat_35U_6U_10U_1_nor_6_nl;
  wire[8:0] inp_lookup_1_FpNormalize_8U_49U_acc_nl;
  wire[10:0] nl_inp_lookup_1_FpNormalize_8U_49U_acc_nl;
  wire[8:0] inp_lookup_2_FpNormalize_8U_49U_acc_nl;
  wire[10:0] nl_inp_lookup_2_FpNormalize_8U_49U_acc_nl;
  wire[8:0] inp_lookup_3_FpNormalize_8U_49U_acc_nl;
  wire[10:0] nl_inp_lookup_3_FpNormalize_8U_49U_acc_nl;
  wire[8:0] inp_lookup_4_FpNormalize_8U_49U_acc_nl;
  wire[10:0] nl_inp_lookup_4_FpNormalize_8U_49U_acc_nl;
  wire[5:0] FpMul_6U_10U_2_else_2_else_acc_nl;
  wire[6:0] nl_FpMul_6U_10U_2_else_2_else_acc_nl;
  wire[5:0] FpMul_6U_10U_2_else_2_else_acc_2_nl;
  wire[6:0] nl_FpMul_6U_10U_2_else_2_else_acc_2_nl;
  wire[5:0] FpMul_6U_10U_2_else_2_else_acc_3_nl;
  wire[6:0] nl_FpMul_6U_10U_2_else_2_else_acc_3_nl;
  wire[5:0] FpMul_6U_10U_2_else_2_else_acc_4_nl;
  wire[6:0] nl_FpMul_6U_10U_2_else_2_else_acc_4_nl;
  wire[22:0] inp_lookup_1_FpMantRNE_49U_24U_else_acc_nl;
  wire[23:0] nl_inp_lookup_1_FpMantRNE_49U_24U_else_acc_nl;
  wire[22:0] inp_lookup_2_FpMantRNE_49U_24U_else_acc_nl;
  wire[23:0] nl_inp_lookup_2_FpMantRNE_49U_24U_else_acc_nl;
  wire[22:0] inp_lookup_3_FpMantRNE_49U_24U_else_acc_nl;
  wire[23:0] nl_inp_lookup_3_FpMantRNE_49U_24U_else_acc_nl;
  wire[22:0] inp_lookup_4_FpMantRNE_49U_24U_else_acc_nl;
  wire[23:0] nl_inp_lookup_4_FpMantRNE_49U_24U_else_acc_nl;
  wire[6:0] FpAdd_6U_10U_1_is_a_greater_acc_3_nl;
  wire[8:0] nl_FpAdd_6U_10U_1_is_a_greater_acc_3_nl;
  wire[6:0] FpAdd_6U_10U_1_is_a_greater_acc_2_nl;
  wire[8:0] nl_FpAdd_6U_10U_1_is_a_greater_acc_2_nl;
  wire[6:0] FpAdd_6U_10U_1_is_a_greater_acc_1_nl;
  wire[8:0] nl_FpAdd_6U_10U_1_is_a_greater_acc_1_nl;
  wire[6:0] FpAdd_6U_10U_1_is_a_greater_acc_nl;
  wire[8:0] nl_FpAdd_6U_10U_1_is_a_greater_acc_nl;
  wire[9:0] FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_nl;
  wire[9:0] FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_mux_1_nl;
  wire[9:0] inp_lookup_1_FpMantRNE_24U_11U_else_acc_nl;
  wire[10:0] nl_inp_lookup_1_FpMantRNE_24U_11U_else_acc_nl;
  wire[9:0] FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_1_nl;
  wire[9:0] FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_mux_14_nl;
  wire[9:0] inp_lookup_2_FpMantRNE_24U_11U_else_acc_nl;
  wire[10:0] nl_inp_lookup_2_FpMantRNE_24U_11U_else_acc_nl;
  wire[9:0] FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_2_nl;
  wire[9:0] FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_mux_27_nl;
  wire[9:0] inp_lookup_3_FpMantRNE_24U_11U_else_acc_nl;
  wire[10:0] nl_inp_lookup_3_FpMantRNE_24U_11U_else_acc_nl;
  wire[9:0] FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_3_nl;
  wire[9:0] FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_mux_40_nl;
  wire[9:0] inp_lookup_4_FpMantRNE_24U_11U_else_acc_nl;
  wire[10:0] nl_inp_lookup_4_FpMantRNE_24U_11U_else_acc_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux_47_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_26_nl;
  wire[0:0] IsZero_5U_10U_1_aelse_not_21_nl;
  wire[7:0] inp_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_1_nl;
  wire[8:0] nl_inp_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_1_nl;
  wire[7:0] inp_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_1_nl;
  wire[8:0] nl_inp_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_1_nl;
  wire[7:0] inp_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_1_nl;
  wire[8:0] nl_inp_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_1_nl;
  wire[7:0] inp_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_1_nl;
  wire[8:0] nl_inp_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_1_nl;
  wire[0:0] FpMul_6U_10U_FpMul_6U_10U_and_16_nl;
  wire[0:0] FpMul_6U_10U_FpMul_6U_10U_and_1_nl;
  wire[0:0] FpMul_6U_10U_FpMul_6U_10U_and_18_nl;
  wire[0:0] FpMul_6U_10U_FpMul_6U_10U_and_4_nl;
  wire[0:0] FpMul_6U_10U_FpMul_6U_10U_and_20_nl;
  wire[0:0] FpMul_6U_10U_FpMul_6U_10U_and_7_nl;
  wire[0:0] FpMul_6U_10U_FpMul_6U_10U_and_22_nl;
  wire[0:0] FpMul_6U_10U_FpMul_6U_10U_and_10_nl;
  wire[0:0] IsNaN_6U_23U_2_aelse_not_11_nl;
  wire[0:0] IsNaN_6U_23U_2_aelse_not_10_nl;
  wire[0:0] IsNaN_6U_23U_2_aelse_not_9_nl;
  wire[0:0] IsNaN_6U_23U_2_aelse_not_8_nl;
  wire[9:0] FpMul_6U_10U_1_nor_nl;
  wire[9:0] mux_2032_nl;
  wire[9:0] inp_lookup_1_FpMantRNE_22U_11U_1_else_acc_nl;
  wire[10:0] nl_inp_lookup_1_FpMantRNE_22U_11U_1_else_acc_nl;
  wire[0:0] or_5857_nl;
  wire[9:0] FpMul_6U_10U_1_nor_4_nl;
  wire[9:0] mux_2033_nl;
  wire[9:0] inp_lookup_2_FpMantRNE_22U_11U_1_else_acc_nl;
  wire[10:0] nl_inp_lookup_2_FpMantRNE_22U_11U_1_else_acc_nl;
  wire[0:0] or_5858_nl;
  wire[9:0] FpMul_6U_10U_1_nor_6_nl;
  wire[9:0] mux_2034_nl;
  wire[9:0] inp_lookup_4_FpMantRNE_22U_11U_1_else_acc_nl;
  wire[10:0] nl_inp_lookup_4_FpMantRNE_22U_11U_1_else_acc_nl;
  wire[0:0] or_5859_nl;
  wire[0:0] or_6166_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_mux_2_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_mux1h_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_2_nl;
  wire[0:0] IsZero_5U_10U_aelse_not_27_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_mux_7_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_1_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_mux1h_1_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_5_nl;
  wire[0:0] IsZero_5U_10U_aelse_not_26_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_mux_12_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_2_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_mux1h_2_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_8_nl;
  wire[0:0] IsZero_5U_10U_aelse_not_25_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_mux_17_nl;
  wire[0:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_3_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_mux1h_3_nl;
  wire[3:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_11_nl;
  wire[0:0] IsZero_5U_10U_aelse_not_24_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_mux_4_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_nl;
  wire[0:0] IsZero_5U_10U_aelse_not_23_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_mux_36_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_3_nl;
  wire[0:0] IsZero_5U_10U_aelse_not_22_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_mux_37_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_6_nl;
  wire[0:0] IsZero_5U_10U_aelse_not_21_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_mux_38_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_9_nl;
  wire[0:0] IsZero_5U_10U_aelse_not_20_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux_43_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_18_nl;
  wire[0:0] IsZero_5U_10U_1_aelse_not_23_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux_45_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_22_nl;
  wire[0:0] IsZero_5U_10U_1_aelse_not_22_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux_49_nl;
  wire[9:0] FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_30_nl;
  wire[0:0] IsZero_5U_10U_1_aelse_not_20_nl;
  wire[0:0] FpAdd_8U_23U_mux_1_nl;
  wire[0:0] FpAdd_8U_23U_mux_17_nl;
  wire[0:0] FpAdd_8U_23U_mux_33_nl;
  wire[0:0] FpAdd_8U_23U_mux_49_nl;
  wire[5:0] inp_lookup_1_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_nl;
  wire[6:0] nl_inp_lookup_1_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_nl;
  wire[5:0] inp_lookup_2_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_nl;
  wire[6:0] nl_inp_lookup_2_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_nl;
  wire[5:0] inp_lookup_3_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_nl;
  wire[6:0] nl_inp_lookup_3_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_nl;
  wire[5:0] inp_lookup_4_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_nl;
  wire[6:0] nl_inp_lookup_4_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_nl;
  wire[7:0] inp_lookup_1_FpMul_6U_10U_1_oelse_1_acc_nl;
  wire[8:0] nl_inp_lookup_1_FpMul_6U_10U_1_oelse_1_acc_nl;
  wire[6:0] FpMul_6U_10U_1_oelse_1_acc_nl;
  wire[7:0] nl_FpMul_6U_10U_1_oelse_1_acc_nl;
  wire[7:0] inp_lookup_2_FpMul_6U_10U_1_oelse_1_acc_nl;
  wire[8:0] nl_inp_lookup_2_FpMul_6U_10U_1_oelse_1_acc_nl;
  wire[6:0] FpMul_6U_10U_1_oelse_1_acc_1_nl;
  wire[7:0] nl_FpMul_6U_10U_1_oelse_1_acc_1_nl;
  wire[7:0] inp_lookup_3_FpMul_6U_10U_1_oelse_1_acc_nl;
  wire[8:0] nl_inp_lookup_3_FpMul_6U_10U_1_oelse_1_acc_nl;
  wire[6:0] FpMul_6U_10U_1_oelse_1_acc_2_nl;
  wire[7:0] nl_FpMul_6U_10U_1_oelse_1_acc_2_nl;
  wire[7:0] inp_lookup_4_FpMul_6U_10U_1_oelse_1_acc_nl;
  wire[8:0] nl_inp_lookup_4_FpMul_6U_10U_1_oelse_1_acc_nl;
  wire[6:0] FpMul_6U_10U_1_oelse_1_acc_3_nl;
  wire[7:0] nl_FpMul_6U_10U_1_oelse_1_acc_3_nl;
  wire[0:0] FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_nl;
  wire[7:0] inp_lookup_1_FpAdd_8U_23U_if_4_if_acc_1_nl;
  wire[8:0] nl_inp_lookup_1_FpAdd_8U_23U_if_4_if_acc_1_nl;
  wire[8:0] FpAdd_8U_23U_1_is_a_greater_acc_nl;
  wire[10:0] nl_FpAdd_8U_23U_1_is_a_greater_acc_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_1_nl;
  wire[0:0] FpNormalize_8U_49U_oelse_not_nl;
  wire[2:0] inp_lookup_1_IntSaturation_51U_32U_if_acc_nl;
  wire[3:0] nl_inp_lookup_1_IntSaturation_51U_32U_if_acc_nl;
  wire[0:0] FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_1_nl;
  wire[7:0] inp_lookup_2_FpAdd_8U_23U_if_4_if_acc_1_nl;
  wire[8:0] nl_inp_lookup_2_FpAdd_8U_23U_if_4_if_acc_1_nl;
  wire[8:0] FpAdd_8U_23U_1_is_a_greater_acc_1_nl;
  wire[10:0] nl_FpAdd_8U_23U_1_is_a_greater_acc_1_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_3_nl;
  wire[0:0] FpNormalize_8U_49U_oelse_not_1_nl;
  wire[2:0] inp_lookup_2_IntSaturation_51U_32U_if_acc_nl;
  wire[3:0] nl_inp_lookup_2_IntSaturation_51U_32U_if_acc_nl;
  wire[0:0] FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_2_nl;
  wire[7:0] inp_lookup_3_FpAdd_8U_23U_if_4_if_acc_1_nl;
  wire[8:0] nl_inp_lookup_3_FpAdd_8U_23U_if_4_if_acc_1_nl;
  wire[8:0] FpAdd_8U_23U_1_is_a_greater_acc_2_nl;
  wire[10:0] nl_FpAdd_8U_23U_1_is_a_greater_acc_2_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_5_nl;
  wire[0:0] FpNormalize_8U_49U_oelse_not_2_nl;
  wire[2:0] inp_lookup_3_IntSaturation_51U_32U_if_acc_nl;
  wire[3:0] nl_inp_lookup_3_IntSaturation_51U_32U_if_acc_nl;
  wire[0:0] FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_3_nl;
  wire[7:0] inp_lookup_4_FpAdd_8U_23U_if_4_if_acc_1_nl;
  wire[8:0] nl_inp_lookup_4_FpAdd_8U_23U_if_4_if_acc_1_nl;
  wire[8:0] FpAdd_8U_23U_1_is_a_greater_acc_3_nl;
  wire[10:0] nl_FpAdd_8U_23U_1_is_a_greater_acc_3_nl;
  wire[48:0] FpNormalize_8U_49U_FpNormalize_8U_49U_and_7_nl;
  wire[0:0] FpNormalize_8U_49U_oelse_not_3_nl;
  wire[2:0] inp_lookup_4_IntSaturation_51U_32U_if_acc_nl;
  wire[3:0] nl_inp_lookup_4_IntSaturation_51U_32U_if_acc_nl;
  wire[5:0] inp_lookup_1_FpMul_6U_10U_1_else_2_else_if_if_acc_nl;
  wire[6:0] nl_inp_lookup_1_FpMul_6U_10U_1_else_2_else_if_if_acc_nl;
  wire[0:0] FpMul_6U_10U_1_or_4_nl;
  wire[0:0] FpMantWidthDec_6U_21U_10U_0U_0U_1_and_1_nl;
  wire[5:0] inp_lookup_2_FpMul_6U_10U_1_else_2_else_if_if_acc_nl;
  wire[6:0] nl_inp_lookup_2_FpMul_6U_10U_1_else_2_else_if_if_acc_nl;
  wire[0:0] FpMul_6U_10U_1_or_5_nl;
  wire[0:0] FpMantWidthDec_6U_21U_10U_0U_0U_1_and_3_nl;
  wire[5:0] inp_lookup_3_FpMul_6U_10U_1_else_2_else_if_if_acc_nl;
  wire[6:0] nl_inp_lookup_3_FpMul_6U_10U_1_else_2_else_if_if_acc_nl;
  wire[0:0] FpMul_6U_10U_1_or_6_nl;
  wire[0:0] FpMantWidthDec_6U_21U_10U_0U_0U_1_and_5_nl;
  wire[5:0] inp_lookup_4_FpMul_6U_10U_1_else_2_else_if_if_acc_nl;
  wire[6:0] nl_inp_lookup_4_FpMul_6U_10U_1_else_2_else_if_if_acc_nl;
  wire[0:0] FpMul_6U_10U_1_FpMul_6U_10U_1_nor_11_nl;
  wire[0:0] FpMul_6U_10U_1_or_7_nl;
  wire[0:0] FpMantWidthDec_6U_21U_10U_0U_0U_1_and_7_nl;
  wire[7:0] inp_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_1_nl;
  wire[8:0] nl_inp_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_1_nl;
  wire[48:0] FpNormalize_8U_49U_1_FpNormalize_8U_49U_1_and_1_nl;
  wire[10:0] FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_nl;
  wire[12:0] nl_FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_nl;
  wire[7:0] inp_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_1_nl;
  wire[8:0] nl_inp_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_1_nl;
  wire[48:0] FpNormalize_8U_49U_1_FpNormalize_8U_49U_1_and_3_nl;
  wire[10:0] FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_1_nl;
  wire[12:0] nl_FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_1_nl;
  wire[7:0] inp_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_1_nl;
  wire[8:0] nl_inp_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_1_nl;
  wire[48:0] FpNormalize_8U_49U_1_FpNormalize_8U_49U_1_and_5_nl;
  wire[10:0] FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_2_nl;
  wire[12:0] nl_FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_2_nl;
  wire[7:0] inp_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_1_nl;
  wire[8:0] nl_inp_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_1_nl;
  wire[48:0] FpNormalize_8U_49U_1_FpNormalize_8U_49U_1_and_7_nl;
  wire[10:0] FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_3_nl;
  wire[12:0] nl_FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_3_nl;
  wire[0:0] FpAdd_8U_23U_1_if_4_FpAdd_8U_23U_1_if_4_or_4_nl;
  wire[7:0] inp_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_nl;
  wire[8:0] nl_inp_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_nl;
  wire[0:0] FpAdd_8U_23U_1_or_1_nl;
  wire[0:0] FpAdd_8U_23U_1_and_13_nl;
  wire[0:0] FpAdd_8U_23U_1_and_30_nl;
  wire[0:0] FpAdd_8U_23U_1_if_4_FpAdd_8U_23U_1_if_4_or_5_nl;
  wire[7:0] inp_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_nl;
  wire[8:0] nl_inp_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_nl;
  wire[0:0] FpAdd_8U_23U_1_or_2_nl;
  wire[0:0] FpAdd_8U_23U_1_and_19_nl;
  wire[0:0] FpAdd_8U_23U_1_and_32_nl;
  wire[0:0] FpAdd_8U_23U_1_if_4_FpAdd_8U_23U_1_if_4_or_6_nl;
  wire[7:0] inp_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_nl;
  wire[8:0] nl_inp_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_nl;
  wire[0:0] FpAdd_8U_23U_1_or_3_nl;
  wire[0:0] FpAdd_8U_23U_1_and_25_nl;
  wire[0:0] FpAdd_8U_23U_1_and_34_nl;
  wire[0:0] FpAdd_8U_23U_1_if_4_FpAdd_8U_23U_1_if_4_or_7_nl;
  wire[0:0] inp_lookup_1_FpMantDecShiftRight_23U_8U_10U_carry_and_nl;
  wire[22:0] inp_lookup_1_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl;
  wire[23:0] nl_inp_lookup_1_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl;
  wire[5:0] inp_lookup_1_FpAdd_6U_10U_1_if_3_if_acc_1_nl;
  wire[6:0] nl_inp_lookup_1_FpAdd_6U_10U_1_if_3_if_acc_1_nl;
  wire[5:0] inp_lookup_1_FpNormalize_6U_23U_1_else_acc_nl;
  wire[7:0] nl_inp_lookup_1_FpNormalize_6U_23U_1_else_acc_nl;
  wire[0:0] inp_lookup_2_FpMantDecShiftRight_23U_8U_10U_carry_and_nl;
  wire[22:0] inp_lookup_2_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl;
  wire[23:0] nl_inp_lookup_2_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl;
  wire[5:0] inp_lookup_2_FpAdd_6U_10U_1_if_3_if_acc_1_nl;
  wire[6:0] nl_inp_lookup_2_FpAdd_6U_10U_1_if_3_if_acc_1_nl;
  wire[5:0] inp_lookup_2_FpNormalize_6U_23U_1_else_acc_nl;
  wire[7:0] nl_inp_lookup_2_FpNormalize_6U_23U_1_else_acc_nl;
  wire[0:0] inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_carry_and_nl;
  wire[22:0] inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl;
  wire[23:0] nl_inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl;
  wire[5:0] inp_lookup_3_FpAdd_6U_10U_1_if_3_if_acc_1_nl;
  wire[6:0] nl_inp_lookup_3_FpAdd_6U_10U_1_if_3_if_acc_1_nl;
  wire[5:0] inp_lookup_3_FpNormalize_6U_23U_1_else_acc_nl;
  wire[7:0] nl_inp_lookup_3_FpNormalize_6U_23U_1_else_acc_nl;
  wire[0:0] inp_lookup_4_FpMantDecShiftRight_23U_8U_10U_carry_and_nl;
  wire[22:0] inp_lookup_4_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl;
  wire[23:0] nl_inp_lookup_4_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl;
  wire[5:0] inp_lookup_4_FpAdd_6U_10U_1_if_3_if_acc_1_nl;
  wire[6:0] nl_inp_lookup_4_FpAdd_6U_10U_1_if_3_if_acc_1_nl;
  wire[5:0] inp_lookup_4_FpNormalize_6U_23U_1_else_acc_nl;
  wire[7:0] nl_inp_lookup_4_FpNormalize_6U_23U_1_else_acc_nl;
  wire[7:0] inp_lookup_1_FpMul_6U_10U_oelse_1_acc_nl;
  wire[8:0] nl_inp_lookup_1_FpMul_6U_10U_oelse_1_acc_nl;
  wire[7:0] inp_lookup_2_FpMul_6U_10U_oelse_1_acc_nl;
  wire[8:0] nl_inp_lookup_2_FpMul_6U_10U_oelse_1_acc_nl;
  wire[7:0] inp_lookup_3_FpMul_6U_10U_oelse_1_acc_nl;
  wire[8:0] nl_inp_lookup_3_FpMul_6U_10U_oelse_1_acc_nl;
  wire[7:0] inp_lookup_4_FpMul_6U_10U_oelse_1_acc_nl;
  wire[8:0] nl_inp_lookup_4_FpMul_6U_10U_oelse_1_acc_nl;
  wire[5:0] inp_lookup_1_FpMul_6U_10U_else_2_else_if_if_acc_1_nl;
  wire[6:0] nl_inp_lookup_1_FpMul_6U_10U_else_2_else_if_if_acc_1_nl;
  wire[5:0] inp_lookup_2_FpMul_6U_10U_else_2_else_if_if_acc_1_nl;
  wire[6:0] nl_inp_lookup_2_FpMul_6U_10U_else_2_else_if_if_acc_1_nl;
  wire[5:0] inp_lookup_3_FpMul_6U_10U_else_2_else_if_if_acc_1_nl;
  wire[6:0] nl_inp_lookup_3_FpMul_6U_10U_else_2_else_if_if_acc_1_nl;
  wire[5:0] inp_lookup_4_FpMul_6U_10U_else_2_else_if_if_acc_1_nl;
  wire[6:0] nl_inp_lookup_4_FpMul_6U_10U_else_2_else_if_if_acc_1_nl;
  wire[0:0] or_5860_nl;
  wire[0:0] IsNaN_6U_23U_aelse_not_8_nl;
  wire[0:0] FpNormalize_6U_23U_oelse_not_16_nl;
  wire[5:0] inp_lookup_1_FpNormalize_6U_23U_else_acc_nl;
  wire[7:0] nl_inp_lookup_1_FpNormalize_6U_23U_else_acc_nl;
  wire[0:0] FpNormalize_6U_23U_oelse_not_8_nl;
  wire[0:0] FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_nl;
  wire[5:0] inp_lookup_1_FpAdd_6U_10U_if_4_if_acc_1_nl;
  wire[6:0] nl_inp_lookup_1_FpAdd_6U_10U_if_4_if_acc_1_nl;
  wire[9:0] FpAdd_6U_10U_FpAdd_6U_10U_or_4_nl;
  wire[9:0] inp_lookup_1_FpMantRNE_23U_11U_else_acc_nl;
  wire[10:0] nl_inp_lookup_1_FpMantRNE_23U_11U_else_acc_nl;
  wire[0:0] or_5861_nl;
  wire[0:0] IsNaN_6U_23U_aelse_not_9_nl;
  wire[0:0] FpNormalize_6U_23U_oelse_not_17_nl;
  wire[5:0] inp_lookup_2_FpNormalize_6U_23U_else_acc_nl;
  wire[7:0] nl_inp_lookup_2_FpNormalize_6U_23U_else_acc_nl;
  wire[0:0] FpNormalize_6U_23U_oelse_not_10_nl;
  wire[0:0] FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_1_nl;
  wire[5:0] inp_lookup_2_FpAdd_6U_10U_if_4_if_acc_1_nl;
  wire[6:0] nl_inp_lookup_2_FpAdd_6U_10U_if_4_if_acc_1_nl;
  wire[9:0] FpAdd_6U_10U_FpAdd_6U_10U_or_6_nl;
  wire[9:0] inp_lookup_2_FpMantRNE_23U_11U_else_acc_nl;
  wire[10:0] nl_inp_lookup_2_FpMantRNE_23U_11U_else_acc_nl;
  wire[0:0] or_5862_nl;
  wire[0:0] IsNaN_6U_23U_aelse_not_10_nl;
  wire[0:0] FpNormalize_6U_23U_oelse_not_18_nl;
  wire[5:0] inp_lookup_3_FpNormalize_6U_23U_else_acc_nl;
  wire[7:0] nl_inp_lookup_3_FpNormalize_6U_23U_else_acc_nl;
  wire[0:0] FpNormalize_6U_23U_oelse_not_12_nl;
  wire[0:0] FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_2_nl;
  wire[5:0] inp_lookup_3_FpAdd_6U_10U_if_4_if_acc_1_nl;
  wire[6:0] nl_inp_lookup_3_FpAdd_6U_10U_if_4_if_acc_1_nl;
  wire[9:0] FpAdd_6U_10U_FpAdd_6U_10U_or_8_nl;
  wire[9:0] inp_lookup_3_FpMantRNE_23U_11U_else_acc_nl;
  wire[10:0] nl_inp_lookup_3_FpMantRNE_23U_11U_else_acc_nl;
  wire[0:0] or_5863_nl;
  wire[0:0] IsNaN_6U_23U_aelse_not_11_nl;
  wire[0:0] FpNormalize_6U_23U_oelse_not_19_nl;
  wire[5:0] inp_lookup_4_FpNormalize_6U_23U_else_acc_nl;
  wire[7:0] nl_inp_lookup_4_FpNormalize_6U_23U_else_acc_nl;
  wire[0:0] FpNormalize_6U_23U_oelse_not_14_nl;
  wire[0:0] FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_3_nl;
  wire[5:0] inp_lookup_4_FpAdd_6U_10U_if_4_if_acc_1_nl;
  wire[6:0] nl_inp_lookup_4_FpAdd_6U_10U_if_4_if_acc_1_nl;
  wire[9:0] FpAdd_6U_10U_FpAdd_6U_10U_or_10_nl;
  wire[9:0] inp_lookup_4_FpMantRNE_23U_11U_else_acc_nl;
  wire[10:0] nl_inp_lookup_4_FpMantRNE_23U_11U_else_acc_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_23_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_25_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_27_nl;
  wire[0:0] FpAdd_8U_23U_is_a_greater_oelse_not_29_nl;
  wire[0:0] inp_lookup_1_IntSignedShiftRight_50U_5U_32U_obits_fixed_and_nl;
  wire[0:0] mux_1980_nl;
  wire[0:0] inp_lookup_2_IntSignedShiftRight_50U_5U_32U_obits_fixed_and_nl;
  wire[0:0] mux_1981_nl;
  wire[0:0] nor_707_nl;
  wire[0:0] or_5639_nl;
  wire[0:0] inp_lookup_3_IntSignedShiftRight_50U_5U_32U_obits_fixed_and_nl;
  wire[0:0] mux_1982_nl;
  wire[0:0] nor_706_nl;
  wire[0:0] or_5638_nl;
  wire[0:0] inp_lookup_4_IntSignedShiftRight_50U_5U_32U_obits_fixed_and_nl;
  wire[0:0] mux_1983_nl;
  wire[0:0] nor_705_nl;
  wire[0:0] or_5637_nl;
  wire[0:0] mux_1984_nl;
  wire[5:0] inp_lookup_1_FpMul_6U_10U_2_else_2_else_if_if_acc_nl;
  wire[6:0] nl_inp_lookup_1_FpMul_6U_10U_2_else_2_else_if_if_acc_nl;
  wire[0:0] FpMul_6U_10U_2_or_4_nl;
  wire[0:0] FpMantWidthDec_6U_21U_10U_0U_0U_2_and_1_nl;
  wire[0:0] mux_1985_nl;
  wire[0:0] nor_704_nl;
  wire[0:0] or_5636_nl;
  wire[5:0] inp_lookup_2_FpMul_6U_10U_2_else_2_else_if_if_acc_nl;
  wire[6:0] nl_inp_lookup_2_FpMul_6U_10U_2_else_2_else_if_if_acc_nl;
  wire[0:0] FpMul_6U_10U_2_or_5_nl;
  wire[0:0] FpMantWidthDec_6U_21U_10U_0U_0U_2_and_3_nl;
  wire[0:0] mux_1986_nl;
  wire[5:0] inp_lookup_3_FpMul_6U_10U_2_else_2_else_if_if_acc_nl;
  wire[6:0] nl_inp_lookup_3_FpMul_6U_10U_2_else_2_else_if_if_acc_nl;
  wire[0:0] FpMul_6U_10U_2_or_6_nl;
  wire[0:0] FpMantWidthDec_6U_21U_10U_0U_0U_2_and_5_nl;
  wire[0:0] mux_1987_nl;
  wire[5:0] inp_lookup_4_FpMul_6U_10U_2_else_2_else_if_if_acc_nl;
  wire[6:0] nl_inp_lookup_4_FpMul_6U_10U_2_else_2_else_if_if_acc_nl;
  wire[0:0] FpMul_6U_10U_2_or_7_nl;
  wire[0:0] FpMantWidthDec_6U_21U_10U_0U_0U_2_and_7_nl;
  wire[7:0] inp_lookup_1_FpAdd_8U_23U_1_b_right_shift_qif_acc_nl;
  wire[9:0] nl_inp_lookup_1_FpAdd_8U_23U_1_b_right_shift_qif_acc_nl;
  wire[7:0] inp_lookup_1_FpAdd_8U_23U_1_a_right_shift_qelse_acc_nl;
  wire[8:0] nl_inp_lookup_1_FpAdd_8U_23U_1_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_8U_23U_1_is_a_greater_oelse_not_23_nl;
  wire[7:0] inp_lookup_2_FpAdd_8U_23U_1_b_right_shift_qif_acc_nl;
  wire[9:0] nl_inp_lookup_2_FpAdd_8U_23U_1_b_right_shift_qif_acc_nl;
  wire[7:0] inp_lookup_2_FpAdd_8U_23U_1_a_right_shift_qelse_acc_nl;
  wire[8:0] nl_inp_lookup_2_FpAdd_8U_23U_1_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_8U_23U_1_is_a_greater_oelse_not_25_nl;
  wire[7:0] inp_lookup_3_FpAdd_8U_23U_1_b_right_shift_qif_acc_nl;
  wire[9:0] nl_inp_lookup_3_FpAdd_8U_23U_1_b_right_shift_qif_acc_nl;
  wire[7:0] inp_lookup_3_FpAdd_8U_23U_1_a_right_shift_qelse_acc_nl;
  wire[8:0] nl_inp_lookup_3_FpAdd_8U_23U_1_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_8U_23U_1_is_a_greater_oelse_not_27_nl;
  wire[7:0] inp_lookup_4_FpAdd_8U_23U_1_b_right_shift_qif_acc_nl;
  wire[9:0] nl_inp_lookup_4_FpAdd_8U_23U_1_b_right_shift_qif_acc_nl;
  wire[7:0] inp_lookup_4_FpAdd_8U_23U_1_a_right_shift_qelse_acc_nl;
  wire[8:0] nl_inp_lookup_4_FpAdd_8U_23U_1_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_8U_23U_1_is_a_greater_oelse_not_29_nl;
  wire[0:0] FpAdd_6U_10U_1_if_4_FpAdd_6U_10U_1_if_4_or_nl;
  wire[0:0] FpAdd_6U_10U_1_if_4_FpAdd_6U_10U_1_if_4_or_1_nl;
  wire[0:0] FpAdd_6U_10U_1_if_4_FpAdd_6U_10U_1_if_4_or_2_nl;
  wire[0:0] FpAdd_6U_10U_1_if_4_FpAdd_6U_10U_1_if_4_or_3_nl;
  wire[5:0] inp_lookup_1_FpMul_6U_10U_else_2_else_if_if_acc_nl;
  wire[6:0] nl_inp_lookup_1_FpMul_6U_10U_else_2_else_if_if_acc_nl;
  wire[0:0] nand_643_nl;
  wire[0:0] FpMul_6U_10U_FpMul_6U_10U_nor_8_nl;
  wire[0:0] FpMul_6U_10U_or_4_nl;
  wire[0:0] FpMantWidthDec_6U_21U_10U_0U_0U_and_1_nl;
  wire[5:0] inp_lookup_2_FpMul_6U_10U_else_2_else_if_if_acc_nl;
  wire[6:0] nl_inp_lookup_2_FpMul_6U_10U_else_2_else_if_if_acc_nl;
  wire[0:0] nand_642_nl;
  wire[0:0] FpMul_6U_10U_FpMul_6U_10U_nor_9_nl;
  wire[0:0] FpMul_6U_10U_or_5_nl;
  wire[0:0] FpMantWidthDec_6U_21U_10U_0U_0U_and_3_nl;
  wire[5:0] inp_lookup_3_FpMul_6U_10U_else_2_else_if_if_acc_nl;
  wire[6:0] nl_inp_lookup_3_FpMul_6U_10U_else_2_else_if_if_acc_nl;
  wire[0:0] nand_641_nl;
  wire[0:0] FpMul_6U_10U_FpMul_6U_10U_nor_10_nl;
  wire[0:0] FpMul_6U_10U_or_6_nl;
  wire[0:0] FpMantWidthDec_6U_21U_10U_0U_0U_and_5_nl;
  wire[5:0] inp_lookup_4_FpMul_6U_10U_else_2_else_if_if_acc_nl;
  wire[6:0] nl_inp_lookup_4_FpMul_6U_10U_else_2_else_if_if_acc_nl;
  wire[0:0] nand_640_nl;
  wire[0:0] FpMul_6U_10U_FpMul_6U_10U_nor_11_nl;
  wire[0:0] FpMul_6U_10U_or_7_nl;
  wire[0:0] FpMantWidthDec_6U_21U_10U_0U_0U_and_7_nl;
  wire[2:0] inp_lookup_1_IntSaturation_51U_32U_else_if_acc_nl;
  wire[3:0] nl_inp_lookup_1_IntSaturation_51U_32U_else_if_acc_nl;
  wire[2:0] inp_lookup_2_IntSaturation_51U_32U_else_if_acc_nl;
  wire[3:0] nl_inp_lookup_2_IntSaturation_51U_32U_else_if_acc_nl;
  wire[2:0] inp_lookup_3_IntSaturation_51U_32U_else_if_acc_nl;
  wire[3:0] nl_inp_lookup_3_IntSaturation_51U_32U_else_if_acc_nl;
  wire[2:0] inp_lookup_4_IntSaturation_51U_32U_else_if_acc_nl;
  wire[3:0] nl_inp_lookup_4_IntSaturation_51U_32U_else_if_acc_nl;
  wire[51:0] inp_lookup_1_else_else_b0_mul_nl;
  wire signed [52:0] nl_inp_lookup_1_else_else_b0_mul_nl;
  wire[51:0] inp_lookup_2_else_else_b0_mul_nl;
  wire signed [52:0] nl_inp_lookup_2_else_else_b0_mul_nl;
  wire[51:0] inp_lookup_3_else_else_b0_mul_nl;
  wire signed [52:0] nl_inp_lookup_3_else_else_b0_mul_nl;
  wire[51:0] inp_lookup_4_else_else_b0_mul_nl;
  wire signed [52:0] nl_inp_lookup_4_else_else_b0_mul_nl;
  wire[8:0] inp_lookup_1_FpNormalize_8U_49U_1_acc_nl;
  wire[10:0] nl_inp_lookup_1_FpNormalize_8U_49U_1_acc_nl;
  wire[8:0] inp_lookup_2_FpNormalize_8U_49U_1_acc_nl;
  wire[10:0] nl_inp_lookup_2_FpNormalize_8U_49U_1_acc_nl;
  wire[8:0] inp_lookup_3_FpNormalize_8U_49U_1_acc_nl;
  wire[10:0] nl_inp_lookup_3_FpNormalize_8U_49U_1_acc_nl;
  wire[8:0] inp_lookup_4_FpNormalize_8U_49U_1_acc_nl;
  wire[10:0] nl_inp_lookup_4_FpNormalize_8U_49U_1_acc_nl;
  wire[6:0] inp_lookup_1_FpNormalize_6U_23U_1_acc_nl;
  wire[8:0] nl_inp_lookup_1_FpNormalize_6U_23U_1_acc_nl;
  wire[6:0] inp_lookup_2_FpNormalize_6U_23U_1_acc_nl;
  wire[8:0] nl_inp_lookup_2_FpNormalize_6U_23U_1_acc_nl;
  wire[6:0] inp_lookup_3_FpNormalize_6U_23U_1_acc_nl;
  wire[8:0] nl_inp_lookup_3_FpNormalize_6U_23U_1_acc_nl;
  wire[6:0] inp_lookup_4_FpNormalize_6U_23U_1_acc_nl;
  wire[8:0] nl_inp_lookup_4_FpNormalize_6U_23U_1_acc_nl;
  wire[0:0] mux_106_nl;
  wire[0:0] and_3402_nl;
  wire[0:0] nor_1710_nl;
  wire[0:0] mux_204_nl;
  wire[0:0] nor_1640_nl;
  wire[0:0] and_132_nl;
  wire[0:0] mux_203_nl;
  wire[0:0] or_454_nl;
  wire[0:0] or_506_nl;
  wire[0:0] mux_242_nl;
  wire[0:0] and_138_nl;
  wire[0:0] mux_240_nl;
  wire[0:0] or_515_nl;
  wire[0:0] or_570_nl;
  wire[0:0] mux_280_nl;
  wire[0:0] mux_278_nl;
  wire[0:0] and_145_nl;
  wire[0:0] or_577_nl;
  wire[0:0] mux_322_nl;
  wire[0:0] mux_321_nl;
  wire[0:0] mux_324_nl;
  wire[0:0] mux_323_nl;
  wire[0:0] or_635_nl;
  wire[0:0] nand_22_nl;
  wire[0:0] mux_326_nl;
  wire[0:0] nand_23_nl;
  wire[0:0] mux_327_nl;
  wire[0:0] or_636_nl;
  wire[0:0] mux_337_nl;
  wire[0:0] or_645_nl;
  wire[0:0] or_647_nl;
  wire[0:0] mux_339_nl;
  wire[0:0] or_968_nl;
  wire[0:0] or_970_nl;
  wire[0:0] nand_568_nl;
  wire[0:0] or_999_nl;
  wire[0:0] mux_502_nl;
  wire[0:0] nand_566_nl;
  wire[0:0] or_1018_nl;
  wire[0:0] or_1022_nl;
  wire[0:0] or_1043_nl;
  wire[0:0] or_1045_nl;
  wire[0:0] or_1280_nl;
  wire[0:0] or_1306_nl;
  wire[0:0] nor_1476_nl;
  wire[0:0] mux_636_nl;
  wire[0:0] and_3289_nl;
  wire[0:0] mux_638_nl;
  wire[0:0] mux_637_nl;
  wire[0:0] nor_1477_nl;
  wire[0:0] or_1319_nl;
  wire[0:0] or_1686_nl;
  wire[0:0] or_1752_nl;
  wire[0:0] or_1805_nl;
  wire[0:0] mux_857_nl;
  wire[0:0] nor_1382_nl;
  wire[0:0] or_5698_nl;
  wire[0:0] or_1866_nl;
  wire[0:0] mux_874_nl;
  wire[0:0] nor_1369_nl;
  wire[0:0] or_5697_nl;
  wire[0:0] or_1904_nl;
  wire[0:0] mux_891_nl;
  wire[0:0] nor_1356_nl;
  wire[0:0] or_5696_nl;
  wire[0:0] or_1942_nl;
  wire[0:0] or_2361_nl;
  wire[0:0] or_2362_nl;
  wire[0:0] or_2398_nl;
  wire[0:0] or_2399_nl;
  wire[0:0] or_2400_nl;
  wire[0:0] or_2401_nl;
  wire[0:0] mux_1057_nl;
  wire[0:0] nor_1175_nl;
  wire[0:0] nor_1176_nl;
  wire[0:0] or_2507_nl;
  wire[0:0] or_2508_nl;
  wire[0:0] nor_1155_nl;
  wire[0:0] nor_1157_nl;
  wire[0:0] mux_1087_nl;
  wire[0:0] or_2509_nl;
  wire[0:0] nand_135_nl;
  wire[0:0] or_2528_nl;
  wire[0:0] or_2530_nl;
  wire[0:0] mux_1100_nl;
  wire[0:0] mux_1099_nl;
  wire[0:0] or_2535_nl;
  wire[0:0] or_2536_nl;
  wire[0:0] or_2544_nl;
  wire[0:0] or_2545_nl;
  wire[0:0] nor_1147_nl;
  wire[0:0] nor_1149_nl;
  wire[0:0] mux_1104_nl;
  wire[0:0] or_2546_nl;
  wire[0:0] nand_139_nl;
  wire[0:0] or_2565_nl;
  wire[0:0] or_2567_nl;
  wire[0:0] mux_1117_nl;
  wire[0:0] mux_1116_nl;
  wire[0:0] or_2572_nl;
  wire[0:0] or_2573_nl;
  wire[0:0] or_2581_nl;
  wire[0:0] or_2582_nl;
  wire[0:0] nor_1139_nl;
  wire[0:0] nor_1141_nl;
  wire[0:0] mux_1121_nl;
  wire[0:0] or_2583_nl;
  wire[0:0] nand_143_nl;
  wire[0:0] or_2602_nl;
  wire[0:0] or_2604_nl;
  wire[0:0] mux_1134_nl;
  wire[0:0] mux_1133_nl;
  wire[0:0] or_2609_nl;
  wire[0:0] or_2610_nl;
  wire[0:0] nor_1131_nl;
  wire[0:0] nor_1133_nl;
  wire[0:0] mux_1138_nl;
  wire[0:0] or_2619_nl;
  wire[0:0] or_2621_nl;
  wire[0:0] or_2640_nl;
  wire[0:0] or_2642_nl;
  wire[0:0] mux_1152_nl;
  wire[0:0] mux_1151_nl;
  wire[0:0] or_2698_nl;
  wire[0:0] mux_1171_nl;
  wire[0:0] or_2701_nl;
  wire[0:0] or_2699_nl;
  wire[0:0] mux_1176_nl;
  wire[0:0] mux_1178_nl;
  wire[0:0] or_2714_nl;
  wire[0:0] mux_1177_nl;
  wire[0:0] and_3195_nl;
  wire[0:0] mux_1180_nl;
  wire[0:0] mux_1181_nl;
  wire[0:0] mux_1236_nl;
  wire[0:0] and_3400_nl;
  wire[0:0] nor_1058_nl;
  wire[0:0] mux_1238_nl;
  wire[0:0] and_3399_nl;
  wire[0:0] nor_1056_nl;
  wire[0:0] mux_1240_nl;
  wire[0:0] and_3398_nl;
  wire[0:0] nor_1054_nl;
  wire[0:0] mux_1242_nl;
  wire[0:0] and_3175_nl;
  wire[0:0] nor_1052_nl;
  wire[0:0] or_3150_nl;
  wire[0:0] or_3198_nl;
  wire[0:0] or_3219_nl;
  wire[0:0] or_3337_nl;
  wire[0:0] or_3339_nl;
  wire[0:0] mux_1449_nl;
  wire[0:0] or_3472_nl;
  wire[0:0] and_3122_nl;
  wire[0:0] nor_500_nl;
  wire[0:0] or_3478_nl;
  wire[0:0] or_3480_nl;
  wire[0:0] mux_1694_nl;
  wire[0:0] or_3781_nl;
  wire[0:0] mux_1821_nl;
  wire[0:0] or_3998_nl;
  wire[0:0] mux_1825_nl;
  wire[0:0] or_4001_nl;
  wire[0:0] nor_689_nl;
  wire[0:0] nor_691_nl;
  wire[0:0] nand_241_nl;
  wire[0:0] and_3053_nl;
  wire[0:0] nor_692_nl;
  wire[0:0] nor_696_nl;
  wire[0:0] mux_1922_nl;
  wire[0:0] mux_1921_nl;
  wire[0:0] mux_1920_nl;
  wire[0:0] nor_725_nl;
  wire[0:0] or_4697_nl;
  wire[0:0] or_4702_nl;
  wire[23:0] FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_nl;
  wire[25:0] nl_FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_nl;
  wire[23:0] FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_1_nl;
  wire[25:0] nl_FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_1_nl;
  wire[23:0] FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_2_nl;
  wire[25:0] nl_FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_2_nl;
  wire[23:0] FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_3_nl;
  wire[25:0] nl_FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_3_nl;
  wire[10:0] FpAdd_6U_10U_is_a_greater_oif_aelse_acc_nl;
  wire[12:0] nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_nl;
  wire[10:0] FpAdd_6U_10U_is_a_greater_oif_aelse_acc_1_nl;
  wire[12:0] nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_1_nl;
  wire[10:0] FpAdd_6U_10U_is_a_greater_oif_aelse_acc_2_nl;
  wire[12:0] nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_2_nl;
  wire[10:0] FpAdd_6U_10U_is_a_greater_oif_aelse_acc_3_nl;
  wire[12:0] nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_3_nl;
  wire[0:0] mux_2130_nl;
  wire[0:0] and_4121_nl;
  wire[0:0] mux_2131_nl;
  wire[0:0] and_4120_nl;
  wire[0:0] mux_2132_nl;
  wire[0:0] and_4119_nl;
  wire[0:0] mux_2133_nl;
  wire[0:0] and_4118_nl;
  wire[50:0] acc_nl;
  wire[51:0] nl_acc_nl;
  wire[48:0] FpAdd_8U_23U_if_2_mux_8_nl;
  wire[0:0] FpAdd_8U_23U_if_2_FpAdd_8U_23U_if_2_nand_4_nl;
  wire[48:0] FpAdd_8U_23U_if_2_mux_9_nl;
  wire[50:0] acc_1_nl;
  wire[51:0] nl_acc_1_nl;
  wire[48:0] FpAdd_8U_23U_if_2_mux_10_nl;
  wire[0:0] FpAdd_8U_23U_if_2_FpAdd_8U_23U_if_2_nand_5_nl;
  wire[48:0] FpAdd_8U_23U_if_2_mux_11_nl;
  wire[50:0] acc_2_nl;
  wire[51:0] nl_acc_2_nl;
  wire[48:0] FpAdd_8U_23U_if_2_mux_12_nl;
  wire[0:0] FpAdd_8U_23U_if_2_FpAdd_8U_23U_if_2_nand_6_nl;
  wire[48:0] FpAdd_8U_23U_if_2_mux_13_nl;
  wire[50:0] acc_3_nl;
  wire[51:0] nl_acc_3_nl;
  wire[48:0] FpAdd_8U_23U_if_2_mux_14_nl;
  wire[0:0] FpAdd_8U_23U_if_2_FpAdd_8U_23U_if_2_nand_7_nl;
  wire[48:0] FpAdd_8U_23U_if_2_mux_15_nl;
  wire[8:0] acc_4_nl;
  wire[9:0] nl_acc_4_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_8_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_9_nl;
  wire[8:0] acc_5_nl;
  wire[9:0] nl_acc_5_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_10_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_11_nl;
  wire[8:0] acc_6_nl;
  wire[9:0] nl_acc_6_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_12_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_13_nl;
  wire[8:0] acc_7_nl;
  wire[9:0] nl_acc_7_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_14_nl;
  wire[7:0] FpAdd_8U_23U_b_right_shift_qif_mux_15_nl;
  wire[0:0] FpMul_6U_10U_oelse_1_FpMul_6U_10U_oelse_1_or_4_nl;
  wire[0:0] FpMul_6U_10U_oelse_1_mux_28_nl;
  wire[3:0] FpMul_6U_10U_oelse_1_mux_29_nl;
  wire[0:0] FpMul_6U_10U_oelse_1_FpMul_6U_10U_oelse_1_or_5_nl;
  wire[0:0] FpMul_6U_10U_oelse_1_mux_30_nl;
  wire[3:0] FpMul_6U_10U_oelse_1_mux_31_nl;
  wire[0:0] FpMul_6U_10U_oelse_1_FpMul_6U_10U_oelse_1_or_6_nl;
  wire[0:0] FpMul_6U_10U_oelse_1_mux_32_nl;
  wire[3:0] FpMul_6U_10U_oelse_1_mux_33_nl;
  wire[0:0] FpMul_6U_10U_oelse_1_FpMul_6U_10U_oelse_1_or_7_nl;
  wire[0:0] FpMul_6U_10U_oelse_1_mux_34_nl;
  wire[3:0] FpMul_6U_10U_oelse_1_mux_35_nl;
  wire[6:0] acc_12_nl;
  wire[7:0] nl_acc_12_nl;
  wire[0:0] FpAdd_6U_10U_a_right_shift_qelse_mux_24_nl;
  wire[0:0] FpAdd_6U_10U_a_right_shift_qelse_mux_25_nl;
  wire[3:0] FpAdd_6U_10U_a_right_shift_qelse_mux_26_nl;
  wire[0:0] FpAdd_6U_10U_a_right_shift_qelse_mux_27_nl;
  wire[0:0] FpAdd_6U_10U_a_right_shift_qelse_mux_28_nl;
  wire[3:0] FpAdd_6U_10U_a_right_shift_qelse_mux_29_nl;
  wire[6:0] acc_13_nl;
  wire[7:0] nl_acc_13_nl;
  wire[0:0] FpAdd_6U_10U_a_right_shift_qelse_mux_30_nl;
  wire[0:0] FpAdd_6U_10U_a_right_shift_qelse_mux_31_nl;
  wire[3:0] FpAdd_6U_10U_a_right_shift_qelse_mux_32_nl;
  wire[0:0] FpAdd_6U_10U_a_right_shift_qelse_mux_33_nl;
  wire[0:0] FpAdd_6U_10U_a_right_shift_qelse_mux_34_nl;
  wire[3:0] FpAdd_6U_10U_a_right_shift_qelse_mux_35_nl;
  wire[6:0] acc_14_nl;
  wire[7:0] nl_acc_14_nl;
  wire[0:0] FpAdd_6U_10U_a_right_shift_qelse_mux_36_nl;
  wire[0:0] FpAdd_6U_10U_a_right_shift_qelse_mux_37_nl;
  wire[3:0] FpAdd_6U_10U_a_right_shift_qelse_mux_38_nl;
  wire[0:0] FpAdd_6U_10U_a_right_shift_qelse_mux_39_nl;
  wire[0:0] FpAdd_6U_10U_a_right_shift_qelse_mux_40_nl;
  wire[3:0] FpAdd_6U_10U_a_right_shift_qelse_mux_41_nl;
  wire[6:0] acc_15_nl;
  wire[7:0] nl_acc_15_nl;
  wire[0:0] FpAdd_6U_10U_a_right_shift_qelse_mux_42_nl;
  wire[0:0] FpAdd_6U_10U_a_right_shift_qelse_mux_43_nl;
  wire[3:0] FpAdd_6U_10U_a_right_shift_qelse_mux_44_nl;
  wire[0:0] FpAdd_6U_10U_a_right_shift_qelse_mux_45_nl;
  wire[0:0] FpAdd_6U_10U_a_right_shift_qelse_mux_46_nl;
  wire[3:0] FpAdd_6U_10U_a_right_shift_qelse_mux_47_nl;
// Interconnect Declarations for Component Instantiations
  wire [48:0] nl_inp_lookup_1_FpNormalize_8U_49U_else_lshift_rg_a;
  assign nl_inp_lookup_1_FpNormalize_8U_49U_else_lshift_rg_a = z_out[48:0];
  wire [48:0] nl_inp_lookup_2_FpNormalize_8U_49U_else_lshift_rg_a;
  assign nl_inp_lookup_2_FpNormalize_8U_49U_else_lshift_rg_a = z_out_1[48:0];
  wire [48:0] nl_inp_lookup_3_FpNormalize_8U_49U_else_lshift_rg_a;
  assign nl_inp_lookup_3_FpNormalize_8U_49U_else_lshift_rg_a = z_out_2[48:0];
  wire [48:0] nl_inp_lookup_4_FpNormalize_8U_49U_else_lshift_rg_a;
  assign nl_inp_lookup_4_FpNormalize_8U_49U_else_lshift_rg_a = z_out_3[48:0];
  wire [10:0] nl_inp_lookup_1_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_1_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_a = {IsZero_6U_10U_1_IsZero_6U_10U_1_and_itm_10
      , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_22};
  wire[5:0] inp_lookup_1_FpAdd_6U_10U_1_a_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl;
  wire[5:0] inp_lookup_1_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_inp_lookup_1_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_1_is_a_greater_oelse_not_23_nl;
  wire [7:0] nl_inp_lookup_1_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_s;
  assign nl_inp_lookup_1_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl = ({FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_7_5_1
      , FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_7_4_1 , FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_7_3_0_1})
      + ({(~ FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_6_5_1) , (~ FpAdd_8U_23U_1_o_sign_1_lpi_1_dfm_5)
      , (~ FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_6_3_0_1)}) + 6'b1;
  assign inp_lookup_1_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl = nl_inp_lookup_1_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_1_is_a_greater_oelse_not_23_nl = ~ FpAdd_6U_10U_1_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0;
  assign inp_lookup_1_FpAdd_6U_10U_1_a_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (inp_lookup_1_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_1_is_a_greater_oelse_not_23_nl)));
  assign nl_inp_lookup_1_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_s = ({1'b1 , (inp_lookup_1_FpAdd_6U_10U_1_a_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_inp_lookup_1_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_1_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_a = {inp_lookup_1_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_itm_3
      , reg_FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_7_itm , reg_FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_7_1_itm};
  wire[5:0] inp_lookup_1_FpAdd_6U_10U_1_b_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl;
  wire[5:0] inp_lookup_1_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl;
  wire[7:0] nl_inp_lookup_1_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl;
  wire [7:0] nl_inp_lookup_1_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_s;
  assign nl_inp_lookup_1_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl = ({FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_6_5_1
      , FpAdd_8U_23U_1_o_sign_1_lpi_1_dfm_5 , FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_6_3_0_1})
      + ({(~ FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_7_5_1) , (~ FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_7_4_1)
      , (~ FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_7_3_0_1)}) + 6'b1;
  assign inp_lookup_1_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl = nl_inp_lookup_1_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl[5:0];
  assign inp_lookup_1_FpAdd_6U_10U_1_b_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (inp_lookup_1_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_1_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0));
  assign nl_inp_lookup_1_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_s = ({1'b1 , (inp_lookup_1_FpAdd_6U_10U_1_b_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_inp_lookup_2_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_2_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_a = {IsZero_6U_10U_1_IsZero_6U_10U_1_and_1_itm_8
      , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_22};
  wire[5:0] inp_lookup_2_FpAdd_6U_10U_1_a_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl;
  wire[5:0] inp_lookup_2_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_inp_lookup_2_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_1_is_a_greater_oelse_not_25_nl;
  wire [7:0] nl_inp_lookup_2_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_s;
  assign nl_inp_lookup_2_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl = ({FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_7_5_1
      , FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_7_4_1 , FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_7_3_0_1})
      + ({(~ FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_6_5_1) , (~ FpAdd_8U_23U_1_o_sign_2_lpi_1_dfm_5)
      , (~ FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_6_3_0_1)}) + 6'b1;
  assign inp_lookup_2_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl = nl_inp_lookup_2_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_1_is_a_greater_oelse_not_25_nl = ~ FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0;
  assign inp_lookup_2_FpAdd_6U_10U_1_a_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (inp_lookup_2_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_1_is_a_greater_oelse_not_25_nl)));
  assign nl_inp_lookup_2_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_s = ({1'b1 , (inp_lookup_2_FpAdd_6U_10U_1_a_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_inp_lookup_2_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_2_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_a = {inp_lookup_2_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_itm_3
      , reg_FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_7_itm , reg_FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_7_1_itm};
  wire[5:0] inp_lookup_2_FpAdd_6U_10U_1_b_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl;
  wire[5:0] inp_lookup_2_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl;
  wire[7:0] nl_inp_lookup_2_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl;
  wire [7:0] nl_inp_lookup_2_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_s;
  assign nl_inp_lookup_2_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl = ({FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_6_5_1
      , FpAdd_8U_23U_1_o_sign_2_lpi_1_dfm_5 , FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_6_3_0_1})
      + ({(~ FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_7_5_1) , (~ FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_7_4_1)
      , (~ FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_7_3_0_1)}) + 6'b1;
  assign inp_lookup_2_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl = nl_inp_lookup_2_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl[5:0];
  assign inp_lookup_2_FpAdd_6U_10U_1_b_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (inp_lookup_2_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0));
  assign nl_inp_lookup_2_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_s = ({1'b1 , (inp_lookup_2_FpAdd_6U_10U_1_b_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_inp_lookup_3_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_3_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_a = {IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_itm_10
      , reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_6_itm , reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_6_1_itm};
  wire[5:0] inp_lookup_3_FpAdd_6U_10U_1_a_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl;
  wire[5:0] inp_lookup_3_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_inp_lookup_3_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_1_is_a_greater_oelse_not_27_nl;
  wire [7:0] nl_inp_lookup_3_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_s;
  assign nl_inp_lookup_3_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl = ({FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_7_5_1
      , FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_7_4_1 , FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_7_3_0_1})
      + ({(~ FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_6_5_1) , (~ FpAdd_8U_23U_1_o_sign_3_lpi_1_dfm_5)
      , (~ FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_6_3_0_1)}) + 6'b1;
  assign inp_lookup_3_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl = nl_inp_lookup_3_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_1_is_a_greater_oelse_not_27_nl = ~ FpAdd_6U_10U_1_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0;
  assign inp_lookup_3_FpAdd_6U_10U_1_a_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (inp_lookup_3_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_1_is_a_greater_oelse_not_27_nl)));
  assign nl_inp_lookup_3_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_s = ({1'b1 , (inp_lookup_3_FpAdd_6U_10U_1_a_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_inp_lookup_3_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_3_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_a = {inp_lookup_3_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_itm_3
      , reg_FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_7_itm , reg_FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_7_1_itm};
  wire[5:0] inp_lookup_3_FpAdd_6U_10U_1_b_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl;
  wire[5:0] inp_lookup_3_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl;
  wire[7:0] nl_inp_lookup_3_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl;
  wire [7:0] nl_inp_lookup_3_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_s;
  assign nl_inp_lookup_3_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl = ({FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_6_5_1
      , FpAdd_8U_23U_1_o_sign_3_lpi_1_dfm_5 , FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_6_3_0_1})
      + ({(~ FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_7_5_1) , (~ FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_7_4_1)
      , (~ FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_7_3_0_1)}) + 6'b1;
  assign inp_lookup_3_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl = nl_inp_lookup_3_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl[5:0];
  assign inp_lookup_3_FpAdd_6U_10U_1_b_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (inp_lookup_3_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_1_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0));
  assign nl_inp_lookup_3_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_s = ({1'b1 , (inp_lookup_3_FpAdd_6U_10U_1_b_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_inp_lookup_4_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_4_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_a = {IsZero_6U_10U_1_IsZero_6U_10U_1_and_3_itm_8
      , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_22};
  wire[5:0] inp_lookup_4_FpAdd_6U_10U_1_a_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl;
  wire[5:0] inp_lookup_4_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl;
  wire[7:0] nl_inp_lookup_4_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl;
  wire[0:0] FpAdd_6U_10U_1_is_a_greater_oelse_not_29_nl;
  wire [7:0] nl_inp_lookup_4_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_s;
  assign nl_inp_lookup_4_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl = ({FpMul_6U_10U_2_o_expo_lpi_1_dfm_7_5_1
      , FpMul_6U_10U_2_o_expo_lpi_1_dfm_7_4_1 , FpMul_6U_10U_2_o_expo_lpi_1_dfm_7_3_0_1})
      + ({(~ FpMul_6U_10U_1_o_expo_lpi_1_dfm_6_5_1) , (~ FpAdd_8U_23U_1_o_sign_lpi_1_dfm_5)
      , (~ FpMul_6U_10U_1_o_expo_lpi_1_dfm_6_3_0_1)}) + 6'b1;
  assign inp_lookup_4_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl = nl_inp_lookup_4_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl[5:0];
  assign FpAdd_6U_10U_1_is_a_greater_oelse_not_29_nl = ~ FpAdd_6U_10U_1_is_a_greater_lor_lpi_1_dfm_1_mx0w0;
  assign inp_lookup_4_FpAdd_6U_10U_1_a_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (inp_lookup_4_FpAdd_6U_10U_1_a_right_shift_qelse_acc_nl),
      (FpAdd_6U_10U_1_is_a_greater_oelse_not_29_nl)));
  assign nl_inp_lookup_4_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_s = ({1'b1 , (inp_lookup_4_FpAdd_6U_10U_1_a_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_inp_lookup_4_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_4_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_a = {inp_lookup_4_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_itm_3
      , reg_FpMul_6U_10U_2_o_mant_lpi_1_dfm_7_reg , reg_FpMul_6U_10U_2_o_mant_lpi_1_dfm_7_1_reg};
  wire[5:0] inp_lookup_4_FpAdd_6U_10U_1_b_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl;
  wire[5:0] inp_lookup_4_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl;
  wire[7:0] nl_inp_lookup_4_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl;
  wire [7:0] nl_inp_lookup_4_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_s;
  assign nl_inp_lookup_4_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl = ({FpMul_6U_10U_1_o_expo_lpi_1_dfm_6_5_1
      , FpAdd_8U_23U_1_o_sign_lpi_1_dfm_5 , FpMul_6U_10U_1_o_expo_lpi_1_dfm_6_3_0_1})
      + ({(~ FpMul_6U_10U_2_o_expo_lpi_1_dfm_7_5_1) , (~ FpMul_6U_10U_2_o_expo_lpi_1_dfm_7_4_1)
      , (~ FpMul_6U_10U_2_o_expo_lpi_1_dfm_7_3_0_1)}) + 6'b1;
  assign inp_lookup_4_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl = nl_inp_lookup_4_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl[5:0];
  assign inp_lookup_4_FpAdd_6U_10U_1_b_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, (inp_lookup_4_FpAdd_6U_10U_1_b_right_shift_qif_acc_nl),
      FpAdd_6U_10U_1_is_a_greater_lor_lpi_1_dfm_1_mx0w0));
  assign nl_inp_lookup_4_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_s = ({1'b1 , (inp_lookup_4_FpAdd_6U_10U_1_b_left_shift_FpAdd_6U_10U_1_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_inp_lookup_1_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_1_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a = {inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_16
      , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_24};
  wire[5:0] inp_lookup_1_FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl;
  wire[0:0] FpAdd_6U_10U_is_a_greater_oelse_not_23_nl;
  wire [7:0] nl_inp_lookup_1_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_s;
  assign FpAdd_6U_10U_is_a_greater_oelse_not_23_nl = ~ FpAdd_6U_10U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0;
  assign inp_lookup_1_FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, z_out_12, (FpAdd_6U_10U_is_a_greater_oelse_not_23_nl)));
  assign nl_inp_lookup_1_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_s = ({1'b1 , (inp_lookup_1_FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_inp_lookup_1_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_1_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a = {inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_3_or_itm_2
      , FpMul_6U_10U_o_mant_1_lpi_1_dfm_7};
  wire[5:0] inp_lookup_1_FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl;
  wire [7:0] nl_inp_lookup_1_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_s;
  assign inp_lookup_1_FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, z_out_12, FpAdd_6U_10U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0));
  assign nl_inp_lookup_1_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_s = ({1'b1 , (inp_lookup_1_FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_inp_lookup_2_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_2_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a = {inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_15
      , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_24};
  wire[5:0] inp_lookup_2_FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl;
  wire[0:0] FpAdd_6U_10U_is_a_greater_oelse_not_25_nl;
  wire [7:0] nl_inp_lookup_2_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_s;
  assign FpAdd_6U_10U_is_a_greater_oelse_not_25_nl = ~ FpAdd_6U_10U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0;
  assign inp_lookup_2_FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, z_out_13, (FpAdd_6U_10U_is_a_greater_oelse_not_25_nl)));
  assign nl_inp_lookup_2_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_s = ({1'b1 , (inp_lookup_2_FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_inp_lookup_2_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_2_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a = {inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_3_or_itm_2
      , FpMul_6U_10U_o_mant_2_lpi_1_dfm_7};
  wire[5:0] inp_lookup_2_FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl;
  wire [7:0] nl_inp_lookup_2_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_s;
  assign inp_lookup_2_FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, z_out_13, FpAdd_6U_10U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0));
  assign nl_inp_lookup_2_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_s = ({1'b1 , (inp_lookup_2_FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_inp_lookup_3_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_3_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a = {inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_16
      , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_27};
  wire[5:0] inp_lookup_3_FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl;
  wire[0:0] FpAdd_6U_10U_is_a_greater_oelse_not_27_nl;
  wire [7:0] nl_inp_lookup_3_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_s;
  assign FpAdd_6U_10U_is_a_greater_oelse_not_27_nl = ~ FpAdd_6U_10U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0;
  assign inp_lookup_3_FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, z_out_14, (FpAdd_6U_10U_is_a_greater_oelse_not_27_nl)));
  assign nl_inp_lookup_3_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_s = ({1'b1 , (inp_lookup_3_FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_inp_lookup_3_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_3_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a = {inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_3_or_itm_2
      , FpMul_6U_10U_o_mant_3_lpi_1_dfm_7};
  wire[5:0] inp_lookup_3_FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl;
  wire [7:0] nl_inp_lookup_3_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_s;
  assign inp_lookup_3_FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, z_out_14, FpAdd_6U_10U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0));
  assign nl_inp_lookup_3_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_s = ({1'b1 , (inp_lookup_3_FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_inp_lookup_4_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_4_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a = {inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_16
      , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_24};
  wire[5:0] inp_lookup_4_FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl;
  wire[0:0] FpAdd_6U_10U_is_a_greater_oelse_not_29_nl;
  wire [7:0] nl_inp_lookup_4_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_s;
  assign FpAdd_6U_10U_is_a_greater_oelse_not_29_nl = ~ FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_1_mx0w0;
  assign inp_lookup_4_FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, z_out_15, (FpAdd_6U_10U_is_a_greater_oelse_not_29_nl)));
  assign nl_inp_lookup_4_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_s = ({1'b1 , (inp_lookup_4_FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [10:0] nl_inp_lookup_4_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_4_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a = {inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_3_or_itm_2
      , FpMul_6U_10U_o_mant_lpi_1_dfm_7};
  wire[5:0] inp_lookup_4_FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl;
  wire [7:0] nl_inp_lookup_4_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_s;
  assign inp_lookup_4_FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl
      = ~(MUX_v_6_2_2(6'b000000, z_out_15, FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_1_mx0w0));
  assign nl_inp_lookup_4_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_s = ({1'b1 , (inp_lookup_4_FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl)})
      + 7'b1101;
  wire [34:0] nl_inp_lookup_1_leading_sign_35_0_1_rg_mantissa;
  assign nl_inp_lookup_1_leading_sign_35_0_1_rg_mantissa = chn_inp_in_rsci_d_mxwt[162:128];
  wire [34:0] nl_inp_lookup_2_leading_sign_35_0_1_rg_mantissa;
  assign nl_inp_lookup_2_leading_sign_35_0_1_rg_mantissa = chn_inp_in_rsci_d_mxwt[197:163];
  wire [34:0] nl_inp_lookup_3_leading_sign_35_0_1_rg_mantissa;
  assign nl_inp_lookup_3_leading_sign_35_0_1_rg_mantissa = chn_inp_in_rsci_d_mxwt[232:198];
  wire [34:0] nl_inp_lookup_4_leading_sign_35_0_1_rg_mantissa;
  assign nl_inp_lookup_4_leading_sign_35_0_1_rg_mantissa = chn_inp_in_rsci_d_mxwt[267:233];
  wire [23:0] nl_inp_lookup_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a = {inp_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2
      , (chn_inp_in_crt_sva_1_739_395_1[235:213])};
  wire[7:0] inp_lookup_1_FpAdd_8U_23U_b_left_shift_acc_nl;
  wire[8:0] nl_inp_lookup_1_FpAdd_8U_23U_b_left_shift_acc_nl;
  wire [8:0] nl_inp_lookup_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s;
  assign nl_inp_lookup_1_FpAdd_8U_23U_b_left_shift_acc_nl = ({1'b1 , (~ (FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign inp_lookup_1_FpAdd_8U_23U_b_left_shift_acc_nl = nl_inp_lookup_1_FpAdd_8U_23U_b_left_shift_acc_nl[7:0];
  assign nl_inp_lookup_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s = {(inp_lookup_1_FpAdd_8U_23U_b_left_shift_acc_nl)
      , (~ (FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm[0]))};
  wire [23:0] nl_inp_lookup_2_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_2_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a = {IsZero_6U_10U_7_IsZero_6U_10U_7_and_1_itm_2
      , (chn_inp_in_crt_sva_1_739_395_1[267:245])};
  wire[7:0] inp_lookup_2_FpAdd_8U_23U_b_left_shift_acc_nl;
  wire[8:0] nl_inp_lookup_2_FpAdd_8U_23U_b_left_shift_acc_nl;
  wire [8:0] nl_inp_lookup_2_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s;
  assign nl_inp_lookup_2_FpAdd_8U_23U_b_left_shift_acc_nl = ({1'b1 , (~ (FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign inp_lookup_2_FpAdd_8U_23U_b_left_shift_acc_nl = nl_inp_lookup_2_FpAdd_8U_23U_b_left_shift_acc_nl[7:0];
  assign nl_inp_lookup_2_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s = {(inp_lookup_2_FpAdd_8U_23U_b_left_shift_acc_nl)
      , (~ (FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm[0]))};
  wire [23:0] nl_inp_lookup_3_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_3_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a = {inp_lookup_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2
      , (chn_inp_in_crt_sva_1_739_395_1[299:277])};
  wire[7:0] inp_lookup_3_FpAdd_8U_23U_b_left_shift_acc_nl;
  wire[8:0] nl_inp_lookup_3_FpAdd_8U_23U_b_left_shift_acc_nl;
  wire [8:0] nl_inp_lookup_3_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s;
  assign nl_inp_lookup_3_FpAdd_8U_23U_b_left_shift_acc_nl = ({1'b1 , (~ (FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign inp_lookup_3_FpAdd_8U_23U_b_left_shift_acc_nl = nl_inp_lookup_3_FpAdd_8U_23U_b_left_shift_acc_nl[7:0];
  assign nl_inp_lookup_3_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s = {(inp_lookup_3_FpAdd_8U_23U_b_left_shift_acc_nl)
      , (~ (FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm[0]))};
  wire [23:0] nl_inp_lookup_4_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_4_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a = {IsZero_6U_10U_7_IsZero_6U_10U_7_and_3_itm_2
      , (chn_inp_in_crt_sva_1_739_395_1[331:309])};
  wire[7:0] inp_lookup_4_FpAdd_8U_23U_b_left_shift_acc_nl;
  wire[8:0] nl_inp_lookup_4_FpAdd_8U_23U_b_left_shift_acc_nl;
  wire [8:0] nl_inp_lookup_4_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s;
  assign nl_inp_lookup_4_FpAdd_8U_23U_b_left_shift_acc_nl = ({1'b1 , (~ (FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign inp_lookup_4_FpAdd_8U_23U_b_left_shift_acc_nl = nl_inp_lookup_4_FpAdd_8U_23U_b_left_shift_acc_nl[7:0];
  assign nl_inp_lookup_4_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s = {(inp_lookup_4_FpAdd_8U_23U_b_left_shift_acc_nl)
      , (~ (FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm[0]))};
  wire [8:0] nl_inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg_a;
  assign nl_inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg_a = chn_inp_in_rsci_d_mxwt[356:348];
  wire [5:0] nl_inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg_s;
  assign nl_inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg_s = conv_u2u_4_5(libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_17)
      + 5'b1;
  wire [8:0] nl_inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg_a;
  assign nl_inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg_a = chn_inp_in_rsci_d_mxwt[388:380];
  wire [5:0] nl_inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg_s;
  assign nl_inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg_s = conv_u2u_4_5(libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_19)
      + 5'b1;
  wire [8:0] nl_inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_a;
  assign nl_inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_a = chn_inp_in_rsci_d_mxwt[308:300];
  wire [5:0] nl_inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_s;
  assign nl_inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_s = conv_u2u_4_5(libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_22)
      + 5'b1;
  wire [8:0] nl_inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_a = chn_inp_in_rsci_d_mxwt[420:412];
  wire [5:0] nl_inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_s = conv_u2u_4_5(libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_25)
      + 5'b1;
  wire [8:0] nl_inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_a;
  assign nl_inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_a = chn_inp_in_rsci_d_mxwt[452:444];
  wire [5:0] nl_inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_s;
  assign nl_inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_s = conv_u2u_4_5(libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_27)
      + 5'b1;
  wire [8:0] nl_inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_a;
  assign nl_inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_a = chn_inp_in_rsci_d_mxwt[276:268];
  wire [5:0] nl_inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_s;
  assign nl_inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_s = conv_u2u_4_5(libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_20)
      + 5'b1;
  wire [8:0] nl_inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_a;
  assign nl_inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_a = chn_inp_in_rsci_d_mxwt[292:284];
  wire [5:0] nl_inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_s;
  assign nl_inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_s = conv_u2u_4_5(libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_21)
      + 5'b1;
  wire [8:0] nl_inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_a;
  assign nl_inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_a = chn_inp_in_rsci_d_mxwt[324:316];
  wire [5:0] nl_inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_s;
  assign nl_inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_s = conv_u2u_4_5(libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_23)
      + 5'b1;
  wire [34:0] nl_inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg_a;
  assign nl_inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg_a
      = chn_inp_in_rsci_d_mxwt[162:128];
  wire [7:0] nl_inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg_s;
  assign nl_inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg_s
      = conv_u2u_6_7(libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_12)
      + 7'b1;
  wire [34:0] nl_inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg_a;
  assign nl_inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg_a
      = chn_inp_in_rsci_d_mxwt[197:163];
  wire [7:0] nl_inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg_s;
  assign nl_inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg_s
      = conv_u2u_6_7(libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_13)
      + 7'b1;
  wire [34:0] nl_inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg_a;
  assign nl_inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg_a
      = chn_inp_in_rsci_d_mxwt[232:198];
  wire [7:0] nl_inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg_s;
  assign nl_inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg_s
      = conv_u2u_6_7(libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_14)
      + 7'b1;
  wire [34:0] nl_inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg_a;
  assign nl_inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg_a
      = chn_inp_in_rsci_d_mxwt[267:233];
  wire [7:0] nl_inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg_s;
  assign nl_inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg_s
      = conv_u2u_6_7(libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_15)
      + 7'b1;
  wire [34:0] nl_inp_lookup_1_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg_a;
  assign nl_inp_lookup_1_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg_a
      = {reg_inp_lookup_1_else_else_a0_acc_1_reg , reg_inp_lookup_1_else_else_a0_acc_2_reg};
  wire [7:0] nl_inp_lookup_1_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg_s;
  assign nl_inp_lookup_1_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg_s
      = conv_u2u_6_7(IntLeadZero_35U_leading_sign_35_0_rtn_1_sva_2) + 7'b1;
  wire [34:0] nl_inp_lookup_2_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg_a;
  assign nl_inp_lookup_2_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg_a
      = {reg_inp_lookup_2_else_else_a0_acc_1_reg , reg_inp_lookup_2_else_else_a0_acc_2_reg};
  wire [7:0] nl_inp_lookup_2_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg_s;
  assign nl_inp_lookup_2_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg_s
      = conv_u2u_6_7(IntLeadZero_35U_leading_sign_35_0_rtn_2_sva_2) + 7'b1;
  wire [34:0] nl_inp_lookup_3_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg_a;
  assign nl_inp_lookup_3_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg_a
      = {reg_inp_lookup_3_else_else_a0_acc_1_reg , reg_inp_lookup_3_else_else_a0_acc_2_reg};
  wire [7:0] nl_inp_lookup_3_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg_s;
  assign nl_inp_lookup_3_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg_s
      = conv_u2u_6_7(IntLeadZero_35U_leading_sign_35_0_rtn_3_sva_2) + 7'b1;
  wire [34:0] nl_inp_lookup_4_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg_a;
  assign nl_inp_lookup_4_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg_a
      = {reg_inp_lookup_4_else_else_a0_acc_1_reg , reg_inp_lookup_4_else_else_a0_acc_2_reg};
  wire [7:0] nl_inp_lookup_4_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg_s;
  assign nl_inp_lookup_4_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg_s
      = conv_u2u_6_7(IntLeadZero_35U_leading_sign_35_0_rtn_sva_2) + 7'b1;
  wire [48:0] nl_inp_lookup_1_leading_sign_49_0_rg_mantissa;
  assign nl_inp_lookup_1_leading_sign_49_0_rg_mantissa = z_out[48:0];
  wire [48:0] nl_inp_lookup_2_leading_sign_49_0_rg_mantissa;
  assign nl_inp_lookup_2_leading_sign_49_0_rg_mantissa = z_out_1[48:0];
  wire [48:0] nl_inp_lookup_3_leading_sign_49_0_rg_mantissa;
  assign nl_inp_lookup_3_leading_sign_49_0_rg_mantissa = z_out_2[48:0];
  wire [48:0] nl_inp_lookup_4_leading_sign_49_0_rg_mantissa;
  assign nl_inp_lookup_4_leading_sign_49_0_rg_mantissa = z_out_3[48:0];
  wire [48:0] nl_inp_lookup_1_leading_sign_49_0_1_rg_mantissa;
  assign nl_inp_lookup_1_leading_sign_49_0_1_rg_mantissa = FpAdd_8U_23U_1_int_mant_p1_1_sva_3[48:0];
  wire [48:0] nl_inp_lookup_1_FpNormalize_8U_49U_1_else_lshift_rg_a;
  assign nl_inp_lookup_1_FpNormalize_8U_49U_1_else_lshift_rg_a = FpAdd_8U_23U_1_int_mant_p1_1_sva_3[48:0];
  wire [48:0] nl_inp_lookup_2_leading_sign_49_0_1_rg_mantissa;
  assign nl_inp_lookup_2_leading_sign_49_0_1_rg_mantissa = FpAdd_8U_23U_1_int_mant_p1_2_sva_3[48:0];
  wire [48:0] nl_inp_lookup_2_FpNormalize_8U_49U_1_else_lshift_rg_a;
  assign nl_inp_lookup_2_FpNormalize_8U_49U_1_else_lshift_rg_a = FpAdd_8U_23U_1_int_mant_p1_2_sva_3[48:0];
  wire [48:0] nl_inp_lookup_3_leading_sign_49_0_1_rg_mantissa;
  assign nl_inp_lookup_3_leading_sign_49_0_1_rg_mantissa = FpAdd_8U_23U_1_int_mant_p1_3_sva_3[48:0];
  wire [48:0] nl_inp_lookup_3_FpNormalize_8U_49U_1_else_lshift_rg_a;
  assign nl_inp_lookup_3_FpNormalize_8U_49U_1_else_lshift_rg_a = FpAdd_8U_23U_1_int_mant_p1_3_sva_3[48:0];
  wire [48:0] nl_inp_lookup_4_leading_sign_49_0_1_rg_mantissa;
  assign nl_inp_lookup_4_leading_sign_49_0_1_rg_mantissa = FpAdd_8U_23U_1_int_mant_p1_sva_3[48:0];
  wire [48:0] nl_inp_lookup_4_FpNormalize_8U_49U_1_else_lshift_rg_a;
  assign nl_inp_lookup_4_FpNormalize_8U_49U_1_else_lshift_rg_a = FpAdd_8U_23U_1_int_mant_p1_sva_3[48:0];
  wire [23:0] nl_inp_lookup_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_a;
  assign nl_inp_lookup_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_a = {1'b1
      , FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_6};
  wire [3:0] nl_inp_lookup_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_s;
  assign nl_inp_lookup_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_s = {reg_FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_8_3_0_1_itm
      , (~ (FpAdd_6U_10U_1_qr_2_lpi_1_dfm_5[0]))};
  wire [5:0] nl_inp_lookup_1_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg_s;
  assign nl_inp_lookup_1_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg_s =
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_1_sva_2 + 5'b11111;
  wire [22:0] nl_inp_lookup_1_FpNormalize_6U_23U_1_else_lshift_rg_a;
  assign nl_inp_lookup_1_FpNormalize_6U_23U_1_else_lshift_rg_a = FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_4[22:0];
  wire [22:0] nl_inp_lookup_1_leading_sign_23_0_1_rg_mantissa;
  assign nl_inp_lookup_1_leading_sign_23_0_1_rg_mantissa = FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_4[22:0];
  wire [23:0] nl_inp_lookup_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_a;
  assign nl_inp_lookup_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_a = {1'b1
      , FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_6};
  wire [3:0] nl_inp_lookup_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_s;
  assign nl_inp_lookup_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_s = {reg_FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_8_3_0_1_itm
      , (~ (FpAdd_6U_10U_1_qr_3_lpi_1_dfm_5[0]))};
  wire [5:0] nl_inp_lookup_2_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg_s;
  assign nl_inp_lookup_2_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg_s =
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_2_sva_2 + 5'b11111;
  wire [22:0] nl_inp_lookup_2_FpNormalize_6U_23U_1_else_lshift_rg_a;
  assign nl_inp_lookup_2_FpNormalize_6U_23U_1_else_lshift_rg_a = FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_4[22:0];
  wire [22:0] nl_inp_lookup_2_leading_sign_23_0_1_rg_mantissa;
  assign nl_inp_lookup_2_leading_sign_23_0_1_rg_mantissa = FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_4[22:0];
  wire [23:0] nl_inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_a;
  assign nl_inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_a = {1'b1
      , FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_6};
  wire [3:0] nl_inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_s;
  assign nl_inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_s = {reg_FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_8_3_0_1_itm
      , (~ (FpAdd_6U_10U_1_qr_4_lpi_1_dfm_5[0]))};
  wire [5:0] nl_inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg_s;
  assign nl_inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg_s =
      reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_8_1_itm + 5'b11111;
  wire [22:0] nl_inp_lookup_3_FpNormalize_6U_23U_1_else_lshift_rg_a;
  assign nl_inp_lookup_3_FpNormalize_6U_23U_1_else_lshift_rg_a = FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_4[22:0];
  wire [22:0] nl_inp_lookup_3_leading_sign_23_0_1_rg_mantissa;
  assign nl_inp_lookup_3_leading_sign_23_0_1_rg_mantissa = FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_4[22:0];
  wire [23:0] nl_inp_lookup_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_a;
  assign nl_inp_lookup_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_a = {1'b1
      , FpAdd_8U_23U_1_o_mant_lpi_1_dfm_6};
  wire [3:0] nl_inp_lookup_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_s;
  assign nl_inp_lookup_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_s = {reg_FpMul_6U_10U_1_o_expo_lpi_1_dfm_8_3_0_1_itm
      , (~ (FpAdd_6U_10U_1_qr_lpi_1_dfm_5[0]))};
  wire [5:0] nl_inp_lookup_4_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg_s;
  assign nl_inp_lookup_4_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg_s =
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva_2 + 5'b11111;
  wire [22:0] nl_inp_lookup_4_FpNormalize_6U_23U_1_else_lshift_rg_a;
  assign nl_inp_lookup_4_FpNormalize_6U_23U_1_else_lshift_rg_a = FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_4[22:0];
  wire [22:0] nl_inp_lookup_4_leading_sign_23_0_1_rg_mantissa;
  assign nl_inp_lookup_4_leading_sign_23_0_1_rg_mantissa = FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_4[22:0];
  wire [22:0] nl_inp_lookup_1_FpNormalize_6U_23U_else_lshift_rg_a;
  assign nl_inp_lookup_1_FpNormalize_6U_23U_else_lshift_rg_a = FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_4[22:0];
  wire [22:0] nl_inp_lookup_2_FpNormalize_6U_23U_else_lshift_rg_a;
  assign nl_inp_lookup_2_FpNormalize_6U_23U_else_lshift_rg_a = FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_4[22:0];
  wire [22:0] nl_inp_lookup_3_FpNormalize_6U_23U_else_lshift_rg_a;
  assign nl_inp_lookup_3_FpNormalize_6U_23U_else_lshift_rg_a = FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_4[22:0];
  wire [22:0] nl_inp_lookup_4_FpNormalize_6U_23U_else_lshift_rg_a;
  assign nl_inp_lookup_4_FpNormalize_6U_23U_else_lshift_rg_a = FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_4[22:0];
  wire [9:0] nl_inp_lookup_1_leading_sign_10_0_3_rg_mantissa;
  assign nl_inp_lookup_1_leading_sign_10_0_3_rg_mantissa = chn_inp_in_rsci_d_mxwt[341:332];
  wire [9:0] nl_inp_lookup_2_leading_sign_10_0_3_rg_mantissa;
  assign nl_inp_lookup_2_leading_sign_10_0_3_rg_mantissa = chn_inp_in_rsci_d_mxwt[357:348];
  wire [9:0] nl_inp_lookup_3_leading_sign_10_0_3_rg_mantissa;
  assign nl_inp_lookup_3_leading_sign_10_0_3_rg_mantissa = chn_inp_in_rsci_d_mxwt[373:364];
  wire [9:0] nl_inp_lookup_4_leading_sign_10_0_3_rg_mantissa;
  assign nl_inp_lookup_4_leading_sign_10_0_3_rg_mantissa = chn_inp_in_rsci_d_mxwt[389:380];
  wire [23:0] nl_inp_lookup_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a = {inp_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_2
      , (chn_inp_in_crt_sva_1_739_395_1[107:85])};
  wire[7:0] inp_lookup_1_FpAdd_8U_23U_a_left_shift_acc_nl;
  wire[8:0] nl_inp_lookup_1_FpAdd_8U_23U_a_left_shift_acc_nl;
  wire [8:0] nl_inp_lookup_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s;
  assign nl_inp_lookup_1_FpAdd_8U_23U_a_left_shift_acc_nl = ({1'b1 , (~ (FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign inp_lookup_1_FpAdd_8U_23U_a_left_shift_acc_nl = nl_inp_lookup_1_FpAdd_8U_23U_a_left_shift_acc_nl[7:0];
  assign nl_inp_lookup_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s = {(inp_lookup_1_FpAdd_8U_23U_a_left_shift_acc_nl)
      , (~ (FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm[0]))};
  wire [23:0] nl_inp_lookup_2_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_2_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a = {inp_lookup_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_2
      , (chn_inp_in_crt_sva_1_739_395_1[139:117])};
  wire[7:0] inp_lookup_2_FpAdd_8U_23U_a_left_shift_acc_nl;
  wire[8:0] nl_inp_lookup_2_FpAdd_8U_23U_a_left_shift_acc_nl;
  wire [8:0] nl_inp_lookup_2_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s;
  assign nl_inp_lookup_2_FpAdd_8U_23U_a_left_shift_acc_nl = ({1'b1 , (~ (FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign inp_lookup_2_FpAdd_8U_23U_a_left_shift_acc_nl = nl_inp_lookup_2_FpAdd_8U_23U_a_left_shift_acc_nl[7:0];
  assign nl_inp_lookup_2_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s = {(inp_lookup_2_FpAdd_8U_23U_a_left_shift_acc_nl)
      , (~ (FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm[0]))};
  wire [23:0] nl_inp_lookup_3_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_3_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a = {inp_lookup_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_2
      , (chn_inp_in_crt_sva_1_739_395_1[171:149])};
  wire[7:0] inp_lookup_3_FpAdd_8U_23U_a_left_shift_acc_nl;
  wire[8:0] nl_inp_lookup_3_FpAdd_8U_23U_a_left_shift_acc_nl;
  wire [8:0] nl_inp_lookup_3_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s;
  assign nl_inp_lookup_3_FpAdd_8U_23U_a_left_shift_acc_nl = ({1'b1 , (~ (FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign inp_lookup_3_FpAdd_8U_23U_a_left_shift_acc_nl = nl_inp_lookup_3_FpAdd_8U_23U_a_left_shift_acc_nl[7:0];
  assign nl_inp_lookup_3_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s = {(inp_lookup_3_FpAdd_8U_23U_a_left_shift_acc_nl)
      , (~ (FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm[0]))};
  wire [23:0] nl_inp_lookup_4_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_4_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a = {inp_lookup_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_2
      , (chn_inp_in_crt_sva_1_739_395_1[203:181])};
  wire[7:0] inp_lookup_4_FpAdd_8U_23U_a_left_shift_acc_nl;
  wire[8:0] nl_inp_lookup_4_FpAdd_8U_23U_a_left_shift_acc_nl;
  wire [8:0] nl_inp_lookup_4_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s;
  assign nl_inp_lookup_4_FpAdd_8U_23U_a_left_shift_acc_nl = ({1'b1 , (~ (FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign inp_lookup_4_FpAdd_8U_23U_a_left_shift_acc_nl = nl_inp_lookup_4_FpAdd_8U_23U_a_left_shift_acc_nl[7:0];
  assign nl_inp_lookup_4_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s = {(inp_lookup_4_FpAdd_8U_23U_a_left_shift_acc_nl)
      , (~ (FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm[0]))};
  wire [23:0] nl_inp_lookup_1_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_1_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a = {inp_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2
      , FpAdd_8U_23U_o_mant_1_lpi_1_dfm_6};
  wire[7:0] inp_lookup_1_FpAdd_8U_23U_1_b_left_shift_acc_nl;
  wire[8:0] nl_inp_lookup_1_FpAdd_8U_23U_1_b_left_shift_acc_nl;
  wire [8:0] nl_inp_lookup_1_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s;
  assign nl_inp_lookup_1_FpAdd_8U_23U_1_b_left_shift_acc_nl = ({1'b1 , (~ (FpAdd_8U_23U_1_b_right_shift_qr_1_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign inp_lookup_1_FpAdd_8U_23U_1_b_left_shift_acc_nl = nl_inp_lookup_1_FpAdd_8U_23U_1_b_left_shift_acc_nl[7:0];
  assign nl_inp_lookup_1_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s = {(inp_lookup_1_FpAdd_8U_23U_1_b_left_shift_acc_nl)
      , (~ (FpAdd_8U_23U_1_b_right_shift_qr_1_lpi_1_dfm[0]))};
  wire [23:0] nl_inp_lookup_1_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_1_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a = {inp_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_7
      , (chn_inp_in_crt_sva_4_127_0_1[22:0])};
  wire[7:0] inp_lookup_1_FpAdd_8U_23U_1_a_left_shift_acc_nl;
  wire[8:0] nl_inp_lookup_1_FpAdd_8U_23U_1_a_left_shift_acc_nl;
  wire [8:0] nl_inp_lookup_1_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s;
  assign nl_inp_lookup_1_FpAdd_8U_23U_1_a_left_shift_acc_nl = ({1'b1 , (~ (FpAdd_8U_23U_1_a_right_shift_qr_1_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign inp_lookup_1_FpAdd_8U_23U_1_a_left_shift_acc_nl = nl_inp_lookup_1_FpAdd_8U_23U_1_a_left_shift_acc_nl[7:0];
  assign nl_inp_lookup_1_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s = {(inp_lookup_1_FpAdd_8U_23U_1_a_left_shift_acc_nl)
      , (~ (FpAdd_8U_23U_1_a_right_shift_qr_1_lpi_1_dfm[0]))};
  wire [23:0] nl_inp_lookup_2_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_2_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a = {inp_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2
      , FpAdd_8U_23U_o_mant_2_lpi_1_dfm_6};
  wire[7:0] inp_lookup_2_FpAdd_8U_23U_1_b_left_shift_acc_nl;
  wire[8:0] nl_inp_lookup_2_FpAdd_8U_23U_1_b_left_shift_acc_nl;
  wire [8:0] nl_inp_lookup_2_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s;
  assign nl_inp_lookup_2_FpAdd_8U_23U_1_b_left_shift_acc_nl = ({1'b1 , (~ (FpAdd_8U_23U_1_b_right_shift_qr_2_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign inp_lookup_2_FpAdd_8U_23U_1_b_left_shift_acc_nl = nl_inp_lookup_2_FpAdd_8U_23U_1_b_left_shift_acc_nl[7:0];
  assign nl_inp_lookup_2_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s = {(inp_lookup_2_FpAdd_8U_23U_1_b_left_shift_acc_nl)
      , (~ (FpAdd_8U_23U_1_b_right_shift_qr_2_lpi_1_dfm[0]))};
  wire [23:0] nl_inp_lookup_2_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_2_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a = {inp_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_6
      , (chn_inp_in_crt_sva_4_127_0_1[54:32])};
  wire[7:0] inp_lookup_2_FpAdd_8U_23U_1_a_left_shift_acc_nl;
  wire[8:0] nl_inp_lookup_2_FpAdd_8U_23U_1_a_left_shift_acc_nl;
  wire [8:0] nl_inp_lookup_2_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s;
  assign nl_inp_lookup_2_FpAdd_8U_23U_1_a_left_shift_acc_nl = ({1'b1 , (~ (FpAdd_8U_23U_1_a_right_shift_qr_2_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign inp_lookup_2_FpAdd_8U_23U_1_a_left_shift_acc_nl = nl_inp_lookup_2_FpAdd_8U_23U_1_a_left_shift_acc_nl[7:0];
  assign nl_inp_lookup_2_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s = {(inp_lookup_2_FpAdd_8U_23U_1_a_left_shift_acc_nl)
      , (~ (FpAdd_8U_23U_1_a_right_shift_qr_2_lpi_1_dfm[0]))};
  wire [23:0] nl_inp_lookup_3_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_3_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a = {inp_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2
      , FpAdd_8U_23U_o_mant_3_lpi_1_dfm_6};
  wire[7:0] inp_lookup_3_FpAdd_8U_23U_1_b_left_shift_acc_nl;
  wire[8:0] nl_inp_lookup_3_FpAdd_8U_23U_1_b_left_shift_acc_nl;
  wire [8:0] nl_inp_lookup_3_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s;
  assign nl_inp_lookup_3_FpAdd_8U_23U_1_b_left_shift_acc_nl = ({1'b1 , (~ (FpAdd_8U_23U_1_b_right_shift_qr_3_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign inp_lookup_3_FpAdd_8U_23U_1_b_left_shift_acc_nl = nl_inp_lookup_3_FpAdd_8U_23U_1_b_left_shift_acc_nl[7:0];
  assign nl_inp_lookup_3_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s = {(inp_lookup_3_FpAdd_8U_23U_1_b_left_shift_acc_nl)
      , (~ (FpAdd_8U_23U_1_b_right_shift_qr_3_lpi_1_dfm[0]))};
  wire [23:0] nl_inp_lookup_3_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_3_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a = {inp_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_7
      , (chn_inp_in_crt_sva_4_127_0_1[86:64])};
  wire[7:0] inp_lookup_3_FpAdd_8U_23U_1_a_left_shift_acc_nl;
  wire[8:0] nl_inp_lookup_3_FpAdd_8U_23U_1_a_left_shift_acc_nl;
  wire [8:0] nl_inp_lookup_3_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s;
  assign nl_inp_lookup_3_FpAdd_8U_23U_1_a_left_shift_acc_nl = ({1'b1 , (~ (FpAdd_8U_23U_1_a_right_shift_qr_3_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign inp_lookup_3_FpAdd_8U_23U_1_a_left_shift_acc_nl = nl_inp_lookup_3_FpAdd_8U_23U_1_a_left_shift_acc_nl[7:0];
  assign nl_inp_lookup_3_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s = {(inp_lookup_3_FpAdd_8U_23U_1_a_left_shift_acc_nl)
      , (~ (FpAdd_8U_23U_1_a_right_shift_qr_3_lpi_1_dfm[0]))};
  wire [23:0] nl_inp_lookup_4_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_4_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a = {inp_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2
      , FpAdd_8U_23U_o_mant_lpi_1_dfm_6};
  wire[7:0] inp_lookup_4_FpAdd_8U_23U_1_b_left_shift_acc_nl;
  wire[8:0] nl_inp_lookup_4_FpAdd_8U_23U_1_b_left_shift_acc_nl;
  wire [8:0] nl_inp_lookup_4_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s;
  assign nl_inp_lookup_4_FpAdd_8U_23U_1_b_left_shift_acc_nl = ({1'b1 , (~ (FpAdd_8U_23U_1_b_right_shift_qr_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign inp_lookup_4_FpAdd_8U_23U_1_b_left_shift_acc_nl = nl_inp_lookup_4_FpAdd_8U_23U_1_b_left_shift_acc_nl[7:0];
  assign nl_inp_lookup_4_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s = {(inp_lookup_4_FpAdd_8U_23U_1_b_left_shift_acc_nl)
      , (~ (FpAdd_8U_23U_1_b_right_shift_qr_lpi_1_dfm[0]))};
  wire [23:0] nl_inp_lookup_4_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a;
  assign nl_inp_lookup_4_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a = {inp_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_6
      , (chn_inp_in_crt_sva_4_127_0_1[118:96])};
  wire[7:0] inp_lookup_4_FpAdd_8U_23U_1_a_left_shift_acc_nl;
  wire[8:0] nl_inp_lookup_4_FpAdd_8U_23U_1_a_left_shift_acc_nl;
  wire [8:0] nl_inp_lookup_4_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s;
  assign nl_inp_lookup_4_FpAdd_8U_23U_1_a_left_shift_acc_nl = ({1'b1 , (~ (FpAdd_8U_23U_1_a_right_shift_qr_lpi_1_dfm[7:1]))})
      + 8'b1101;
  assign inp_lookup_4_FpAdd_8U_23U_1_a_left_shift_acc_nl = nl_inp_lookup_4_FpAdd_8U_23U_1_a_left_shift_acc_nl[7:0];
  assign nl_inp_lookup_4_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s = {(inp_lookup_4_FpAdd_8U_23U_1_a_left_shift_acc_nl)
      , (~ (FpAdd_8U_23U_1_a_right_shift_qr_lpi_1_dfm[0]))};
  wire [22:0] nl_inp_lookup_1_leading_sign_23_0_rg_mantissa;
  assign nl_inp_lookup_1_leading_sign_23_0_rg_mantissa = FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_mx0[22:0];
  wire [22:0] nl_inp_lookup_2_leading_sign_23_0_rg_mantissa;
  assign nl_inp_lookup_2_leading_sign_23_0_rg_mantissa = FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_mx0[22:0];
  wire [22:0] nl_inp_lookup_3_leading_sign_23_0_rg_mantissa;
  assign nl_inp_lookup_3_leading_sign_23_0_rg_mantissa = FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_mx0[22:0];
  wire [22:0] nl_inp_lookup_4_leading_sign_23_0_rg_mantissa;
  assign nl_inp_lookup_4_leading_sign_23_0_rg_mantissa = FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_mx0[22:0];
  wire[49:0] inp_lookup_1_if_else_b_mul_nl;
  wire [64:0] nl_inp_lookup_1_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg_a;
  assign inp_lookup_1_if_else_b_mul_nl = conv_s2u_50_50($signed((reg_inp_lookup_1_else_else_a0_acc_2_reg))
      * $signed((chn_inp_in_crt_sva_1_739_395_1[16:1])));
  assign nl_inp_lookup_1_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg_a =
      {(inp_lookup_1_if_else_b_mul_nl) , 15'b0};
  wire [4:0] nl_inp_lookup_1_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg_s;
  assign nl_inp_lookup_1_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg_s =
      chn_inp_in_crt_sva_1_739_395_1[69:65];
  wire[49:0] inp_lookup_2_if_else_b_mul_nl;
  wire [64:0] nl_inp_lookup_2_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg_a;
  assign inp_lookup_2_if_else_b_mul_nl = conv_s2u_50_50($signed((reg_inp_lookup_2_else_else_a0_acc_2_reg))
      * $signed((chn_inp_in_crt_sva_1_739_395_1[32:17])));
  assign nl_inp_lookup_2_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg_a =
      {(inp_lookup_2_if_else_b_mul_nl) , 15'b0};
  wire [4:0] nl_inp_lookup_2_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg_s;
  assign nl_inp_lookup_2_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg_s =
      chn_inp_in_crt_sva_1_739_395_1[74:70];
  wire[49:0] inp_lookup_3_if_else_b_mul_nl;
  wire [64:0] nl_inp_lookup_3_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg_a;
  assign inp_lookup_3_if_else_b_mul_nl = conv_s2u_50_50($signed((reg_inp_lookup_3_else_else_a0_acc_2_reg))
      * $signed((chn_inp_in_crt_sva_1_739_395_1[48:33])));
  assign nl_inp_lookup_3_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg_a =
      {(inp_lookup_3_if_else_b_mul_nl) , 15'b0};
  wire [4:0] nl_inp_lookup_3_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg_s;
  assign nl_inp_lookup_3_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg_s =
      chn_inp_in_crt_sva_1_739_395_1[79:75];
  wire[49:0] inp_lookup_4_if_else_b_mul_nl;
  wire [64:0] nl_inp_lookup_4_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg_a;
  assign inp_lookup_4_if_else_b_mul_nl = conv_s2u_50_50($signed((reg_inp_lookup_4_else_else_a0_acc_2_reg))
      * $signed((chn_inp_in_crt_sva_1_739_395_1[64:49])));
  assign nl_inp_lookup_4_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg_a =
      {(inp_lookup_4_if_else_b_mul_nl) , 15'b0};
  wire [4:0] nl_inp_lookup_4_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg_s;
  assign nl_inp_lookup_4_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg_s =
      chn_inp_in_crt_sva_1_739_395_1[84:80];
  wire [9:0] nl_inp_lookup_1_leading_sign_10_0_2_rg_mantissa;
  assign nl_inp_lookup_1_leading_sign_10_0_2_rg_mantissa = chn_inp_in_rsci_d_mxwt[277:268];
  wire [9:0] nl_inp_lookup_2_leading_sign_10_0_2_rg_mantissa;
  assign nl_inp_lookup_2_leading_sign_10_0_2_rg_mantissa = chn_inp_in_rsci_d_mxwt[293:284];
  wire [9:0] nl_inp_lookup_3_leading_sign_10_0_2_rg_mantissa;
  assign nl_inp_lookup_3_leading_sign_10_0_2_rg_mantissa = chn_inp_in_rsci_d_mxwt[309:300];
  wire [9:0] nl_inp_lookup_4_leading_sign_10_0_2_rg_mantissa;
  assign nl_inp_lookup_4_leading_sign_10_0_2_rg_mantissa = chn_inp_in_rsci_d_mxwt[325:316];
  wire [9:0] nl_inp_lookup_1_leading_sign_10_0_rg_mantissa;
  assign nl_inp_lookup_1_leading_sign_10_0_rg_mantissa = chn_inp_in_rsci_d_mxwt[405:396];
  wire [9:0] nl_inp_lookup_2_leading_sign_10_0_rg_mantissa;
  assign nl_inp_lookup_2_leading_sign_10_0_rg_mantissa = chn_inp_in_rsci_d_mxwt[421:412];
  wire [9:0] nl_inp_lookup_3_leading_sign_10_0_rg_mantissa;
  assign nl_inp_lookup_3_leading_sign_10_0_rg_mantissa = chn_inp_in_rsci_d_mxwt[437:428];
  wire [9:0] nl_inp_lookup_4_leading_sign_10_0_rg_mantissa;
  assign nl_inp_lookup_4_leading_sign_10_0_rg_mantissa = chn_inp_in_rsci_d_mxwt[453:444];
  wire [8:0] nl_inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg_a;
  assign nl_inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg_a = MUX_v_9_2_2((chn_inp_in_rsci_d_mxwt[340:332]),
      (chn_inp_in_rsci_d_mxwt[404:396]), FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_and_tmp);
  wire[4:0] inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_1_nl;
  wire[5:0] nl_inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_1_nl;
  wire[4:0] inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_1_nl;
  wire[5:0] nl_inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_1_nl;
  wire [4:0] nl_inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg_s;
  assign nl_inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_1_nl = conv_u2u_4_5(libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_24)
      + 5'b1;
  assign inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_1_nl = nl_inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_1_nl[4:0];
  assign nl_inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_1_nl = conv_u2u_4_5(libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_16)
      + 5'b1;
  assign inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_1_nl = nl_inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_1_nl[4:0];
  assign nl_inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg_s = MUX_v_5_2_2((inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_1_nl),
      (inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_1_nl), FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_and_tmp);
  wire [8:0] nl_inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg_a;
  assign nl_inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg_a = MUX_v_9_2_2((chn_inp_in_rsci_d_mxwt[372:364]),
      (chn_inp_in_rsci_d_mxwt[436:428]), FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_and_tmp_1);
  wire[4:0] inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_1_nl;
  wire[5:0] nl_inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_1_nl;
  wire[4:0] inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_1_nl;
  wire[5:0] nl_inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_1_nl;
  wire [4:0] nl_inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg_s;
  assign nl_inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_1_nl = conv_u2u_4_5(libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_26)
      + 5'b1;
  assign inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_1_nl = nl_inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_1_nl[4:0];
  assign nl_inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_1_nl = conv_u2u_4_5(libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_18)
      + 5'b1;
  assign inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_1_nl = nl_inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_1_nl[4:0];
  assign nl_inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg_s = MUX_v_5_2_2((inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_1_nl),
      (inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_1_nl), FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_and_tmp_1);
  wire [127:0] nl_NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_out_rsci_inst_chn_inp_out_rsci_d;
  assign nl_NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_out_rsci_inst_chn_inp_out_rsci_d
      = {chn_inp_out_rsci_d_127 , chn_inp_out_rsci_d_126_124 , chn_inp_out_rsci_d_123
      , chn_inp_out_rsci_d_122_119 , chn_inp_out_rsci_d_118_109 , chn_inp_out_rsci_d_108_106
      , chn_inp_out_rsci_d_105_97 , chn_inp_out_rsci_d_96 , chn_inp_out_rsci_d_95
      , chn_inp_out_rsci_d_94_92 , chn_inp_out_rsci_d_91 , chn_inp_out_rsci_d_90_87
      , chn_inp_out_rsci_d_86_77 , chn_inp_out_rsci_d_76_74 , chn_inp_out_rsci_d_73_65
      , chn_inp_out_rsci_d_64 , chn_inp_out_rsci_d_63 , chn_inp_out_rsci_d_62_60
      , chn_inp_out_rsci_d_59 , chn_inp_out_rsci_d_58_55 , chn_inp_out_rsci_d_54_45
      , chn_inp_out_rsci_d_44_42 , chn_inp_out_rsci_d_41_33 , chn_inp_out_rsci_d_32
      , chn_inp_out_rsci_d_31 , chn_inp_out_rsci_d_30_28 , chn_inp_out_rsci_d_27
      , chn_inp_out_rsci_d_26_23 , chn_inp_out_rsci_d_22_13 , chn_inp_out_rsci_d_12_10
      , chn_inp_out_rsci_d_9_1 , chn_inp_out_rsci_d_0};
  SDP_Y_INP_mgc_in_wire_v1 #(.rscid(32'sd2),
  .width(32'sd2)) cfg_precision_rsci (
      .d(cfg_precision_rsci_d),
      .z(cfg_precision_rsc_z)
    );
  SDP_Y_INP_leading_sign_35_0 inp_lookup_1_leading_sign_35_0_rg (
      .mantissa(inp_lookup_else_if_a0_frac_1_sva_mx0w0),
      .rtn(libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_8)
    );
  SDP_Y_INP_leading_sign_35_0 inp_lookup_2_leading_sign_35_0_rg (
      .mantissa(inp_lookup_else_if_a0_frac_2_sva_mx0w0),
      .rtn(libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_9)
    );
  SDP_Y_INP_leading_sign_35_0 inp_lookup_3_leading_sign_35_0_rg (
      .mantissa(inp_lookup_else_if_a0_frac_3_sva_mx0w0),
      .rtn(libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_10)
    );
  SDP_Y_INP_leading_sign_35_0 inp_lookup_4_leading_sign_35_0_rg (
      .mantissa(inp_lookup_else_if_a0_frac_sva_mx0w0),
      .rtn(libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_11)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) inp_lookup_1_FpNormalize_8U_49U_else_lshift_rg (
      .a(nl_inp_lookup_1_FpNormalize_8U_49U_else_lshift_rg_a[48:0]),
      .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_8),
      .z(inp_lookup_1_FpNormalize_8U_49U_else_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) inp_lookup_2_FpNormalize_8U_49U_else_lshift_rg (
      .a(nl_inp_lookup_2_FpNormalize_8U_49U_else_lshift_rg_a[48:0]),
      .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_9),
      .z(inp_lookup_2_FpNormalize_8U_49U_else_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) inp_lookup_3_FpNormalize_8U_49U_else_lshift_rg (
      .a(nl_inp_lookup_3_FpNormalize_8U_49U_else_lshift_rg_a[48:0]),
      .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_10),
      .z(inp_lookup_3_FpNormalize_8U_49U_else_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) inp_lookup_4_FpNormalize_8U_49U_else_lshift_rg (
      .a(nl_inp_lookup_4_FpNormalize_8U_49U_else_lshift_rg_a[48:0]),
      .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_11),
      .z(inp_lookup_4_FpNormalize_8U_49U_else_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) inp_lookup_1_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_1_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_inp_lookup_1_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(inp_lookup_1_FpAdd_6U_10U_1_a_int_mant_p1_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) inp_lookup_1_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_1_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_inp_lookup_1_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(inp_lookup_1_FpAdd_6U_10U_1_b_int_mant_p1_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) inp_lookup_2_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_2_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_inp_lookup_2_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(inp_lookup_2_FpAdd_6U_10U_1_a_int_mant_p1_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) inp_lookup_2_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_2_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_inp_lookup_2_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(inp_lookup_2_FpAdd_6U_10U_1_b_int_mant_p1_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) inp_lookup_3_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_3_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_inp_lookup_3_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(inp_lookup_3_FpAdd_6U_10U_1_a_int_mant_p1_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) inp_lookup_3_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_3_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_inp_lookup_3_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(inp_lookup_3_FpAdd_6U_10U_1_b_int_mant_p1_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) inp_lookup_4_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_4_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_inp_lookup_4_FpAdd_6U_10U_1_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(inp_lookup_4_FpAdd_6U_10U_1_a_int_mant_p1_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) inp_lookup_4_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_4_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_inp_lookup_4_FpAdd_6U_10U_1_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(inp_lookup_4_FpAdd_6U_10U_1_b_int_mant_p1_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) inp_lookup_1_FpAdd_6U_10U_a_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_1_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_inp_lookup_1_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(inp_lookup_1_FpAdd_6U_10U_a_int_mant_p1_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) inp_lookup_1_FpAdd_6U_10U_b_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_1_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_inp_lookup_1_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(inp_lookup_1_FpAdd_6U_10U_b_int_mant_p1_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) inp_lookup_2_FpAdd_6U_10U_a_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_2_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_inp_lookup_2_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(inp_lookup_2_FpAdd_6U_10U_a_int_mant_p1_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) inp_lookup_2_FpAdd_6U_10U_b_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_2_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_inp_lookup_2_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(inp_lookup_2_FpAdd_6U_10U_b_int_mant_p1_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) inp_lookup_3_FpAdd_6U_10U_a_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_3_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_inp_lookup_3_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(inp_lookup_3_FpAdd_6U_10U_a_int_mant_p1_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) inp_lookup_3_FpAdd_6U_10U_b_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_3_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_inp_lookup_3_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(inp_lookup_3_FpAdd_6U_10U_b_int_mant_p1_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) inp_lookup_4_FpAdd_6U_10U_a_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_4_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_inp_lookup_4_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_s[6:0]),
      .z(inp_lookup_4_FpAdd_6U_10U_a_int_mant_p1_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) inp_lookup_4_FpAdd_6U_10U_b_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_4_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(nl_inp_lookup_4_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_s[6:0]),
      .z(inp_lookup_4_FpAdd_6U_10U_b_int_mant_p1_lshift_itm)
    );
  SDP_Y_INP_leading_sign_35_0 inp_lookup_1_leading_sign_35_0_1_rg (
      .mantissa(nl_inp_lookup_1_leading_sign_35_0_1_rg_mantissa[34:0]),
      .rtn(libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_12)
    );
  SDP_Y_INP_leading_sign_35_0 inp_lookup_2_leading_sign_35_0_1_rg (
      .mantissa(nl_inp_lookup_2_leading_sign_35_0_1_rg_mantissa[34:0]),
      .rtn(libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_13)
    );
  SDP_Y_INP_leading_sign_35_0 inp_lookup_3_leading_sign_35_0_1_rg (
      .mantissa(nl_inp_lookup_3_leading_sign_35_0_1_rg_mantissa[34:0]),
      .rtn(libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_14)
    );
  SDP_Y_INP_leading_sign_35_0 inp_lookup_4_leading_sign_35_0_1_rg (
      .mantissa(nl_inp_lookup_4_leading_sign_35_0_1_rg_mantissa[34:0]),
      .rtn(libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_15)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) inp_lookup_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_inp_lookup_1_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_19_mx0w1)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) inp_lookup_2_FpAdd_8U_23U_b_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_2_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_inp_lookup_2_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_13_mx0w1)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) inp_lookup_3_FpAdd_8U_23U_b_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_3_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_inp_lookup_3_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_7_mx0w1)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) inp_lookup_4_FpAdd_8U_23U_b_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_4_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_inp_lookup_4_FpAdd_8U_23U_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_addend_larger_asn_1_mx0w1)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd9),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd10)) inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg
      (
      .a(nl_inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg_a[8:0]),
      .s(nl_inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg_s[4:0]),
      .z(inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd9),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd10)) inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg
      (
      .a(nl_inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg_a[8:0]),
      .s(nl_inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg_s[4:0]),
      .z(inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd9),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd10)) inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg
      (
      .a(nl_inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_a[8:0]),
      .s(nl_inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_s[4:0]),
      .z(inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd9),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd10)) inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg
      (
      .a(nl_inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_a[8:0]),
      .s(nl_inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_s[4:0]),
      .z(inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd9),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd10)) inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg
      (
      .a(nl_inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_a[8:0]),
      .s(nl_inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_rg_s[4:0]),
      .z(inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd9),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd10)) inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg
      (
      .a(nl_inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_a[8:0]),
      .s(nl_inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_s[4:0]),
      .z(inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd9),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd10)) inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg
      (
      .a(nl_inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_a[8:0]),
      .s(nl_inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_s[4:0]),
      .z(inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd9),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd10)) inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg
      (
      .a(nl_inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_a[8:0]),
      .s(nl_inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_rg_s[4:0]),
      .z(inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd35),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd36)) inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg
      (
      .a(nl_inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg_a[34:0]),
      .s(nl_inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg_s[6:0]),
      .z(inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd35),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd36)) inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg
      (
      .a(nl_inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg_a[34:0]),
      .s(nl_inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg_s[6:0]),
      .z(inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd35),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd36)) inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg
      (
      .a(nl_inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg_a[34:0]),
      .s(nl_inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg_s[6:0]),
      .z(inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd35),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd36)) inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg
      (
      .a(nl_inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg_a[34:0]),
      .s(nl_inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_rg_s[6:0]),
      .z(inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd35),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd36)) inp_lookup_1_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg
      (
      .a(nl_inp_lookup_1_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg_a[34:0]),
      .s(nl_inp_lookup_1_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg_s[6:0]),
      .z(FpMantRNE_36U_11U_i_data_2_sva)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd35),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd36)) inp_lookup_2_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg
      (
      .a(nl_inp_lookup_2_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg_a[34:0]),
      .s(nl_inp_lookup_2_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg_s[6:0]),
      .z(FpMantRNE_36U_11U_i_data_3_sva)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd35),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd36)) inp_lookup_3_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg
      (
      .a(nl_inp_lookup_3_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg_a[34:0]),
      .s(nl_inp_lookup_3_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg_s[6:0]),
      .z(FpMantRNE_36U_11U_i_data_4_sva)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd35),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd36)) inp_lookup_4_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg
      (
      .a(nl_inp_lookup_4_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg_a[34:0]),
      .s(nl_inp_lookup_4_FpFractionToFloat_35U_6U_10U_if_shifted_frac_p1_lshift_rg_s[6:0]),
      .z(FpMantRNE_36U_11U_i_data_sva)
    );
  SDP_Y_INP_leading_sign_49_0 inp_lookup_1_leading_sign_49_0_rg (
      .mantissa(nl_inp_lookup_1_leading_sign_49_0_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_8)
    );
  SDP_Y_INP_leading_sign_49_0 inp_lookup_2_leading_sign_49_0_rg (
      .mantissa(nl_inp_lookup_2_leading_sign_49_0_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_9)
    );
  SDP_Y_INP_leading_sign_49_0 inp_lookup_3_leading_sign_49_0_rg (
      .mantissa(nl_inp_lookup_3_leading_sign_49_0_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_10)
    );
  SDP_Y_INP_leading_sign_49_0 inp_lookup_4_leading_sign_49_0_rg (
      .mantissa(nl_inp_lookup_4_leading_sign_49_0_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_11)
    );
  SDP_Y_INP_leading_sign_49_0 inp_lookup_1_leading_sign_49_0_1_rg (
      .mantissa(nl_inp_lookup_1_leading_sign_49_0_1_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_12)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) inp_lookup_1_FpNormalize_8U_49U_1_else_lshift_rg (
      .a(nl_inp_lookup_1_FpNormalize_8U_49U_1_else_lshift_rg_a[48:0]),
      .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_12),
      .z(inp_lookup_1_FpNormalize_8U_49U_1_else_lshift_itm)
    );
  SDP_Y_INP_leading_sign_49_0 inp_lookup_2_leading_sign_49_0_1_rg (
      .mantissa(nl_inp_lookup_2_leading_sign_49_0_1_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_13)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) inp_lookup_2_FpNormalize_8U_49U_1_else_lshift_rg (
      .a(nl_inp_lookup_2_FpNormalize_8U_49U_1_else_lshift_rg_a[48:0]),
      .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_13),
      .z(inp_lookup_2_FpNormalize_8U_49U_1_else_lshift_itm)
    );
  SDP_Y_INP_leading_sign_49_0 inp_lookup_3_leading_sign_49_0_1_rg (
      .mantissa(nl_inp_lookup_3_leading_sign_49_0_1_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_14)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) inp_lookup_3_FpNormalize_8U_49U_1_else_lshift_rg (
      .a(nl_inp_lookup_3_FpNormalize_8U_49U_1_else_lshift_rg_a[48:0]),
      .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_14),
      .z(inp_lookup_3_FpNormalize_8U_49U_1_else_lshift_itm)
    );
  SDP_Y_INP_leading_sign_49_0 inp_lookup_4_leading_sign_49_0_1_rg (
      .mantissa(nl_inp_lookup_4_leading_sign_49_0_1_rg_mantissa[48:0]),
      .rtn(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_15)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd49),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd49)) inp_lookup_4_FpNormalize_8U_49U_1_else_lshift_rg (
      .a(nl_inp_lookup_4_FpNormalize_8U_49U_1_else_lshift_rg_a[48:0]),
      .s(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_15),
      .z(inp_lookup_4_FpNormalize_8U_49U_1_else_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_r_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd24)) inp_lookup_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg
      (
      .a(nl_inp_lookup_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_a[23:0]),
      .s(nl_inp_lookup_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_s[3:0]),
      .z(inp_lookup_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_itm)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) inp_lookup_1_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_inp_lookup_1_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg_s[4:0]),
      .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_1_sva)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) inp_lookup_1_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_rg
      (
      .a(1'b1),
      .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_1_sva_2),
      .z(FpMantDecShiftRight_23U_8U_10U_least_mask_1_sva)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) inp_lookup_1_FpNormalize_6U_23U_1_else_lshift_rg (
      .a(nl_inp_lookup_1_FpNormalize_6U_23U_1_else_lshift_rg_a[22:0]),
      .s(libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_8),
      .z(inp_lookup_1_FpNormalize_6U_23U_1_else_lshift_itm)
    );
  SDP_Y_INP_leading_sign_23_0 inp_lookup_1_leading_sign_23_0_1_rg (
      .mantissa(nl_inp_lookup_1_leading_sign_23_0_1_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_8)
    );
  SDP_Y_INP_mgc_shift_r_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd24)) inp_lookup_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg
      (
      .a(nl_inp_lookup_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_a[23:0]),
      .s(nl_inp_lookup_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_s[3:0]),
      .z(inp_lookup_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_itm)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) inp_lookup_2_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_inp_lookup_2_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg_s[4:0]),
      .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_2_sva)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) inp_lookup_2_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_rg
      (
      .a(1'b1),
      .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_2_sva_2),
      .z(FpMantDecShiftRight_23U_8U_10U_least_mask_2_sva)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) inp_lookup_2_FpNormalize_6U_23U_1_else_lshift_rg (
      .a(nl_inp_lookup_2_FpNormalize_6U_23U_1_else_lshift_rg_a[22:0]),
      .s(libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_9),
      .z(inp_lookup_2_FpNormalize_6U_23U_1_else_lshift_itm)
    );
  SDP_Y_INP_leading_sign_23_0 inp_lookup_2_leading_sign_23_0_1_rg (
      .mantissa(nl_inp_lookup_2_leading_sign_23_0_1_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_9)
    );
  SDP_Y_INP_mgc_shift_r_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd24)) inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg
      (
      .a(nl_inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_a[23:0]),
      .s(nl_inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_s[3:0]),
      .z(inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_itm)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg_s[4:0]),
      .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_3_sva)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_rg
      (
      .a(1'b1),
      .s(reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_8_1_itm),
      .z(FpMantDecShiftRight_23U_8U_10U_least_mask_3_sva)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) inp_lookup_3_FpNormalize_6U_23U_1_else_lshift_rg (
      .a(nl_inp_lookup_3_FpNormalize_6U_23U_1_else_lshift_rg_a[22:0]),
      .s(libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_10),
      .z(inp_lookup_3_FpNormalize_6U_23U_1_else_lshift_itm)
    );
  SDP_Y_INP_leading_sign_23_0 inp_lookup_3_leading_sign_23_0_1_rg (
      .mantissa(nl_inp_lookup_3_leading_sign_23_0_1_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_10)
    );
  SDP_Y_INP_mgc_shift_r_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd24)) inp_lookup_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg
      (
      .a(nl_inp_lookup_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_a[23:0]),
      .s(nl_inp_lookup_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_s[3:0]),
      .z(inp_lookup_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_itm)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) inp_lookup_4_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg
      (
      .a(1'b1),
      .s(nl_inp_lookup_4_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg_s[4:0]),
      .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_sva)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) inp_lookup_4_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_rg
      (
      .a(1'b1),
      .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva_2),
      .z(FpMantDecShiftRight_23U_8U_10U_least_mask_sva)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) inp_lookup_4_FpNormalize_6U_23U_1_else_lshift_rg (
      .a(nl_inp_lookup_4_FpNormalize_6U_23U_1_else_lshift_rg_a[22:0]),
      .s(libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_11),
      .z(inp_lookup_4_FpNormalize_6U_23U_1_else_lshift_itm)
    );
  SDP_Y_INP_leading_sign_23_0 inp_lookup_4_leading_sign_23_0_1_rg (
      .mantissa(nl_inp_lookup_4_leading_sign_23_0_1_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_11)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) inp_lookup_1_FpNormalize_6U_23U_else_lshift_rg (
      .a(nl_inp_lookup_1_FpNormalize_6U_23U_else_lshift_rg_a[22:0]),
      .s(IntLeadZero_23U_leading_sign_23_0_rtn_1_sva_2),
      .z(inp_lookup_1_FpNormalize_6U_23U_else_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) inp_lookup_2_FpNormalize_6U_23U_else_lshift_rg (
      .a(nl_inp_lookup_2_FpNormalize_6U_23U_else_lshift_rg_a[22:0]),
      .s(IntLeadZero_23U_leading_sign_23_0_rtn_2_sva_2),
      .z(inp_lookup_2_FpNormalize_6U_23U_else_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) inp_lookup_3_FpNormalize_6U_23U_else_lshift_rg (
      .a(nl_inp_lookup_3_FpNormalize_6U_23U_else_lshift_rg_a[22:0]),
      .s(IntLeadZero_23U_leading_sign_23_0_rtn_3_sva_2),
      .z(inp_lookup_3_FpNormalize_6U_23U_else_lshift_itm)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) inp_lookup_4_FpNormalize_6U_23U_else_lshift_rg (
      .a(nl_inp_lookup_4_FpNormalize_6U_23U_else_lshift_rg_a[22:0]),
      .s(IntLeadZero_23U_leading_sign_23_0_rtn_sva_2),
      .z(inp_lookup_4_FpNormalize_6U_23U_else_lshift_itm)
    );
  SDP_Y_INP_leading_sign_10_0 inp_lookup_1_leading_sign_10_0_3_rg (
      .mantissa(nl_inp_lookup_1_leading_sign_10_0_3_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_16)
    );
  SDP_Y_INP_leading_sign_10_0 inp_lookup_2_leading_sign_10_0_3_rg (
      .mantissa(nl_inp_lookup_2_leading_sign_10_0_3_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_17)
    );
  SDP_Y_INP_leading_sign_10_0 inp_lookup_3_leading_sign_10_0_3_rg (
      .mantissa(nl_inp_lookup_3_leading_sign_10_0_3_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_18)
    );
  SDP_Y_INP_leading_sign_10_0 inp_lookup_4_leading_sign_10_0_3_rg (
      .mantissa(nl_inp_lookup_4_leading_sign_10_0_3_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_19)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) inp_lookup_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_inp_lookup_1_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_1_sva)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) inp_lookup_2_FpAdd_8U_23U_a_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_2_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_inp_lookup_2_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_2_sva)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) inp_lookup_3_FpAdd_8U_23U_a_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_3_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_inp_lookup_3_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_3_sva)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) inp_lookup_4_FpAdd_8U_23U_a_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_4_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_inp_lookup_4_FpAdd_8U_23U_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_a_int_mant_p1_sva)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) inp_lookup_1_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_1_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_inp_lookup_1_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_1_addend_larger_asn_19_mx0w1)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) inp_lookup_1_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_1_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_inp_lookup_1_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_1_a_int_mant_p1_1_sva)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) inp_lookup_2_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_2_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_inp_lookup_2_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_1_addend_larger_asn_13_mx0w1)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) inp_lookup_2_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_2_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_inp_lookup_2_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_1_a_int_mant_p1_2_sva)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) inp_lookup_3_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_3_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_inp_lookup_3_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_1_addend_larger_asn_7_mx0w1)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) inp_lookup_3_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_3_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_inp_lookup_3_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_1_a_int_mant_p1_3_sva)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) inp_lookup_4_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_4_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_inp_lookup_4_FpAdd_8U_23U_1_b_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_1_addend_larger_asn_1_mx0w1)
    );
  SDP_Y_INP_mgc_shift_bl_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd9),
  .width_z(32'sd49)) inp_lookup_4_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg (
      .a(nl_inp_lookup_4_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_a[23:0]),
      .s(nl_inp_lookup_4_FpAdd_8U_23U_1_a_int_mant_p1_lshift_rg_s[8:0]),
      .z(FpAdd_8U_23U_1_a_int_mant_p1_sva)
    );
  SDP_Y_INP_leading_sign_23_0 inp_lookup_1_leading_sign_23_0_rg (
      .mantissa(nl_inp_lookup_1_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_12)
    );
  SDP_Y_INP_leading_sign_23_0 inp_lookup_2_leading_sign_23_0_rg (
      .mantissa(nl_inp_lookup_2_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_13)
    );
  SDP_Y_INP_leading_sign_23_0 inp_lookup_3_leading_sign_23_0_rg (
      .mantissa(nl_inp_lookup_3_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_14)
    );
  SDP_Y_INP_leading_sign_23_0 inp_lookup_4_leading_sign_23_0_rg (
      .mantissa(nl_inp_lookup_4_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_15)
    );
  SDP_Y_INP_mgc_shift_br_v4 #(.width_a(32'sd65),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd81)) inp_lookup_1_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg
      (
      .a(nl_inp_lookup_1_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg_a[64:0]),
      .s(nl_inp_lookup_1_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg_s[4:0]),
      .z(IntSignedShiftRight_50U_5U_32U_mbits_fixed_1_sva)
    );
  SDP_Y_INP_mgc_shift_br_v4 #(.width_a(32'sd65),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd81)) inp_lookup_2_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg
      (
      .a(nl_inp_lookup_2_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg_a[64:0]),
      .s(nl_inp_lookup_2_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg_s[4:0]),
      .z(IntSignedShiftRight_50U_5U_32U_mbits_fixed_2_sva)
    );
  SDP_Y_INP_mgc_shift_br_v4 #(.width_a(32'sd65),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd81)) inp_lookup_3_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg
      (
      .a(nl_inp_lookup_3_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg_a[64:0]),
      .s(nl_inp_lookup_3_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg_s[4:0]),
      .z(IntSignedShiftRight_50U_5U_32U_mbits_fixed_3_sva)
    );
  SDP_Y_INP_mgc_shift_br_v4 #(.width_a(32'sd65),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd81)) inp_lookup_4_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg
      (
      .a(nl_inp_lookup_4_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg_a[64:0]),
      .s(nl_inp_lookup_4_IntSignedShiftRight_50U_5U_32U_mbits_fixed_rshift_rg_s[4:0]),
      .z(IntSignedShiftRight_50U_5U_32U_mbits_fixed_sva)
    );
  SDP_Y_INP_leading_sign_10_0 inp_lookup_1_leading_sign_10_0_2_rg (
      .mantissa(nl_inp_lookup_1_leading_sign_10_0_2_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_20)
    );
  SDP_Y_INP_leading_sign_10_0 inp_lookup_2_leading_sign_10_0_2_rg (
      .mantissa(nl_inp_lookup_2_leading_sign_10_0_2_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_21)
    );
  SDP_Y_INP_leading_sign_10_0 inp_lookup_3_leading_sign_10_0_2_rg (
      .mantissa(nl_inp_lookup_3_leading_sign_10_0_2_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_22)
    );
  SDP_Y_INP_leading_sign_10_0 inp_lookup_4_leading_sign_10_0_2_rg (
      .mantissa(nl_inp_lookup_4_leading_sign_10_0_2_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_23)
    );
  SDP_Y_INP_leading_sign_10_0 inp_lookup_1_leading_sign_10_0_rg (
      .mantissa(nl_inp_lookup_1_leading_sign_10_0_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_24)
    );
  SDP_Y_INP_leading_sign_10_0 inp_lookup_2_leading_sign_10_0_rg (
      .mantissa(nl_inp_lookup_2_leading_sign_10_0_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_25)
    );
  SDP_Y_INP_leading_sign_10_0 inp_lookup_3_leading_sign_10_0_rg (
      .mantissa(nl_inp_lookup_3_leading_sign_10_0_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_26)
    );
  SDP_Y_INP_leading_sign_10_0 inp_lookup_4_leading_sign_10_0_rg (
      .mantissa(nl_inp_lookup_4_leading_sign_10_0_rg_mantissa[9:0]),
      .rtn(libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_27)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd9),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd10)) inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg
      (
      .a(nl_inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg_a[8:0]),
      .s(nl_inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg_s[4:0]),
      .z(z_out_16)
    );
  SDP_Y_INP_mgc_shift_l_v4 #(.width_a(32'sd9),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd10)) inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg
      (
      .a(nl_inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg_a[8:0]),
      .s(nl_inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_rg_s[4:0]),
      .z(z_out_17)
    );
  NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_in_rsci NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_in_rsci_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_inp_in_rsc_z(chn_inp_in_rsc_z),
      .chn_inp_in_rsc_vz(chn_inp_in_rsc_vz),
      .chn_inp_in_rsc_lz(chn_inp_in_rsc_lz),
      .chn_inp_in_rsci_oswt(chn_inp_in_rsci_oswt),
      .core_wen(core_wen),
      .chn_inp_in_rsci_iswt0(chn_inp_in_rsci_iswt0),
      .chn_inp_in_rsci_bawt(chn_inp_in_rsci_bawt),
      .chn_inp_in_rsci_wen_comp(chn_inp_in_rsci_wen_comp),
      .chn_inp_in_rsci_ld_core_psct(chn_inp_in_rsci_ld_core_psct),
      .chn_inp_in_rsci_d_mxwt(chn_inp_in_rsci_d_mxwt),
      .core_wten(core_wten)
    );
  NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_out_rsci NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_out_rsci_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_inp_out_rsc_z(chn_inp_out_rsc_z),
      .chn_inp_out_rsc_vz(chn_inp_out_rsc_vz),
      .chn_inp_out_rsc_lz(chn_inp_out_rsc_lz),
      .chn_inp_out_rsci_oswt(chn_inp_out_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_inp_out_rsci_iswt0(chn_inp_out_rsci_iswt0),
      .chn_inp_out_rsci_bawt(chn_inp_out_rsci_bawt),
      .chn_inp_out_rsci_wen_comp(chn_inp_out_rsci_wen_comp),
      .chn_inp_out_rsci_ld_core_psct(reg_chn_inp_out_rsci_ld_core_psct_cse),
      .chn_inp_out_rsci_d(nl_NV_NVDLA_SDP_CORE_Y_inp_core_chn_inp_out_rsci_inst_chn_inp_out_rsci_d[127:0])
    );
  NV_NVDLA_SDP_CORE_Y_inp_core_staller NV_NVDLA_SDP_CORE_Y_inp_core_staller_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .chn_inp_in_rsci_wen_comp(chn_inp_in_rsci_wen_comp),
      .core_wten(core_wten),
      .chn_inp_out_rsci_wen_comp(chn_inp_out_rsci_wen_comp)
    );
  NV_NVDLA_SDP_CORE_Y_inp_core_core_fsm NV_NVDLA_SDP_CORE_Y_inp_core_core_fsm_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign and_44 = main_stage_v_7 & (cfg_precision_1_sva_st_84==2'b10) & (~ inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs)
      & inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2
      & (~ inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2)
      & (chn_inp_in_crt_sva_7_739_736_1[0]) & or_11_cse;
  assign shift_0_prb = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ reg_FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_8_3_0_1_itm)
      , (FpAdd_6U_10U_1_qr_2_lpi_1_dfm_5[0])}) + 5'b1)), and_44);
// assert(shift > 0) - ../include/nvdla_float.h: line 286
// PSL inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln286_assert_shift_gt_0 : assert { shift_0_prb } @rose(nvdla_core_clk);
  assign and_51 = and_dcpl_21 & (~ (cfg_precision_1_sva_st_84[0])) & inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2
      & (~(inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
      | inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2))
      & or_11_cse;
  assign shift_0_prb_1 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ reg_FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_8_3_0_1_itm)
      , (FpAdd_6U_10U_1_qr_3_lpi_1_dfm_5[0])}) + 5'b1)), and_51);
// assert(shift > 0) - ../include/nvdla_float.h: line 286
// PSL inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln286_assert_shift_gt_0 : assert { shift_0_prb_1 } @rose(nvdla_core_clk);
  assign and_58 = main_stage_v_7 & (cfg_precision_1_sva_st_84==2'b10) & (chn_inp_in_crt_sva_7_739_736_1[2])
      & inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2
      & (~(inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
      | inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2))
      & or_11_cse;
  assign shift_0_prb_2 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ reg_FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_8_3_0_1_itm)
      , (FpAdd_6U_10U_1_qr_4_lpi_1_dfm_5[0])}) + 5'b1)), and_58);
// assert(shift > 0) - ../include/nvdla_float.h: line 286
// PSL inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln286_assert_shift_gt_0 : assert { shift_0_prb_2 } @rose(nvdla_core_clk);
  assign and_65 = main_stage_v_7 & (cfg_precision_1_sva_st_84==2'b10) & inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2
      & (~ inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs)
      & (chn_inp_in_crt_sva_7_739_736_1[3]) & (~ inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2)
      & or_11_cse;
  assign shift_0_prb_3 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ reg_FpMul_6U_10U_1_o_expo_lpi_1_dfm_8_3_0_1_itm)
      , (FpAdd_6U_10U_1_qr_lpi_1_dfm_5[0])}) + 5'b1)), and_65);
// assert(shift > 0) - ../include/nvdla_float.h: line 286
// PSL inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln286_assert_shift_gt_0 : assert { shift_0_prb_3 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb = inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iMantWidth >= oMantWidth) - ../include/nvdla_float.h: line 669
// PSL inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln669_assert_iMantWidth_ge_oMantWidth : assert { iMantWidth_oMantWidth_prb } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb = inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iExpoWidth >= oExpoWidth) - ../include/nvdla_float.h: line 670
// PSL inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_1 = inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_1 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_1 = inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth : assert { iMantWidth_oMantWidth_prb_1 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_2 = inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_2 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_3 = inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_3 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_2 = inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_2 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_3 = inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_3 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_4 = inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2 : assert { iExpoWidth_oExpoWidth_prb_4 } @rose(nvdla_core_clk);
  assign or_4171 = (and_dcpl_42 & and_dcpl_38 & (fsm_output[1])) | (and_dcpl_42 &
      (chn_inp_in_rsci_d_mxwt[736]) & chn_inp_out_rsci_bawt & reg_chn_inp_out_rsci_ld_core_psct_cse);
  assign oWidth_iWidth_prb = MUX1HOT_s_1_1_2(1'b1, or_4171);
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth : assert { oWidth_iWidth_prb } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_5 = inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_3 : assert { iExpoWidth_oExpoWidth_prb_5 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_6 = inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_4 : assert { iExpoWidth_oExpoWidth_prb_6 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_4 = inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_4 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_5 = inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_2 : assert { iMantWidth_oMantWidth_prb_5 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_7 = inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_7 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_6 = inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_6 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_7 = inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_7 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_8 = inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5 : assert { iExpoWidth_oExpoWidth_prb_8 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_8 = inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iMantWidth >= oMantWidth) - ../include/nvdla_float.h: line 669
// PSL inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln669_assert_iMantWidth_ge_oMantWidth : assert { iMantWidth_oMantWidth_prb_8 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_9 = inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iExpoWidth >= oExpoWidth) - ../include/nvdla_float.h: line 670
// PSL inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_9 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_10 = inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_10 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_9 = inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth : assert { iMantWidth_oMantWidth_prb_9 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_11 = inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_11 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_12 = inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_12 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_10 = inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_10 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_11 = inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_11 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_13 = inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2 : assert { iExpoWidth_oExpoWidth_prb_13 } @rose(nvdla_core_clk);
  assign or_4174 = (and_dcpl_42 & and_dcpl_49 & (fsm_output[1])) | (and_dcpl_42 &
      (chn_inp_in_rsci_d_mxwt[737]) & chn_inp_out_rsci_bawt & reg_chn_inp_out_rsci_ld_core_psct_cse);
  assign oWidth_iWidth_prb_1 = MUX1HOT_s_1_1_2(1'b1, or_4174);
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth : assert { oWidth_iWidth_prb_1 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_14 = inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_3 : assert { iExpoWidth_oExpoWidth_prb_14 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_15 = inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_4 : assert { iExpoWidth_oExpoWidth_prb_15 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_12 = inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_12 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_13 = inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_2 : assert { iMantWidth_oMantWidth_prb_13 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_16 = inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_16 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_14 = inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_14 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_15 = inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_15 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_17 = inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5 : assert { iExpoWidth_oExpoWidth_prb_17 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_16 = inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iMantWidth >= oMantWidth) - ../include/nvdla_float.h: line 669
// PSL inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln669_assert_iMantWidth_ge_oMantWidth : assert { iMantWidth_oMantWidth_prb_16 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_18 = inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iExpoWidth >= oExpoWidth) - ../include/nvdla_float.h: line 670
// PSL inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_18 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_19 = inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_19 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_17 = inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth : assert { iMantWidth_oMantWidth_prb_17 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_20 = inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_20 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_21 = inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_21 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_18 = inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_18 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_19 = inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_19 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_22 = inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2 : assert { iExpoWidth_oExpoWidth_prb_22 } @rose(nvdla_core_clk);
  assign or_4177 = (and_dcpl_42 & and_dcpl_57 & (fsm_output[1])) | (and_dcpl_42 &
      (chn_inp_in_rsci_d_mxwt[738]) & chn_inp_out_rsci_bawt & reg_chn_inp_out_rsci_ld_core_psct_cse);
  assign oWidth_iWidth_prb_2 = MUX1HOT_s_1_1_2(1'b1, or_4177);
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth : assert { oWidth_iWidth_prb_2 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_23 = inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_3 : assert { iExpoWidth_oExpoWidth_prb_23 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_24 = inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_4 : assert { iExpoWidth_oExpoWidth_prb_24 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_20 = inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_20 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_21 = inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_2 : assert { iMantWidth_oMantWidth_prb_21 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_25 = inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_25 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_22 = inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_22 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_23 = inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_23 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_26 = inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5 : assert { iExpoWidth_oExpoWidth_prb_26 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_24 = inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iMantWidth >= oMantWidth) - ../include/nvdla_float.h: line 669
// PSL inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln669_assert_iMantWidth_ge_oMantWidth : assert { iMantWidth_oMantWidth_prb_24 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_27 = inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iExpoWidth >= oExpoWidth) - ../include/nvdla_float.h: line 670
// PSL inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_27 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_28 = inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_28 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_25 = inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth : assert { iMantWidth_oMantWidth_prb_25 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_29 = inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_29 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_30 = inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb_30 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_26 = inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_26 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_27 = inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth : assert { iMantWidth_oMantWidth_prb_27 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_31 = inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2 : assert { iExpoWidth_oExpoWidth_prb_31 } @rose(nvdla_core_clk);
  assign or_4180 = (and_dcpl_42 & and_dcpl_65 & (fsm_output[1])) | (and_dcpl_42 &
      (chn_inp_in_rsci_d_mxwt[739]) & chn_inp_out_rsci_bawt & reg_chn_inp_out_rsci_ld_core_psct_cse);
  assign oWidth_iWidth_prb_3 = MUX1HOT_s_1_1_2(1'b1, or_4180);
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth : assert { oWidth_iWidth_prb_3 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_32 = inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_3 : assert { iExpoWidth_oExpoWidth_prb_32 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_33 = inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_4 : assert { iExpoWidth_oExpoWidth_prb_33 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_28 = inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_28 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_29 = inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iMantWidth > oMantWidth) - ../include/nvdla_float.h: line 334
// PSL inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln334_assert_iMantWidth_gt_oMantWidth_2 : assert { iMantWidth_oMantWidth_prb_29 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_34 = inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 556
// PSL inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln556_assert_iExpoWidth_le_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_34 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_30 = inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 557
// PSL inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln557_assert_iMantWidth_le_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_30 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_31 = inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iMantWidth <= oMantWidth) - ../include/nvdla_float.h: line 508
// PSL inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln508_assert_iMantWidth_le_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_31 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_35 = inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1;
// assert(iExpoWidth <= oExpoWidth) - ../include/nvdla_float.h: line 433
// PSL inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5 : assert { iExpoWidth_oExpoWidth_prb_35 } @rose(nvdla_core_clk);
  assign chn_inp_out_and_cse = core_wen & (~ or_dcpl_4);
  assign or_5836_tmp = inp_lookup_asn_106 | inp_lookup_and_8_m1c;
  assign and_3545_tmp = ((~ IsInf_6U_23U_land_1_lpi_1_dfm_mx0w0) | IsNaN_6U_23U_land_1_lpi_1_dfm_mx2)
      & inp_lookup_and_10_m1c;
  assign or_5838_tmp = inp_lookup_asn_122 | inp_lookup_and_28_m1c;
  assign and_3546_tmp = ((~ IsInf_6U_23U_land_2_lpi_1_dfm_mx0w0) | IsNaN_6U_23U_land_2_lpi_1_dfm_mx2)
      & inp_lookup_and_30_m1c;
  assign or_5840_tmp = inp_lookup_asn_114 | inp_lookup_and_48_m1c;
  assign and_3547_tmp = ((~ IsInf_6U_23U_land_3_lpi_1_dfm_mx0w0) | IsNaN_6U_23U_land_3_lpi_1_dfm_mx1)
      & inp_lookup_and_50_m1c;
  assign or_5842_tmp = inp_lookup_asn_98 | inp_lookup_and_68_m1c;
  assign and_3548_tmp = ((~ IsInf_6U_23U_land_lpi_1_dfm_mx0w0) | IsNaN_6U_23U_land_lpi_1_dfm_mx1)
      & inp_lookup_and_70_m1c;
  assign mux_78_nl = MUX_s_1_2_2(nand_694_cse, nand_602_cse_1, or_11_cse);
  assign IsNaN_8U_23U_aelse_and_cse = core_wen & (~ and_dcpl_78) & (~ (mux_78_nl));
  assign FpAdd_8U_23U_is_a_greater_oelse_and_cse = core_wen & (and_dcpl_38 | and_dcpl_105)
      & (~ mux_93_cse);
  assign or_11_cse = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt;
  assign IntLeadZero_35U_1_leading_sign_35_0_rtn_and_4_cse = core_wen & (and_dcpl_106
      | and_dcpl_141) & (~ mux_81_itm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_12_cse = core_wen & (and_dcpl_144
      | and_dcpl_145) & mux_tmp_6;
  assign FpFractionToFloat_35U_6U_10U_1_if_else_else_and_cse = core_wen & (~ and_dcpl_78)
      & (~ mux_81_itm);
  assign cfg_precision_and_cse = core_wen & (~ and_dcpl_78) & mux_tmp_6;
  assign FpAdd_8U_23U_is_a_greater_oelse_FpAdd_8U_23U_is_a_greater_oelse_or_19_cse
      = and_dcpl_49 | and_dcpl_176;
  assign FpAdd_8U_23U_is_a_greater_oelse_and_1_cse = core_wen & FpAdd_8U_23U_is_a_greater_oelse_FpAdd_8U_23U_is_a_greater_oelse_or_19_cse
      & (~ mux_93_cse);
  assign IntLeadZero_35U_1_leading_sign_35_0_rtn_and_5_cse = core_wen & (and_dcpl_177
      | and_dcpl_212) & (~ mux_87_itm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_15_cse = core_wen & (and_dcpl_214
      | and_dcpl_215) & mux_tmp_6;
  assign FpFractionToFloat_35U_6U_10U_1_if_else_else_and_1_cse = core_wen & (~ and_dcpl_78)
      & (~ mux_87_itm);
  assign mux_93_cse = MUX_s_1_2_2(or_tmp_8, or_tmp_6, or_11_cse);
  assign FpAdd_8U_23U_is_a_greater_oelse_and_2_cse = core_wen & (and_dcpl_57 | and_dcpl_246)
      & (~ mux_93_cse);
  assign or_82_cse = (inp_lookup_3_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_3!=35'b00000000000000000000000000000000000);
  assign or_79_cse = (chn_inp_in_rsci_d_mxwt[232:198]!=35'b00000000000000000000000000000000000);
  assign IntLeadZero_35U_1_leading_sign_35_0_rtn_and_6_cse = core_wen & (and_dcpl_247
      | and_dcpl_282) & (~ mux_95_itm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_18_cse = core_wen & (and_dcpl_284
      | and_dcpl_285) & mux_tmp_6;
  assign FpFractionToFloat_35U_6U_10U_1_if_else_else_and_2_cse = core_wen & (~ and_dcpl_78)
      & (~ mux_95_itm);
  assign FpAdd_8U_23U_is_a_greater_oelse_FpAdd_8U_23U_is_a_greater_oelse_or_17_cse
      = and_dcpl_65 | and_dcpl_316;
  assign FpAdd_8U_23U_is_a_greater_oelse_and_3_cse = core_wen & FpAdd_8U_23U_is_a_greater_oelse_FpAdd_8U_23U_is_a_greater_oelse_or_17_cse
      & (~ mux_93_cse);
  assign nor_1713_cse = ~((inp_lookup_4_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_3!=35'b00000000000000000000000000000000000));
  assign IntLeadZero_35U_1_leading_sign_35_0_rtn_and_7_cse = core_wen & (and_dcpl_317
      | and_dcpl_352) & (~ mux_100_itm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_21_cse = core_wen & (and_dcpl_354
      | and_dcpl_355) & mux_tmp_6;
  assign FpFractionToFloat_35U_6U_10U_1_if_else_else_and_3_cse = core_wen & (~ and_dcpl_78)
      & (~ mux_100_itm);
  assign nand_772_cse = ~(main_stage_v_2 & (chn_inp_in_crt_sva_2_739_736_1[0]) &
      (cfg_precision_1_sva_st_91==2'b10));
  assign mux_108_nl = MUX_s_1_2_2(nand_772_cse, nand_tmp_3, or_11_cse);
  assign FpAdd_8U_23U_addend_larger_and_cse = core_wen & ((or_11_cse & FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_5)
      | and_dcpl_390) & (~ (mux_108_nl));
  assign mux_110_nl = MUX_s_1_2_2(nand_772_cse, nand_694_cse, or_11_cse);
  assign FpAdd_8U_23U_is_addition_and_cse = core_wen & (~ and_dcpl_78) & (~ (mux_110_nl));
  assign and_861_rgt = or_11_cse & (~ inp_lookup_1_FpMantRNE_36U_11U_else_and_tmp);
  assign and_3393_cse = (chn_inp_in_crt_sva_2_739_736_1[0]) & main_stage_v_2 & (cfg_precision_1_sva_st_91==2'b10);
  assign FpFractionToFloat_35U_6U_10U_is_zero_FpFractionToFloat_35U_6U_10U_is_zero_or_3_cse
      = and_dcpl_393 | and_dcpl_394;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_cse = core_wen & FpFractionToFloat_35U_6U_10U_is_zero_FpFractionToFloat_35U_6U_10U_is_zero_or_3_cse
      & (~ mux_115_itm);
  assign mux_116_nl = MUX_s_1_2_2(or_5800_cse, or_tmp_21, or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_17_cse = core_wen & (~ and_dcpl_78)
      & (~ (mux_116_nl));
  assign and_3369_nl = nor_1380_cse & (~(((~ inp_lookup_1_FpMul_6U_10U_2_else_2_if_acc_itm_6)
      | or_5873_cse) & or_178_cse));
  assign nor_1700_nl = ~((~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[0])
      | (cfg_precision_1_sva_st_91[0]) | (~((cfg_precision_1_sva_st_91[1]) & (IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_14
      | nor_44_cse))));
  assign mux_119_nl = MUX_s_1_2_2((nor_1700_nl), (and_3369_nl), or_11_cse);
  assign FpFractionToFloat_35U_6U_10U_1_o_mant_and_12_cse = core_wen & (~ and_dcpl_78)
      & (mux_119_nl);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_asn_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_conc_40_cgspt_7_mux_nl
      = MUX_v_8_2_2((chn_inp_in_crt_sva_1_739_395_1[115:108]), (chn_inp_in_crt_sva_1_739_395_1[243:236]),
      and_dcpl_390);
  assign mux_1866_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_2_739_736_1[0]), (chn_inp_in_crt_sva_1_739_395_1[341]),
      or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_mux1h_1_itm = MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_8,
      ({2'b0 , (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_asn_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_conc_40_cgspt_7_mux_nl)}),
      mux_1866_nl);
  assign or_5873_cse = IsZero_6U_10U_6_IsZero_6U_10U_6_nor_tmp | inp_lookup_1_FpMul_6U_10U_2_oelse_1_acc_itm_7
      | IsZero_6U_10U_7_IsZero_6U_10U_7_and_itm_2;
  assign nor_1896_cse = ~(chn_inp_out_rsci_bawt | (~ reg_chn_inp_out_rsci_ld_core_psct_cse));
  assign or_5882_cse = (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_8!=10'b0000000000);
  assign cfg_precision_and_4_cse = core_wen & (~ and_dcpl_78) & mux_tmp_50;
  assign mux_129_nl = MUX_s_1_2_2(nand_358_cse, nand_tmp_5, or_11_cse);
  assign FpAdd_8U_23U_addend_larger_and_1_cse = core_wen & ((or_11_cse & FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_5)
      | and_dcpl_398) & (~ (mux_129_nl));
  assign mux_133_nl = MUX_s_1_2_2(nand_358_cse, or_tmp_213, or_11_cse);
  assign FpAdd_8U_23U_is_addition_and_2_cse = core_wen & (~ and_dcpl_78) & (~ (mux_133_nl));
  assign and_869_rgt = or_11_cse & (~ inp_lookup_2_FpMantRNE_36U_11U_else_and_tmp);
  assign and_3391_cse = (chn_inp_in_crt_sva_2_739_736_1[1]) & main_stage_v_2 & (cfg_precision_1_sva_st_91==2'b10);
  assign FpFractionToFloat_35U_6U_10U_is_zero_FpFractionToFloat_35U_6U_10U_is_zero_or_2_cse
      = and_dcpl_401 | and_dcpl_402;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_18_cse = core_wen & FpFractionToFloat_35U_6U_10U_is_zero_FpFractionToFloat_35U_6U_10U_is_zero_or_2_cse
      & (~ mux_115_itm);
  assign mux_139_nl = MUX_s_1_2_2(or_tmp_234, or_tmp_52, or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_19_cse = core_wen & (~ and_dcpl_78)
      & (~ (mux_139_nl));
  assign nor_1683_nl = ~(inp_lookup_2_FpMul_6U_10U_2_else_2_if_acc_itm_6 | (~ or_tmp_241));
  assign mux_141_nl = MUX_s_1_2_2((nor_1683_nl), or_tmp_241, or_5890_cse);
  assign nor_1682_nl = ~((~ main_stage_v_1) | (chn_inp_in_crt_sva_1_739_395_1[342])
      | (cfg_precision_1_sva_st_90!=2'b10) | (mux_141_nl));
  assign nor_1684_nl = ~((~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[1])
      | (cfg_precision_1_sva_st_91[0]) | (~((cfg_precision_1_sva_st_91[1]) & (IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_14
      | nor_268_cse))));
  assign mux_142_nl = MUX_s_1_2_2((nor_1684_nl), (nor_1682_nl), or_11_cse);
  assign FpFractionToFloat_35U_6U_10U_1_o_mant_and_13_cse = core_wen & (~ and_dcpl_78)
      & (mux_142_nl);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_asn_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_conc_41_cgspt_7_mux_nl
      = MUX_v_8_2_2((chn_inp_in_crt_sva_1_739_395_1[147:140]), (chn_inp_in_crt_sva_1_739_395_1[275:268]),
      and_dcpl_398);
  assign mux_1867_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_2_739_736_1[1]), (chn_inp_in_crt_sva_1_739_395_1[342]),
      or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_mux1h_3_itm = MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_8,
      ({2'b0 , (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_asn_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_conc_41_cgspt_7_mux_nl)}),
      mux_1867_nl);
  assign or_5889_cse = (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_8!=10'b0000000000);
  assign or_5890_cse = inp_lookup_2_FpMul_6U_10U_2_oelse_1_acc_itm_7 | IsZero_6U_10U_7_IsZero_6U_10U_7_and_1_itm_2
      | IsZero_6U_10U_6_IsZero_6U_10U_6_nor_1_tmp;
  assign or_5896_cse = inp_lookup_2_FpMul_6U_10U_2_oelse_1_acc_itm_7 | IsZero_6U_10U_7_IsZero_6U_10U_7_and_1_itm_2
      | IsZero_6U_10U_6_IsZero_6U_10U_6_nor_1_tmp | (~ inp_lookup_2_FpMul_6U_10U_2_else_2_if_acc_itm_6);
  assign and_4145_cse = or_5889_cse & FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_6_1_1
      & FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_6_0_1 & (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_9==4'b1111);
  assign mux_151_nl = MUX_s_1_2_2(or_tmp_277, nand_tmp_8, or_11_cse);
  assign FpAdd_8U_23U_addend_larger_and_2_cse = core_wen & ((or_11_cse & FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_5)
      | and_dcpl_406) & (~ (mux_151_nl));
  assign mux_155_nl = MUX_s_1_2_2(or_tmp_277, nand_693_cse, or_11_cse);
  assign FpAdd_8U_23U_is_addition_and_4_cse = core_wen & (~ and_dcpl_78) & (~ (mux_155_nl));
  assign and_877_rgt = or_11_cse & (~ inp_lookup_3_FpMantRNE_36U_11U_else_and_tmp);
  assign and_3401_cse = (chn_inp_in_crt_sva_2_739_736_1[2]) & main_stage_v_2 & (cfg_precision_1_sva_st_91==2'b10);
  assign and_3389_cse = (chn_inp_in_crt_sva_1_739_395_1[343]) & main_stage_v_1 &
      (cfg_precision_1_sva_st_90==2'b10);
  assign FpFractionToFloat_35U_6U_10U_is_zero_FpFractionToFloat_35U_6U_10U_is_zero_or_1_cse
      = and_dcpl_409 | and_dcpl_410;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_20_cse = core_wen & FpFractionToFloat_35U_6U_10U_is_zero_FpFractionToFloat_35U_6U_10U_is_zero_or_1_cse
      & (~ mux_115_itm);
  assign mux_161_nl = MUX_s_1_2_2(or_tmp_306, or_tmp_85, or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_21_cse = core_wen & (~ and_dcpl_78)
      & (~ (mux_161_nl));
  assign and_3364_nl = nor_1354_cse & (~(((~ inp_lookup_3_FpMul_6U_10U_2_else_2_if_acc_itm_6_1)
      | FpMul_6U_10U_2_if_2_FpMul_6U_10U_2_if_2_or_5_tmp) & nand_616_cse));
  assign nor_1662_nl = ~((~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[2])
      | (cfg_precision_1_sva_st_91[0]) | (~((cfg_precision_1_sva_st_91[1]) & (IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_14
      | nor_67_cse))));
  assign mux_164_nl = MUX_s_1_2_2((nor_1662_nl), (and_3364_nl), or_11_cse);
  assign FpFractionToFloat_35U_6U_10U_1_o_mant_and_14_cse = core_wen & (~ and_dcpl_78)
      & (mux_164_nl);
  assign nor_1661_nl = ~((cfg_precision_1_sva_st_90!=2'b10) | (chn_inp_in_crt_sva_1_739_395_1[343])
      | (~(main_stage_v_1 & (nor_301_cse | (inp_lookup_3_IsNaN_6U_10U_7_aif_IsNaN_6U_10U_7_aelse_IsNaN_6U_10U_7_aelse_or_tmp
      & FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_6_1_1 & FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_6_0_1
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_3_lpi_1_dfm_9==4'b1111) & nand_616_cse)))));
  assign and_3363_nl = (~((~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[2])
      | (cfg_precision_1_sva_st_91!=2'b10))) & (~(((~ IsNaN_6U_10U_7_land_3_lpi_1_dfm_5)
      | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_14) & (FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_3
      | (~ inp_lookup_3_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs))));
  assign mux_165_nl = MUX_s_1_2_2((and_3363_nl), (nor_1661_nl), or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_and_cse = core_wen & (~ and_dcpl_78)
      & (mux_165_nl);
  assign mux_170_nl = MUX_s_1_2_2(nand_701_cse, nand_tmp_12, or_11_cse);
  assign FpAdd_8U_23U_addend_larger_and_3_cse = core_wen & ((or_11_cse & FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2)
      | and_dcpl_412) & (~ (mux_170_nl));
  assign mux_174_nl = MUX_s_1_2_2(nand_701_cse, or_tmp_347, or_11_cse);
  assign FpAdd_8U_23U_is_addition_and_6_cse = core_wen & (~ and_dcpl_78) & (~ (mux_174_nl));
  assign or_356_cse = (inp_lookup_4_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_4!=35'b00000000000000000000000000000000000);
  assign and_883_rgt = or_11_cse & (~ inp_lookup_4_FpMantRNE_36U_11U_else_and_tmp);
  assign FpFractionToFloat_35U_6U_10U_is_zero_FpFractionToFloat_35U_6U_10U_is_zero_or_cse
      = and_dcpl_415 | and_dcpl_416;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_22_cse = core_wen & FpFractionToFloat_35U_6U_10U_is_zero_FpFractionToFloat_35U_6U_10U_is_zero_or_cse
      & (~ mux_115_itm);
  assign mux_179_nl = MUX_s_1_2_2(or_5809_cse, or_tmp_114, or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_24_cse = core_wen & (~ and_dcpl_78)
      & (~ (mux_179_nl));
  assign nor_1650_nl = ~((chn_inp_in_crt_sva_1_739_395_1[344]) | (~ main_stage_v_1)
      | (cfg_precision_1_sva_st_90!=2'b10));
  assign and_3388_nl = (IntLeadZero_35U_1_leading_sign_35_0_rtn_sva_2[5]) & inp_lookup_4_FpMantRNE_36U_11U_1_else_and_svs_2
      & FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2 & (~ IsNaN_6U_10U_6_nor_3_tmp)
      & (FpFractionToFloat_35U_6U_10U_1_mux_42_tmp==5'b11111) & (~ (chn_inp_in_crt_sva_1_739_395_1[344]))
      & main_stage_v_1 & (cfg_precision_1_sva_st_90==2'b10);
  assign mux_181_nl = MUX_s_1_2_2((and_3388_nl), (nor_1650_nl), nor_29_cse);
  assign nor_1652_nl = ~((~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[3])
      | (cfg_precision_1_sva_st_91[0]) | (~((cfg_precision_1_sva_st_91[1]) & (IsNaN_6U_10U_2_land_lpi_1_dfm_st_14
      | (~(FpMul_6U_10U_2_lor_1_lpi_1_dfm_st_3 | (~ inp_lookup_4_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs)))))));
  assign mux_182_nl = MUX_s_1_2_2((nor_1652_nl), (mux_181_nl), or_11_cse);
  assign FpFractionToFloat_35U_6U_10U_1_o_mant_and_15_cse = core_wen & (~ and_dcpl_78)
      & (mux_182_nl);
  assign and_3361_cse_1 = or_5904_cse & FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_6_1_1
      & FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_6_0_1 & (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_9==4'b1111);
  assign nor_29_cse = ~(FpMul_6U_10U_2_if_2_FpMul_6U_10U_2_if_2_or_7_tmp | (~ inp_lookup_4_FpMul_6U_10U_2_else_2_if_acc_itm_6));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_asn_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_conc_42_cgspt_7_mux_nl
      = MUX_v_8_2_2((chn_inp_in_crt_sva_1_739_395_1[211:204]), (chn_inp_in_crt_sva_1_739_395_1[339:332]),
      and_dcpl_412);
  assign mux_1868_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_2_739_736_1[3]), (chn_inp_in_crt_sva_1_739_395_1[344]),
      or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_mux1h_6_itm = MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_8,
      ({2'b0 , (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_asn_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_conc_42_cgspt_7_mux_nl)}),
      mux_1868_nl);
  assign or_6160_cse = (FpFractionToFloat_35U_6U_10U_1_o_mant_lpi_1_dfm_6!=10'b0000000000);
  assign or_5904_cse = (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_8!=10'b0000000000);
  assign mux_190_nl = MUX_s_1_2_2(main_stage_v_3, main_stage_v_2, or_11_cse);
  assign and_3624_cse = core_wen & (~ and_dcpl_78) & (mux_190_nl);
  assign nand_602_cse_1 = ~((chn_inp_in_rsci_d_mxwt[736]) & chn_inp_in_rsci_bawt
      & (cfg_precision_rsci_d==2'b10));
  assign nand_694_cse = ~(main_stage_v_1 & (chn_inp_in_crt_sva_1_739_395_1[341])
      & (cfg_precision_1_sva_st_90==2'b10));
  assign and_3463_cse = (fsm_output[1]) & core_wen;
  assign or_4340_cse = (~ (chn_inp_in_crt_sva_3_739_736_1[0])) | (cfg_precision_1_sva_st_80!=2'b10);
  assign nor_1961_cse = ~((~ (chn_inp_in_crt_sva_2_739_736_1[0])) | (cfg_precision_1_sva_st_91!=2'b10));
  assign or_6241_cse = (~ (chn_inp_in_crt_sva_1_739_395_1[341])) | (cfg_precision_1_sva_st_90[0]);
  assign nor_1978_cse = ~((cfg_precision_1_sva_st_91[1]) | (~ (fsm_output[0])));
  assign and_899_rgt = and_dcpl_428 & (~ IsNaN_6U_10U_7_land_1_lpi_1_dfm_5) & or_11_cse;
  assign and_901_rgt = and_dcpl_428 & IsNaN_6U_10U_7_land_1_lpi_1_dfm_5 & or_11_cse;
  assign and_903_rgt = and_dcpl_433 & or_11_cse;
  assign FpAdd_8U_23U_o_expo_and_cse = core_wen & (~ (fsm_output[0]));
  assign and_907_rgt = and_dcpl_437 & or_11_cse & (~ (z_out[49]));
  assign and_912_rgt = nand_772_cse & (cfg_precision_1_sva_st_80==2'b10) & (chn_inp_in_crt_sva_3_739_736_1[0])
      & main_stage_v_3 & or_11_cse;
  assign and_915_rgt = and_dcpl_437 & (z_out[49]) & inp_lookup_1_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1
      & or_11_cse;
  assign and_918_rgt = and_dcpl_437 & (z_out[49]) & (~ inp_lookup_1_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1)
      & or_11_cse;
  assign and_131_cse = main_stage_v_3 & (chn_inp_in_crt_sva_3_739_736_1[0]) & or_tmp_440;
  assign mux_202_nl = MUX_s_1_2_2(and_131_cse, and_tmp_29, or_11_cse);
  assign IntSignedShiftRight_50U_5U_32U_obits_fixed_and_cse = core_wen & (~ and_dcpl_78)
      & (mux_202_nl);
  assign and_3358_cse = IsNaN_8U_23U_land_1_lpi_1_dfm_st_4 & (~ IsNaN_6U_10U_4_nor_tmp)
      & inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_5_1 & (inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_4_0_1==5'b11111);
  assign nor_35_cse = ~(inp_lookup_1_FpMul_6U_10U_1_oelse_1_acc_itm_7_1 | FpMul_6U_10U_1_if_2_FpMul_6U_10U_1_if_2_or_tmp
      | (~ inp_lookup_1_FpMul_6U_10U_1_else_2_if_acc_itm_6_1));
  assign and_920_rgt = and_dcpl_423 & or_11_cse;
  assign or_456_nl = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[0]) | (cfg_precision_1_sva_st_80[0])
      | not_tmp_182;
  assign mux_212_nl = MUX_s_1_2_2((or_456_nl), mux_tmp_133, and_3358_cse);
  assign mux_213_nl = MUX_s_1_2_2((mux_212_nl), mux_tmp_133, nor_35_cse);
  assign inp_lookup_else_if_a0_and_8_cse = core_wen & (~ and_dcpl_78) & (~ (mux_213_nl));
  assign or_457_cse = inp_lookup_1_FpMul_6U_10U_1_oelse_1_acc_itm_7_1 | FpMul_6U_10U_1_if_2_FpMul_6U_10U_1_if_2_or_tmp;
  assign or_461_cse = (chn_inp_in_crt_sva_2_739_736_1[0]) | (cfg_precision_1_sva_st_91[0]);
  assign or_471_cse = (chn_inp_in_rsci_d_mxwt[736]) | (cfg_precision_rsci_d!=2'b10)
      | (~ chn_inp_in_rsci_bawt);
  assign FpMul_6U_10U_2_else_2_else_if_FpMul_6U_10U_2_else_2_else_if_or_3_cse = and_dcpl_453
      | and_dcpl_458;
  assign nor_44_cse = ~(FpMul_6U_10U_2_lor_6_lpi_1_dfm_st_3 | (~ inp_lookup_1_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs));
  assign FpMul_6U_10U_2_oelse_1_FpMul_6U_10U_2_oelse_1_or_11_cse = and_dcpl_459 |
      and_dcpl_427;
  assign FpMul_6U_10U_2_oelse_1_and_4_cse = core_wen & FpMul_6U_10U_2_oelse_1_FpMul_6U_10U_2_oelse_1_or_11_cse
      & (~ mux_197_itm);
  assign nand_728_cse_1 = ~((chn_inp_in_rsci_d_mxwt[737]) & chn_inp_in_rsci_bawt
      & (cfg_precision_rsci_d==2'b10));
  assign or_6252_cse = (~ (chn_inp_in_crt_sva_2_739_736_1[1])) | (cfg_precision_1_sva_st_91!=2'b10);
  assign or_6257_cse = (~ (chn_inp_in_crt_sva_1_739_395_1[342])) | (cfg_precision_1_sva_st_90[0]);
  assign and_936_rgt = and_dcpl_465 & (~ (chn_inp_in_crt_sva_2_739_736_1[1])) & or_11_cse;
  assign and_939_rgt = and_dcpl_468 & (~ (chn_inp_in_crt_sva_2_739_736_1[1])) & or_11_cse;
  assign and_941_rgt = and_dcpl_471 & or_11_cse;
  assign and_3056_cse = main_stage_v_2 & (chn_inp_in_crt_sva_2_739_736_1[1]);
  assign and_945_rgt = and_920_rgt & and_3056_cse & (~ (z_out_1[49]));
  assign and_950_rgt = nand_358_cse & (cfg_precision_1_sva_st_80==2'b10) & (chn_inp_in_crt_sva_3_739_736_1[1])
      & main_stage_v_3 & or_11_cse;
  assign and_953_rgt = and_920_rgt & and_3056_cse & (z_out_1[49]) & inp_lookup_2_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1;
  assign and_956_rgt = and_920_rgt & and_3056_cse & (z_out_1[49]) & (~ inp_lookup_2_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1);
  assign and_137_cse = main_stage_v_3 & (chn_inp_in_crt_sva_3_739_736_1[1]) & or_tmp_440;
  assign mux_239_nl = MUX_s_1_2_2(and_137_cse, and_tmp_35, or_11_cse);
  assign IntSignedShiftRight_50U_5U_32U_obits_fixed_and_3_cse = core_wen & (~ and_dcpl_78)
      & (mux_239_nl);
  assign and_3355_cse = (~ IsNaN_6U_10U_4_nor_1_tmp) & inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_6_5_1
      & (inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_6_4_0_1==5'b11111) & IsNaN_8U_23U_land_2_lpi_1_dfm_st_4;
  assign or_507_cse = (~ inp_lookup_2_FpMul_6U_10U_1_else_2_if_acc_itm_6_1) | inp_lookup_2_FpMul_6U_10U_1_oelse_1_acc_itm_7_1
      | FpMul_6U_10U_1_if_2_FpMul_6U_10U_1_if_2_or_2_tmp;
  assign IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_2_cse
      = and_dcpl_464 | and_dcpl_488;
  assign or_518_nl = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[1]) | mux_tmp_163;
  assign mux_250_nl = MUX_s_1_2_2(mux_tmp_171, (or_518_nl), or_507_cse);
  assign mux_251_nl = MUX_s_1_2_2((mux_250_nl), mux_tmp_171, and_3355_cse);
  assign inp_lookup_else_if_a0_and_9_cse = core_wen & (~ and_dcpl_78) & (~ (mux_251_nl));
  assign or_519_cse = inp_lookup_2_FpMul_6U_10U_1_oelse_1_acc_itm_7_1 | FpMul_6U_10U_1_if_2_FpMul_6U_10U_1_if_2_or_2_tmp;
  assign or_523_cse = (chn_inp_in_crt_sva_2_739_736_1[1]) | (cfg_precision_1_sva_st_91[0]);
  assign FpMul_6U_10U_2_else_2_else_if_FpMul_6U_10U_2_else_2_else_if_or_2_cse = (and_dcpl_423
      & (~ (chn_inp_in_crt_sva_2_739_736_1[1])) & and_dcpl_419) | and_dcpl_495;
  assign FpMul_6U_10U_2_oelse_1_and_5_cse = core_wen & IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_2_cse
      & (~ mux_197_itm);
  assign nand_693_cse = ~(main_stage_v_1 & (chn_inp_in_crt_sva_1_739_395_1[343])
      & (cfg_precision_1_sva_st_90==2'b10));
  assign nand_598_cse = ~((chn_inp_in_rsci_d_mxwt[738]) & chn_inp_in_rsci_bawt &
      (cfg_precision_rsci_d==2'b10));
  assign nor_1967_cse = ~((~ (chn_inp_in_crt_sva_2_739_736_1[2])) | (cfg_precision_1_sva_st_91!=2'b10));
  assign or_6272_cse = (~ (chn_inp_in_crt_sva_1_739_395_1[343])) | (cfg_precision_1_sva_st_90[0]);
  assign and_973_rgt = nor_1017_cse & (~ (chn_inp_in_crt_sva_2_739_736_1[2])) & or_11_cse;
  assign and_976_rgt = and_dcpl_504 & (~ (chn_inp_in_crt_sva_2_739_736_1[2])) & or_11_cse;
  assign and_978_rgt = IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_14 & (~ (chn_inp_in_crt_sva_2_739_736_1[2]))
      & or_11_cse;
  assign and_3054_cse = (chn_inp_in_crt_sva_2_739_736_1[2]) & main_stage_v_2;
  assign and_982_rgt = and_920_rgt & and_3054_cse & (~ (z_out_2[49]));
  assign and_987_rgt = or_tmp_277 & (cfg_precision_1_sva_st_80==2'b10) & (chn_inp_in_crt_sva_3_739_736_1[2])
      & main_stage_v_3 & or_11_cse;
  assign and_990_rgt = and_920_rgt & and_3054_cse & (z_out_2[49]) & inp_lookup_3_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1;
  assign and_993_rgt = and_920_rgt & and_3054_cse & (z_out_2[49]) & (~ inp_lookup_3_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1);
  assign and_144_cse = main_stage_v_3 & (chn_inp_in_crt_sva_3_739_736_1[2]) & or_tmp_440;
  assign mux_277_nl = MUX_s_1_2_2(and_144_cse, and_tmp_42, or_11_cse);
  assign IntSignedShiftRight_50U_5U_32U_obits_fixed_and_6_cse = core_wen & (~ and_dcpl_78)
      & (mux_277_nl);
  assign and_3351_cse = (~ IsNaN_6U_10U_4_nor_2_tmp) & inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_6_5_1
      & (inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_6_4_0_1==5'b11111) & IsNaN_8U_23U_land_3_lpi_1_dfm_st_4;
  assign nor_55_cse = ~(inp_lookup_3_FpMul_6U_10U_1_oelse_1_acc_itm_7_1 | FpMul_6U_10U_1_if_2_FpMul_6U_10U_1_if_2_or_4_tmp
      | (~ inp_lookup_3_FpMul_6U_10U_1_else_2_if_acc_itm_6_1));
  assign IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_1_cse
      = and_dcpl_496 | and_dcpl_524;
  assign or_579_nl = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[2]) | mux_tmp_201;
  assign mux_288_nl = MUX_s_1_2_2((or_579_nl), mux_tmp_209, nor_55_cse);
  assign mux_289_nl = MUX_s_1_2_2((mux_288_nl), mux_tmp_209, and_3351_cse);
  assign inp_lookup_else_if_a0_and_10_cse = core_wen & (~ and_dcpl_78) & (~ (mux_289_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_or_cse
      = (and_dcpl_498 & and_dcpl_524) | and_dcpl_530;
  assign or_582_nl = nor_55_cse | and_348_cse;
  assign mux_290_nl = MUX_s_1_2_2(and_tmp_48, (or_582_nl), or_11_cse);
  assign mux_291_nl = MUX_s_1_2_2(nand_tmp_18, (mux_290_nl), nor_275_cse);
  assign nor_1634_nl = ~((~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ and_tmp_48));
  assign mux_292_nl = MUX_s_1_2_2(nand_tmp_18, (nor_1634_nl), cfg_precision_1_sva_st_90[1]);
  assign mux_293_nl = MUX_s_1_2_2((mux_292_nl), nand_tmp_18, or_604_cse);
  assign nor_1635_nl = ~((~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (main_stage_v_3 & (~ or_tmp_584)));
  assign mux_294_nl = MUX_s_1_2_2((nor_1635_nl), nand_tmp_18, or_802_cse);
  assign mux_295_nl = MUX_s_1_2_2((mux_294_nl), (mux_293_nl), main_stage_v_1);
  assign mux_296_nl = MUX_s_1_2_2((mux_295_nl), (mux_291_nl), main_stage_v_2);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_and_cse = FpAdd_8U_23U_o_expo_and_cse
      & FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_or_cse
      & (mux_296_nl);
  assign or_593_cse = inp_lookup_3_FpMul_6U_10U_1_oelse_1_acc_itm_7_1 | FpMul_6U_10U_1_if_2_FpMul_6U_10U_1_if_2_or_4_tmp;
  assign or_597_cse = (chn_inp_in_crt_sva_2_739_736_1[2]) | (cfg_precision_1_sva_st_91[0]);
  assign or_604_cse = (chn_inp_in_crt_sva_1_739_395_1[343]) | (cfg_precision_1_sva_st_90[0]);
  assign nor_67_cse = ~(FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_3 | (~ inp_lookup_3_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs));
  assign FpMul_6U_10U_2_oelse_1_and_6_cse = core_wen & IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_1_cse
      & (~ mux_197_itm);
  assign mux_74_nl = MUX_v_23_2_2(FpAdd_8U_23U_FpAdd_8U_23U_or_7_itm, reg_chn_inp_in_crt_sva_3_606_576_1_reg,
      IsNaN_6U_10U_7_land_lpi_1_dfm_6);
  assign FpAdd_8U_23U_o_mant_not_3_nl = ~ (fsm_output[0]);
  assign and_3424_nl = MUX_v_23_2_2(23'b00000000000000000000000, (mux_74_nl), (FpAdd_8U_23U_o_mant_not_3_nl));
  assign and_1004_nl = and_dcpl_423 & (chn_inp_in_crt_sva_2_739_736_1[3]) & and_dcpl_419;
  assign mux_1993_rgt = MUX_v_31_2_2(({8'b0 , (and_3424_nl)}), ({reg_chn_inp_in_crt_sva_2_606_576_itm
      , reg_chn_inp_in_crt_sva_2_606_576_1_itm}), and_1004_nl);
  assign nand_701_cse = ~(main_stage_v_2 & (chn_inp_in_crt_sva_2_739_736_1[3]) &
      (cfg_precision_1_sva_st_91==2'b10));
  assign nor_1743_rgt = ~(IsNaN_6U_10U_2_land_lpi_1_dfm_st_14 | IsNaN_6U_10U_7_land_lpi_1_dfm_5
      | (chn_inp_in_crt_sva_2_739_736_1[3]) | (~ or_11_cse));
  assign and_1012_rgt = and_dcpl_539 & (~ (chn_inp_in_crt_sva_2_739_736_1[3])) &
      or_11_cse;
  assign and_1014_rgt = IsNaN_6U_10U_2_land_lpi_1_dfm_st_14 & (~ (chn_inp_in_crt_sva_2_739_736_1[3]))
      & or_11_cse;
  assign and_1018_rgt = and_920_rgt & and_3346_cse & (~ (z_out_3[49]));
  assign and_1023_rgt = nand_701_cse & (cfg_precision_1_sva_st_80==2'b10) & (chn_inp_in_crt_sva_3_739_736_1[3])
      & main_stage_v_3 & or_11_cse;
  assign and_1026_rgt = and_920_rgt & and_3346_cse & (z_out_3[49]) & inp_lookup_4_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1;
  assign and_1029_rgt = and_920_rgt & and_3346_cse & (z_out_3[49]) & (~ inp_lookup_4_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1);
  assign and_152_cse = main_stage_v_3 & (chn_inp_in_crt_sva_3_739_736_1[3]) & or_tmp_440;
  assign mux_320_nl = MUX_s_1_2_2(and_152_cse, and_tmp_50, or_11_cse);
  assign IntSignedShiftRight_50U_5U_32U_obits_fixed_and_9_cse = core_wen & (~ and_dcpl_78)
      & (mux_320_nl);
  assign and_3345_cse = (~ IsNaN_6U_10U_4_nor_3_tmp) & inp_lookup_else_if_a0_15_10_lpi_1_dfm_6_5_1
      & (inp_lookup_else_if_a0_15_10_lpi_1_dfm_6_4_0_1==5'b11111) & IsNaN_8U_23U_land_lpi_1_dfm_st_4;
  assign IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_cse
      = and_dcpl_535 | and_dcpl_559;
  assign and_3344_nl = inp_lookup_else_if_a0_15_10_lpi_1_dfm_6_5_1 & (inp_lookup_else_if_a0_15_10_lpi_1_dfm_6_4_0_1==5'b11111)
      & IsNaN_8U_23U_land_lpi_1_dfm_st_4;
  assign mux_341_nl = MUX_s_1_2_2(mux_tmp_262, (~ mux_tmp_260), and_3344_nl);
  assign mux_342_nl = MUX_s_1_2_2((mux_341_nl), mux_tmp_262, IsNaN_6U_10U_4_nor_3_tmp);
  assign mux_343_nl = MUX_s_1_2_2(nand_tmp_24, (mux_342_nl), nor_74_cse);
  assign inp_lookup_else_if_a0_and_11_cse = core_wen & (~ and_dcpl_78) & (~ (mux_343_nl));
  assign or_648_cse = inp_lookup_4_FpMul_6U_10U_1_oelse_1_acc_itm_7_1 | FpMul_6U_10U_1_if_2_FpMul_6U_10U_1_if_2_or_6_tmp;
  assign FpMul_6U_10U_2_oelse_1_and_7_cse = core_wen & IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_cse
      & (~ mux_197_itm);
  assign FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_or_6_cse = and_dcpl_564
      | and_dcpl_565;
  assign or_671_nl = (cfg_precision_1_sva_st_80!=2'b10) | IsNaN_6U_10U_5_land_1_lpi_1_dfm_5
      | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_15;
  assign mux_352_nl = MUX_s_1_2_2((or_671_nl), or_tmp_440, chn_inp_in_crt_sva_3_739_736_1[0]);
  assign and_3340_nl = main_stage_v_3 & (~ (mux_352_nl));
  assign or_672_nl = (~ (chn_inp_in_crt_sva_4_739_736_1[0])) | (cfg_precision_1_sva_st_81!=2'b10);
  assign or_674_nl = (cfg_precision_1_sva_st_81!=2'b10) | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_16;
  assign mux_353_nl = MUX_s_1_2_2((or_674_nl), or_3379_cse, chn_inp_in_crt_sva_4_739_736_1[0]);
  assign mux_354_nl = MUX_s_1_2_2((mux_353_nl), (or_672_nl), IsNaN_6U_10U_5_land_1_lpi_1_dfm_6);
  assign and_3341_nl = main_stage_v_4 & (~ (mux_354_nl));
  assign mux_355_nl = MUX_s_1_2_2((and_3341_nl), (and_3340_nl), or_11_cse);
  assign FpAdd_8U_23U_1_is_a_greater_oelse_and_cse = core_wen & FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_or_6_cse
      & (mux_355_nl);
  assign cfg_precision_and_12_cse = core_wen & (~ and_dcpl_78) & mux_tmp_278;
  assign FpMul_6U_10U_2_o_expo_and_cse = core_wen & ((and_dcpl_567 & or_11_cse) |
      and_dcpl_575) & mux_tmp_278;
  assign nor_1622_nl = ~((~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[0])
      | (cfg_precision_1_sva_st_80[0]) | not_tmp_282);
  assign nor_1623_nl = ~((~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[0])
      | (cfg_precision_1_sva_st_81!=2'b10) | (~ IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_16));
  assign mux_367_nl = MUX_s_1_2_2((nor_1623_nl), (nor_1622_nl), or_11_cse);
  assign inp_lookup_else_if_a0_and_12_cse = core_wen & (~ and_dcpl_78) & (mux_367_nl);
  assign or_683_cse = (chn_inp_in_crt_sva_1_739_395_1[341]) | (cfg_precision_1_sva_st_90!=2'b10);
  assign and_1049_rgt = IsNaN_6U_10U_5_land_1_lpi_1_dfm_5 & (cfg_precision_1_sva_st_80[1])
      & and_dcpl_454 & and_dcpl_560;
  assign and_1052_rgt = (~ IsNaN_6U_10U_5_land_1_lpi_1_dfm_5) & (cfg_precision_1_sva_st_80[1])
      & and_dcpl_454 & and_dcpl_560;
  assign IsNaN_6U_10U_5_aelse_and_4_cse = core_wen & (~ and_dcpl_78) & (~ mux_461_cse);
  assign FpMul_6U_10U_1_oelse_1_and_5_cse = core_wen & FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_or_6_cse
      & (~ mux_461_cse);
  assign FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_or_5_cse = and_dcpl_582
      | and_dcpl_583;
  assign or_720_nl = IsNaN_6U_10U_5_land_2_lpi_1_dfm_5 | (cfg_precision_1_sva_st_80!=2'b10)
      | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_15;
  assign mux_383_nl = MUX_s_1_2_2((or_720_nl), or_tmp_440, chn_inp_in_crt_sva_3_739_736_1[1]);
  assign and_3335_nl = main_stage_v_3 & (~ (mux_383_nl));
  assign or_721_nl = (~ (chn_inp_in_crt_sva_4_739_736_1[1])) | (cfg_precision_1_sva_st_81!=2'b10);
  assign or_723_nl = (cfg_precision_1_sva_st_81!=2'b10) | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_16;
  assign mux_384_nl = MUX_s_1_2_2((or_723_nl), or_3379_cse, chn_inp_in_crt_sva_4_739_736_1[1]);
  assign mux_385_nl = MUX_s_1_2_2((mux_384_nl), (or_721_nl), IsNaN_6U_10U_5_land_2_lpi_1_dfm_6);
  assign and_3336_nl = main_stage_v_4 & (~ (mux_385_nl));
  assign mux_386_nl = MUX_s_1_2_2((and_3336_nl), (and_3335_nl), or_11_cse);
  assign FpAdd_8U_23U_1_is_a_greater_oelse_and_1_cse = core_wen & FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_or_5_cse
      & (mux_386_nl);
  assign FpMul_6U_10U_2_o_expo_and_3_cse = core_wen & ((and_dcpl_585 & or_11_cse)
      | and_dcpl_593) & mux_tmp_278;
  assign nor_1615_nl = ~((~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[1])
      | (cfg_precision_1_sva_st_80!=2'b10) | (~ IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_15));
  assign nor_1616_nl = ~((~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[1])
      | (cfg_precision_1_sva_st_81!=2'b10) | (~ IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_16));
  assign mux_407_nl = MUX_s_1_2_2((nor_1616_nl), (nor_1615_nl), or_11_cse);
  assign inp_lookup_else_if_a0_and_14_cse = core_wen & (~ and_dcpl_78) & (mux_407_nl);
  assign or_740_cse = (chn_inp_in_crt_sva_1_739_395_1[342]) | (cfg_precision_1_sva_st_90!=2'b10);
  assign mux_400_cse = MUX_s_1_2_2(or_763_cse, or_740_cse, main_stage_v_1);
  assign and_1068_rgt = and_dcpl_584 & IsNaN_6U_10U_5_land_2_lpi_1_dfm_5 & (~ (chn_inp_in_crt_sva_3_739_736_1[1]))
      & and_dcpl_560;
  assign and_1071_rgt = and_dcpl_584 & and_dcpl_597 & and_dcpl_560;
  assign or_763_cse = (~ chn_inp_in_rsci_bawt) | (cfg_precision_rsci_d!=2'b10) |
      (chn_inp_in_rsci_d_mxwt[737]);
  assign FpMul_6U_10U_1_oelse_1_and_7_cse = core_wen & FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_or_5_cse
      & (~ mux_461_cse);
  assign FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_or_4_cse = and_dcpl_600
      | and_dcpl_601;
  assign or_772_nl = IsNaN_6U_10U_5_land_3_lpi_1_dfm_5 | (cfg_precision_1_sva_st_80!=2'b10)
      | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_15;
  assign mux_423_nl = MUX_s_1_2_2((or_772_nl), or_tmp_440, chn_inp_in_crt_sva_3_739_736_1[2]);
  assign and_3330_nl = main_stage_v_3 & (~ (mux_423_nl));
  assign or_774_nl = IsNaN_6U_10U_5_land_3_lpi_1_dfm_6 | (cfg_precision_1_sva_st_81!=2'b10)
      | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_16;
  assign mux_424_nl = MUX_s_1_2_2((or_774_nl), or_3379_cse, chn_inp_in_crt_sva_4_739_736_1[2]);
  assign and_3331_nl = main_stage_v_4 & (~ (mux_424_nl));
  assign mux_425_nl = MUX_s_1_2_2((and_3331_nl), (and_3330_nl), or_11_cse);
  assign FpAdd_8U_23U_1_is_a_greater_oelse_and_2_cse = core_wen & FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_or_4_cse
      & (mux_425_nl);
  assign FpMul_6U_10U_2_o_expo_and_6_cse = core_wen & ((and_dcpl_603 & or_11_cse)
      | and_dcpl_611) & mux_tmp_278;
  assign nor_1608_nl = ~((~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[2])
      | (cfg_precision_1_sva_st_80!=2'b10) | (~ IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_15));
  assign nor_1609_nl = ~((~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[2])
      | (cfg_precision_1_sva_st_81!=2'b10) | (~ IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_16));
  assign mux_439_nl = MUX_s_1_2_2((nor_1609_nl), (nor_1608_nl), or_11_cse);
  assign inp_lookup_else_if_a0_and_16_cse = core_wen & (~ and_dcpl_78) & (mux_439_nl);
  assign or_792_cse = (chn_inp_in_crt_sva_3_739_736_1[2]) | (cfg_precision_1_sva_st_80[0]);
  assign or_801_cse = (cfg_precision_1_sva_st_90!=2'b10) | (chn_inp_in_crt_sva_1_739_395_1[343]);
  assign or_802_cse = (~ chn_inp_in_rsci_bawt) | (cfg_precision_rsci_d!=2'b10) |
      (chn_inp_in_rsci_d_mxwt[738]);
  assign and_1099_rgt = and_dcpl_584 & IsNaN_6U_10U_5_land_3_lpi_1_dfm_5 & (~ (chn_inp_in_crt_sva_3_739_736_1[2]))
      & and_dcpl_560;
  assign and_1102_rgt = and_dcpl_584 & and_dcpl_627 & and_dcpl_560;
  assign FpMul_6U_10U_1_oelse_1_and_9_cse = core_wen & FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_or_4_cse
      & (~ mux_461_cse);
  assign FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_4_cse = and_dcpl_630 | and_dcpl_631;
  assign mux_461_cse = MUX_s_1_2_2(or_3850_cse, or_2282_cse, or_11_cse);
  assign IsNaN_8U_23U_2_aelse_and_cse = core_wen & FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_4_cse
      & (~ mux_461_cse);
  assign and_3327_nl = main_stage_v_3 & (~((~((~(IsNaN_6U_10U_5_land_lpi_1_dfm_5
      | IsNaN_6U_10U_2_land_lpi_1_dfm_st_15)) | (chn_inp_in_crt_sva_3_739_736_1[3])))
      | (cfg_precision_1_sva_st_80!=2'b10)));
  assign or_833_nl = IsNaN_6U_10U_4_land_lpi_1_dfm_5 | IsNaN_6U_10U_5_land_lpi_1_dfm_6
      | (cfg_precision_1_sva_st_81!=2'b10);
  assign mux_465_nl = MUX_s_1_2_2((or_833_nl), or_3379_cse, chn_inp_in_crt_sva_4_739_736_1[3]);
  assign and_3328_nl = main_stage_v_4 & (~ (mux_465_nl));
  assign mux_466_nl = MUX_s_1_2_2((and_3328_nl), (and_3327_nl), or_11_cse);
  assign FpAdd_8U_23U_1_is_a_greater_oelse_and_3_cse = core_wen & FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_4_cse
      & (mux_466_nl);
  assign FpMul_6U_10U_2_o_expo_and_9_cse = core_wen & ((and_dcpl_633 & or_11_cse)
      | and_dcpl_641) & mux_tmp_278;
  assign or_654_nl = (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[3]) | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_467_nl = MUX_s_1_2_2(nand_tmp_50, (or_654_nl), or_11_cse);
  assign mux_468_nl = MUX_s_1_2_2(nand_tmp_50, or_2282_cse, or_11_cse);
  assign mux_469_nl = MUX_s_1_2_2((mux_468_nl), (mux_467_nl), FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_3);
  assign IsNaN_6U_10U_4_aelse_and_cse = core_wen & FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_4_cse
      & (~ (mux_469_nl));
  assign nor_1596_nl = ~((~ main_stage_v_3) | (~ IsNaN_6U_10U_2_land_lpi_1_dfm_st_15)
      | (chn_inp_in_crt_sva_3_739_736_1[3]) | (cfg_precision_1_sva_st_80!=2'b10));
  assign nor_1597_nl = ~((~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[3])
      | (~ IsNaN_6U_10U_4_land_lpi_1_dfm_5) | (cfg_precision_1_sva_st_81!=2'b10));
  assign mux_470_nl = MUX_s_1_2_2((nor_1597_nl), (nor_1596_nl), or_11_cse);
  assign inp_lookup_else_if_a0_and_18_cse = core_wen & (~ and_dcpl_78) & (mux_470_nl);
  assign FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_3_cse = and_dcpl_654 | and_dcpl_655;
  assign and_1131_rgt = or_11_cse & inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5;
  assign mux_475_nl = MUX_s_1_2_2(main_stage_v_5, main_stage_v_4, or_11_cse);
  assign cfg_precision_and_16_cse = core_wen & (~ and_dcpl_78) & (mux_475_nl);
  assign mux_476_cse = MUX_s_1_2_2((~ chn_inp_in_crt_sva_4_411_1), chn_inp_in_crt_sva_4_411_1,
      inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5);
  assign nor_1593_cse = ~((~ IsNaN_8U_23U_2_land_1_lpi_1_dfm_st_7) | chn_inp_in_crt_sva_5_411_1);
  assign and_1127_nl = or_11_cse & (~ FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5);
  assign FpMul_6U_10U_2_o_mant_asn_FpMul_6U_10U_2_o_mant_conc_80_cgspt_7_mux_nl =
      MUX_v_8_2_2((chn_inp_in_crt_sva_4_127_0_1[30:23]), ({reg_FpAdd_8U_23U_o_expo_1_lpi_1_dfm_11_reg
      , reg_FpAdd_8U_23U_o_expo_1_lpi_1_dfm_11_1_reg}), and_1127_nl);
  assign mux_1897_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_5_739_736_1[0]), (chn_inp_in_crt_sva_4_739_736_1[0]),
      or_11_cse);
  assign FpMul_6U_10U_2_o_mant_mux1h_1_itm = MUX_v_10_2_2(FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_8,
      ({2'b0 , (FpMul_6U_10U_2_o_mant_asn_FpMul_6U_10U_2_o_mant_conc_80_cgspt_7_mux_nl)}),
      mux_1897_nl);
  assign or_5950_cse = (FpMul_6U_10U_1_o_mant_1_lpi_1_dfm_3!=10'b0000000000);
  assign and_4141_cse = (FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_3_3_0_mx1w1==4'b1111);
  assign and_3637_cse = inp_lookup_1_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp &
      (~ FpAdd_6U_10U_1_is_a_greater_acc_itm_6);
  assign xnor_6_cse = ~(chn_inp_in_crt_sva_4_411_1 ^ inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5);
  assign and_4164_cse = (~(inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_8_5_1 & (inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_8_4_0_1[4])))
      & or_tmp_4675;
  assign and_4165_cse = (~(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_9_1
      & FpAdd_8U_23U_o_sign_1_lpi_1_dfm_8)) & or_tmp_4675;
  assign nor_1883_cse = ~(nor_1896_cse | (cfg_precision_1_sva_st_81[0]));
  assign FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_2_cse = and_dcpl_662 | and_dcpl_663;
  assign and_1139_rgt = or_11_cse & inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5;
  assign mux_485_cse = MUX_s_1_2_2((~ chn_inp_in_crt_sva_4_427_1), chn_inp_in_crt_sva_4_427_1,
      inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5);
  assign nor_1587_cse = ~((~ IsNaN_8U_23U_2_land_2_lpi_1_dfm_st_7) | chn_inp_in_crt_sva_5_427_1);
  assign and_1135_nl = or_11_cse & (~ FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5);
  assign FpMul_6U_10U_2_o_mant_asn_FpMul_6U_10U_2_o_mant_conc_81_cgspt_7_mux_nl =
      MUX_v_8_2_2((chn_inp_in_crt_sva_4_127_0_1[62:55]), ({reg_FpAdd_8U_23U_o_expo_2_lpi_1_dfm_11_reg
      , reg_FpAdd_8U_23U_o_expo_2_lpi_1_dfm_11_1_reg}), and_1135_nl);
  assign mux_1898_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_5_739_736_1[1]), (chn_inp_in_crt_sva_4_739_736_1[1]),
      or_11_cse);
  assign FpMul_6U_10U_2_o_mant_mux1h_3_itm = MUX_v_10_2_2(FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_8,
      ({2'b0 , (FpMul_6U_10U_2_o_mant_asn_FpMul_6U_10U_2_o_mant_conc_81_cgspt_7_mux_nl)}),
      mux_1898_nl);
  assign or_5967_cse = (FpMul_6U_10U_1_o_mant_2_lpi_1_dfm_3!=10'b0000000000);
  assign and_4136_cse = (FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_3_3_0_mx1w1==4'b1111);
  assign and_3663_cse = inp_lookup_2_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp &
      (~ FpAdd_6U_10U_1_is_a_greater_acc_1_itm_6);
  assign xnor_4_cse = ~(chn_inp_in_crt_sva_4_427_1 ^ inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5);
  assign and_4159_cse = (~(inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_8_5_1 & (inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_8_4_0_1[4])))
      & or_tmp_4685;
  assign and_4160_cse = (~(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_9_1
      & FpAdd_8U_23U_o_sign_2_lpi_1_dfm_8)) & or_tmp_4685;
  assign FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_1_cse = and_dcpl_670 | and_dcpl_671;
  assign and_1147_rgt = or_11_cse & inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5;
  assign mux_500_cse = MUX_s_1_2_2((~ chn_inp_in_crt_sva_4_443_1), chn_inp_in_crt_sva_4_443_1,
      inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5);
  assign nor_1584_cse = ~((~ IsNaN_8U_23U_2_land_3_lpi_1_dfm_st_7) | chn_inp_in_crt_sva_5_443_1);
  assign FpMul_6U_10U_1_o_mant_mux1h_1_itm = MUX_v_10_2_2(FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_3_mx0w1,
      ({2'b0 , reg_FpAdd_8U_23U_o_expo_3_lpi_1_dfm_11_reg , reg_FpAdd_8U_23U_o_expo_3_lpi_1_dfm_11_1_reg}),
      mux_tmp_1821);
  assign or_5985_cse = (FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_3_mx0w1!=10'b0000000000);
  assign and_3689_cse = inp_lookup_3_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp &
      (~ FpAdd_6U_10U_1_is_a_greater_acc_2_itm_6);
  assign xnor_2_cse = ~(chn_inp_in_crt_sva_4_443_1 ^ inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5);
  assign nor_1877_cse = ~(nor_1896_cse | (chn_inp_in_crt_sva_4_739_736_1[2]));
  assign and_1143_nl = or_11_cse & (~ FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5);
  assign FpMul_6U_10U_2_o_mant_asn_FpMul_6U_10U_2_o_mant_conc_82_cgspt_7_mux_nl =
      MUX_v_8_2_2((chn_inp_in_crt_sva_4_127_0_1[94:87]), ({reg_FpAdd_8U_23U_o_expo_3_lpi_1_dfm_11_reg
      , reg_FpAdd_8U_23U_o_expo_3_lpi_1_dfm_11_1_reg}), and_1143_nl);
  assign FpMul_6U_10U_2_o_mant_mux1h_5_itm = MUX_v_10_2_2(FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_8,
      ({2'b0 , (FpMul_6U_10U_2_o_mant_asn_FpMul_6U_10U_2_o_mant_conc_82_cgspt_7_mux_nl)}),
      mux_tmp_1821);
  assign and_4126_cse = (FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_3_0_mx1w1==4'b1111);
  assign and_4154_cse = (~(inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_8_5_1 & (inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_8_4_0_1[4])))
      & or_tmp_4703;
  assign and_4155_cse = (~(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_9_1
      & FpAdd_8U_23U_o_sign_3_lpi_1_dfm_9)) & or_tmp_4703;
  assign IsNaN_8U_23U_2_aelse_IsNaN_8U_23U_2_aelse_or_cse = and_dcpl_678 | and_dcpl_679;
  assign nand_579_cse = ~(main_stage_v_4 & (chn_inp_in_crt_sva_4_739_736_1[3]) &
      (cfg_precision_1_sva_st_81==2'b10));
  assign and_1155_rgt = or_11_cse & inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4;
  assign and_1151_nl = or_11_cse & (~ FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5);
  assign mux_2004_nl = MUX_v_8_2_2((chn_inp_in_crt_sva_4_127_0_1[126:119]), ({reg_FpAdd_8U_23U_o_expo_lpi_1_dfm_11_reg
      , reg_FpAdd_8U_23U_o_expo_lpi_1_dfm_11_1_reg}), and_1151_nl);
  assign mux_1900_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_5_739_736_1[3]), (chn_inp_in_crt_sva_4_739_736_1[3]),
      or_11_cse);
  assign FpMul_6U_10U_2_o_mant_FpMul_6U_10U_2_o_mant_mux_rgt = MUX_v_10_2_2(FpMul_6U_10U_2_o_mant_lpi_1_dfm_7,
      ({2'b0 , (mux_2004_nl)}), mux_1900_nl);
  assign and_3483_cse = or_11_cse & core_wen;
  assign nor_126_cse = ~(inp_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_1_itm_7_1 | (~ (FpAdd_8U_23U_1_int_mant_p1_1_sva_3[49])));
  assign and_1163_rgt = or_11_cse & IsNaN_8U_23U_3_land_1_lpi_1_dfm_6;
  assign IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_4_cse = and_dcpl_690 | and_dcpl_691;
  assign IsNaN_8U_23U_3_aelse_and_cse = core_wen & IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_4_cse
      & (~ mux_516_itm);
  assign and_1166_nl = IsNaN_8U_23U_2_land_1_lpi_1_dfm_9 & (chn_inp_in_crt_sva_5_739_736_1[0]);
  assign and_3443_nl = IsNaN_6U_10U_8_land_1_lpi_1_dfm_st_3 & (chn_inp_in_crt_sva_6_739_736_1[0]);
  assign mux_1901_tmp = MUX_s_1_2_2((and_3443_nl), (and_1166_nl), or_11_cse);
  assign mux_517_nl = MUX_s_1_2_2(or_tmp_962, or_tmp_850, or_11_cse);
  assign FpMantRNE_49U_24U_1_else_and_cse = core_wen & (~ and_dcpl_78) & (~ (mux_517_nl));
  assign mux_518_nl = MUX_s_1_2_2(main_stage_v_6, main_stage_v_5, or_11_cse);
  assign cfg_precision_and_20_cse = core_wen & (~ and_dcpl_78) & (mux_518_nl);
  assign and_1174_rgt = or_11_cse & IsNaN_8U_23U_3_land_2_lpi_1_dfm_6;
  assign IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_3_cse = and_dcpl_701 | and_dcpl_702;
  assign IsNaN_8U_23U_3_aelse_and_1_cse = core_wen & IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_3_cse
      & (~ mux_530_itm);
  assign and_1177_nl = IsNaN_8U_23U_2_land_2_lpi_1_dfm_9 & (chn_inp_in_crt_sva_5_739_736_1[1]);
  assign and_3444_nl = IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_4 & (chn_inp_in_crt_sva_6_739_736_1[1]);
  assign mux_1902_tmp = MUX_s_1_2_2((and_3444_nl), (and_1177_nl), or_11_cse);
  assign mux_531_nl = MUX_s_1_2_2(or_tmp_992, or_tmp_880, or_11_cse);
  assign FpMantRNE_49U_24U_1_else_and_2_cse = core_wen & (~ and_dcpl_78) & (~ (mux_531_nl));
  assign FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_1_cse = ~(inp_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_1_itm_7_1
      | (~ (FpAdd_8U_23U_1_int_mant_p1_2_sva_3[49])));
  assign IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_2_cse = and_dcpl_712 | and_dcpl_713;
  assign IsNaN_8U_23U_3_aelse_and_2_cse = core_wen & IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_2_cse
      & (~ mux_540_itm);
  assign and_1188_nl = IsNaN_8U_23U_2_land_3_lpi_1_dfm_9 & (chn_inp_in_crt_sva_5_739_736_1[2]);
  assign mux_1903_tmp = MUX_s_1_2_2(nor_tmp_686, (and_1188_nl), or_11_cse);
  assign mux_541_nl = MUX_s_1_2_2(or_tmp_1009, or_tmp_899, or_11_cse);
  assign FpMantRNE_49U_24U_1_else_and_4_cse = core_wen & (~ and_dcpl_78) & (~ (mux_541_nl));
  assign FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_2_cse = ~(inp_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_1_itm_7
      | (~ (FpAdd_8U_23U_1_int_mant_p1_3_sva_3[49])));
  assign nor_136_cse = ~(inp_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_1_itm_7_1 | (~ (FpAdd_8U_23U_1_int_mant_p1_sva_3[49])));
  assign and_1192_rgt = or_11_cse & IsNaN_8U_23U_3_land_lpi_1_dfm_5;
  assign IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_1_cse = and_dcpl_719 | and_dcpl_720;
  assign IsNaN_8U_23U_3_aelse_and_3_cse = core_wen & IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_1_cse
      & (~ mux_516_itm);
  assign and_1195_nl = IsNaN_8U_23U_2_land_lpi_1_dfm_9 & (chn_inp_in_crt_sva_5_739_736_1[3]);
  assign and_3446_nl = IsNaN_6U_10U_8_land_lpi_1_dfm_st_4 & (chn_inp_in_crt_sva_6_739_736_1[3]);
  assign mux_1904_tmp = MUX_s_1_2_2((and_3446_nl), (and_1195_nl), or_11_cse);
  assign mux_552_nl = MUX_s_1_2_2(or_tmp_1038, or_tmp_945, or_11_cse);
  assign FpMantRNE_49U_24U_1_else_and_6_cse = core_wen & (~ and_dcpl_78) & (~ (mux_552_nl));
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_and_cse = core_wen & (~ and_dcpl_78)
      & (~ mux_559_itm);
  assign and_1209_rgt = ((~ inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8)
      | inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7 | (~ inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8))
      & or_11_cse;
  assign nor_1546_cse = ~((~ inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2)
      | inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
      | (~ (chn_inp_in_crt_sva_7_739_736_1[0])) | (cfg_precision_1_sva_st_84!=2'b10)
      | (~ main_stage_v_7));
  assign and_1211_rgt = or_11_cse & (~ IsNaN_6U_10U_8_land_1_lpi_1_dfm_st_3);
  assign and_1213_rgt = or_11_cse & (~ inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8);
  assign mux_567_nl = MUX_s_1_2_2(main_stage_v_7, main_stage_v_6, or_11_cse);
  assign cfg_precision_and_24_cse = core_wen & (~ and_dcpl_78) & (mux_567_nl);
  assign or_4591_tmp = (cfg_precision_1_sva_st_83[0]) | (~ (chn_inp_in_crt_sva_6_739_736_1[0]))
      | (~ (cfg_precision_1_sva_st_83[1]));
  assign FpAdd_6U_10U_1_and_47_rgt = (~ or_4591_tmp) & and_dcpl_741;
  assign and_1217_rgt = or_11_cse & (~ IsNaN_8U_23U_3_land_1_lpi_1_dfm_7);
  assign FpNormalize_6U_23U_1_if_FpNormalize_6U_23U_1_if_or_3_cse = and_dcpl_740
      | and_dcpl_741;
  assign and_1221_rgt = ((~ inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8)
      | inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7 | (~ inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8))
      & or_11_cse;
  assign and_1223_rgt = or_11_cse & (~ IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_4);
  assign and_1225_rgt = or_11_cse & (~ inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_if_and_2_cse = core_wen & (~ and_dcpl_78)
      & (~ mux_573_itm);
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_14_cse = and_dcpl_752 | and_dcpl_753;
  assign and_1229_rgt = or_11_cse & (~ IsNaN_8U_23U_3_land_2_lpi_1_dfm_7);
  assign IsNaN_6U_10U_8_aelse_and_cse = core_wen & FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_14_cse
      & (~ mux_586_itm);
  assign and_1233_rgt = ((~ inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8)
      | inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7 | (~ inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8))
      & or_11_cse;
  assign nor_1517_cse = ~(inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
      | (~ inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2)
      | (~ main_stage_v_7) | (~ (chn_inp_in_crt_sva_7_739_736_1[2])) | (cfg_precision_1_sva_st_84!=2'b10));
  assign and_1235_rgt = or_11_cse & (~ IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_4);
  assign and_1237_rgt = or_11_cse & (~ inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_if_and_4_cse = core_wen & (~ and_dcpl_78)
      & (~ mux_587_itm);
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_13_cse = and_dcpl_764 | and_dcpl_765;
  assign and_1241_rgt = or_11_cse & (~ IsNaN_8U_23U_3_land_3_lpi_1_dfm_7);
  assign IsNaN_6U_10U_8_aelse_and_1_cse = core_wen & FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_13_cse
      & (~ mux_854_cse);
  assign and_1245_rgt = ((~ inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8)
      | inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7 | (~ inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8))
      & or_11_cse;
  assign and_1247_rgt = or_11_cse & (~ IsNaN_6U_10U_8_land_lpi_1_dfm_st_4);
  assign and_1249_rgt = or_11_cse & (~ inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_if_and_6_cse = core_wen & (~ and_dcpl_78)
      & (~ mux_599_itm);
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_12_cse = and_dcpl_776 | and_dcpl_777;
  assign and_1253_rgt = or_11_cse & (~ IsNaN_8U_23U_3_land_lpi_1_dfm_6);
  assign IsNaN_6U_10U_8_aelse_and_2_cse = core_wen & FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_12_cse
      & (~ mux_854_cse);
  assign nand_62_nl = ~((chn_inp_in_crt_sva_7_739_736_1[0]) & (~((~(IsNaN_6U_10U_IsNaN_6U_10U_nor_tmp
      | (~ FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_tmp))) | (cfg_precision_1_sva_st_84!=2'b10)
      | (~ main_stage_v_7))));
  assign mux_614_nl = MUX_s_1_2_2(or_tmp_1255, or_tmp_1253, reg_FpMul_6U_10U_lor_3_lpi_1_dfm_3_cse);
  assign mux_615_cse = MUX_s_1_2_2((mux_614_nl), (nand_62_nl), or_11_cse);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_and_cse = core_wen & (~ and_dcpl_78)
      & (~ mux_615_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_or_15_cse
      = and_dcpl_784 | and_dcpl_785;
  assign nor_1493_cse = ~((~ main_stage_v_8) | (cfg_precision_1_sva_st_85!=2'b10));
  assign and_3293_nl = (~(inp_lookup_1_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp
      & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_12_1_1 & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_12_0_1
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_21==4'b1111))) & nor_tmp_161;
  assign mux_616_nl = MUX_s_1_2_2((and_3293_nl), nor_tmp_161, IsNaN_6U_10U_IsNaN_6U_10U_nor_tmp);
  assign nor_1491_nl = ~((~ (cfg_precision_1_sva_st_84[1])) | (~ main_stage_v_7)
      | (cfg_precision_1_sva_st_84[0]) | (mux_616_nl));
  assign nor_1492_nl = ~((chn_inp_in_crt_sva_8_739_736_1[0]) | (~ main_stage_v_8)
      | (cfg_precision_1_sva_st_85!=2'b10));
  assign mux_617_nl = MUX_s_1_2_2(nor_1493_cse, (nor_1492_nl), reg_FpMul_6U_10U_lor_3_lpi_1_dfm_3_cse);
  assign mux_618_nl = MUX_s_1_2_2(nor_1493_cse, (mux_617_nl), or_2797_cse);
  assign mux_619_nl = MUX_s_1_2_2((mux_618_nl), (nor_1491_nl), or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_12_cse = core_wen & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_or_15_cse
      & (mux_619_nl);
  assign nor_1490_cse = ~(reg_FpMul_6U_10U_lor_3_lpi_1_dfm_3_cse | (~ (chn_inp_in_crt_sva_8_739_736_1[0]))
      | (cfg_precision_1_sva_st_85!=2'b10) | (~ main_stage_v_8));
  assign mux_621_nl = MUX_s_1_2_2(or_tmp_1255, or_tmp_1058, or_11_cse);
  assign FpMul_6U_10U_oelse_and_cse = core_wen & (~ and_dcpl_78) & (~ (mux_621_nl));
  assign mux_622_nl = MUX_s_1_2_2(main_stage_v_8, main_stage_v_7, or_11_cse);
  assign cfg_precision_and_28_cse = core_wen & (~ and_dcpl_78) & (mux_622_nl);
  assign and_1270_rgt = (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_21==4'b1111)
      & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_12_0_1 & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_12_1_1
      & inp_lookup_1_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp
      & (~ IsNaN_6U_10U_IsNaN_6U_10U_nor_tmp) & (chn_inp_in_crt_sva_7_739_736_1[0])
      & or_11_cse;
  assign and_1273_rgt = ((FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_21!=4'b1111)
      | (~(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_12_0_1 & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_12_1_1
      & inp_lookup_1_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp)))
      & and_dcpl_798;
  assign and_1277_rgt = or_11_cse & (~ IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_19) & and_dcpl_801;
  assign and_1279_rgt = or_11_cse & IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_19 & and_dcpl_801;
  assign and_1280_rgt = ((chn_inp_in_crt_sva_7_739_736_1[0]) | IsNaN_6U_10U_8_land_1_lpi_1_dfm_7
      | IsNaN_6U_10U_9_land_1_lpi_1_dfm_8) & or_11_cse;
  assign nor_1488_cse = ~(reg_FpMul_6U_10U_lor_4_lpi_1_dfm_3_cse | (~ main_stage_v_8)
      | (~ (chn_inp_in_crt_sva_8_739_736_1[1])) | (cfg_precision_1_sva_st_85!=2'b10));
  assign nor_1486_nl = ~((cfg_precision_1_sva_st_84[0]) | (~((cfg_precision_1_sva_st_84[1])
      & (chn_inp_in_crt_sva_7_739_736_1[1]) & main_stage_v_7 & (IsNaN_6U_10U_IsNaN_6U_10U_nor_1_tmp
      | (~ FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_2_tmp)))));
  assign or_1284_nl = (~ reg_FpMul_6U_10U_lor_4_lpi_1_dfm_3_cse) | IsNaN_6U_10U_land_2_lpi_1_dfm_5;
  assign mux_624_nl = MUX_s_1_2_2(nor_1488_cse, and_3374_cse, or_1284_nl);
  assign mux_625_nl = MUX_s_1_2_2((mux_624_nl), (nor_1486_nl), or_11_cse);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_and_2_cse = core_wen & (~ and_dcpl_78)
      & (mux_625_nl);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_or_14_cse
      = and_dcpl_807 | and_dcpl_808;
  assign and_3291_nl = (~(inp_lookup_2_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp
      & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_12_1_1 & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_12_0_1
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_21==4'b1111))) & nor_tmp_166;
  assign mux_626_nl = MUX_s_1_2_2((and_3291_nl), nor_tmp_166, IsNaN_6U_10U_IsNaN_6U_10U_nor_1_tmp);
  assign nor_1482_nl = ~((cfg_precision_1_sva_st_84!=2'b10) | (~ main_stage_v_7)
      | (mux_626_nl));
  assign nor_1483_nl = ~((chn_inp_in_crt_sva_8_739_736_1[1]) | (~ main_stage_v_8)
      | (cfg_precision_1_sva_st_85!=2'b10));
  assign mux_627_nl = MUX_s_1_2_2(nor_1493_cse, (nor_1483_nl), reg_FpMul_6U_10U_lor_4_lpi_1_dfm_3_cse);
  assign mux_628_nl = MUX_s_1_2_2(nor_1493_cse, (mux_627_nl), or_2810_cse);
  assign mux_629_nl = MUX_s_1_2_2((mux_628_nl), (nor_1482_nl), or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_13_cse = core_wen & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_or_14_cse
      & (mux_629_nl);
  assign mux_631_nl = MUX_s_1_2_2(or_tmp_1302, or_tmp_1106, or_11_cse);
  assign FpMul_6U_10U_oelse_and_2_cse = core_wen & (~ and_dcpl_78) & (~ (mux_631_nl));
  assign and_1293_rgt = (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_21==4'b1111)
      & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_12_0_1 & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_12_1_1
      & inp_lookup_2_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp
      & (chn_inp_in_crt_sva_7_739_736_1[1]) & (~ IsNaN_6U_10U_IsNaN_6U_10U_nor_1_tmp)
      & or_11_cse;
  assign and_1296_rgt = ((FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_21!=4'b1111)
      | (~(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_12_0_1 & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_12_1_1
      & inp_lookup_2_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp)))
      & and_dcpl_821;
  assign nor_1733_rgt = ~((~ and_dcpl_825) | (chn_inp_in_crt_sva_7_739_736_1[1])
      | IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_5 | IsNaN_6U_10U_9_land_2_lpi_1_dfm_8);
  assign and_1303_rgt = and_dcpl_825 & (~ (chn_inp_in_crt_sva_7_739_736_1[1])) &
      IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_5 & (~ IsNaN_6U_10U_9_land_2_lpi_1_dfm_8);
  assign and_1304_rgt = (IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_19 | (chn_inp_in_crt_sva_7_739_736_1[1])
      | IsNaN_6U_10U_9_land_2_lpi_1_dfm_8) & or_11_cse;
  assign nand_561_nl = ~((IsNaN_6U_10U_IsNaN_6U_10U_nor_2_tmp | (~ FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_4_tmp))
      & (chn_inp_in_crt_sva_7_739_736_1[2]) & (cfg_precision_1_sva_st_84==2'b10)
      & main_stage_v_7);
  assign mux_634_nl = MUX_s_1_2_2(or_tmp_1312, or_tmp_1310, reg_FpMul_6U_10U_lor_5_lpi_1_dfm_3_cse);
  assign mux_635_cse = MUX_s_1_2_2((mux_634_nl), (nand_561_nl), or_11_cse);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_and_4_cse = core_wen & (~ and_dcpl_78)
      & (~ mux_635_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_or_13_cse
      = and_dcpl_831 | and_dcpl_832;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_14_cse = core_wen & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_or_13_cse
      & not_tmp_546;
  assign mux_641_nl = MUX_s_1_2_2(or_tmp_1312, or_tmp_1151, or_11_cse);
  assign FpMul_6U_10U_oelse_and_4_cse = core_wen & (~ and_dcpl_78) & (~ (mux_641_nl));
  assign and_1317_rgt = (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_21==4'b1111)
      & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_12_0_1 & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_12_1_1
      & inp_lookup_3_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp
      & (chn_inp_in_crt_sva_7_739_736_1[2]) & (~ IsNaN_6U_10U_IsNaN_6U_10U_nor_2_tmp)
      & or_11_cse;
  assign and_1320_rgt = ((FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_21!=4'b1111)
      | (~(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_12_0_1 & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_12_1_1
      & inp_lookup_3_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp)))
      & and_dcpl_845;
  assign nor_1732_rgt = ~(IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_19 | IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_5
      | (chn_inp_in_crt_sva_7_739_736_1[2]) | (~ and_dcpl_847));
  assign and_1327_rgt = (~ IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_19) & IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_5
      & (~ (chn_inp_in_crt_sva_7_739_736_1[2])) & and_dcpl_847;
  assign and_1329_rgt = FpAdd_6U_10U_1_or_16_cse & (~ (chn_inp_in_crt_sva_7_739_736_1[2]))
      & or_11_cse;
  assign nand_560_nl = ~((IsNaN_6U_10U_IsNaN_6U_10U_nor_3_tmp | (~ FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_6_tmp))
      & (chn_inp_in_crt_sva_7_739_736_1[3]) & (cfg_precision_1_sva_st_84==2'b10)
      & main_stage_v_7);
  assign mux_644_nl = MUX_s_1_2_2(or_tmp_1340, or_tmp_1338, reg_FpMul_6U_10U_lor_lpi_1_dfm_3_cse);
  assign mux_645_cse = MUX_s_1_2_2((mux_644_nl), (nand_560_nl), or_11_cse);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_and_6_cse = core_wen & (~ and_dcpl_78)
      & (~ mux_645_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_or_12_cse
      = and_dcpl_856 | and_dcpl_857;
  assign and_3287_nl = (~(inp_lookup_4_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp
      & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_12_1_1 & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_12_0_1
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_21==4'b1111))) & nor_tmp_176;
  assign mux_646_nl = MUX_s_1_2_2((and_3287_nl), nor_tmp_176, IsNaN_6U_10U_IsNaN_6U_10U_nor_3_tmp);
  assign nor_1470_nl = ~((~ (cfg_precision_1_sva_st_84[1])) | (~ main_stage_v_7)
      | (cfg_precision_1_sva_st_84[0]) | (mux_646_nl));
  assign nor_1471_nl = ~((chn_inp_in_crt_sva_8_739_736_1[3]) | (~ main_stage_v_8)
      | (cfg_precision_1_sva_st_85!=2'b10));
  assign mux_647_nl = MUX_s_1_2_2(nor_1493_cse, (nor_1471_nl), reg_FpMul_6U_10U_lor_lpi_1_dfm_3_cse);
  assign mux_648_nl = MUX_s_1_2_2(nor_1493_cse, (mux_647_nl), or_2822_cse);
  assign mux_649_nl = MUX_s_1_2_2((mux_648_nl), (nor_1470_nl), or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_15_cse = core_wen & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_or_12_cse
      & (mux_649_nl);
  assign nor_1469_cse = ~(reg_FpMul_6U_10U_lor_lpi_1_dfm_3_cse | (~ (chn_inp_in_crt_sva_8_739_736_1[3]))
      | (cfg_precision_1_sva_st_85!=2'b10) | (~ main_stage_v_8));
  assign mux_651_nl = MUX_s_1_2_2(or_tmp_1340, or_tmp_1198, or_11_cse);
  assign FpMul_6U_10U_oelse_and_6_cse = core_wen & (~ and_dcpl_78) & (~ (mux_651_nl));
  assign and_1342_rgt = (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_21==4'b1111)
      & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_12_0_1 & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_12_1_1
      & inp_lookup_4_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp
      & (chn_inp_in_crt_sva_7_739_736_1[3]) & (~ IsNaN_6U_10U_IsNaN_6U_10U_nor_3_tmp)
      & or_11_cse;
  assign and_1345_rgt = ((FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_21!=4'b1111)
      | (~(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_12_0_1 & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_12_1_1
      & inp_lookup_4_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp)))
      & and_dcpl_870;
  assign and_1349_rgt = and_dcpl_874 & and_dcpl_872 & (~ IsNaN_6U_10U_8_land_lpi_1_dfm_st_5);
  assign and_1351_rgt = and_dcpl_874 & and_dcpl_872 & IsNaN_6U_10U_8_land_lpi_1_dfm_st_5;
  assign and_1352_rgt = (FpAdd_6U_10U_1_or_18_cse | (chn_inp_in_crt_sva_7_739_736_1[3]))
      & or_11_cse;
  assign IsNaN_6U_10U_2_aelse_and_cse = core_wen & (~ and_dcpl_78) & (~ mux_659_itm);
  assign and_1360_rgt = (inp_lookup_1_FpMul_6U_10U_oelse_1_acc_itm_7_1 | reg_FpMul_6U_10U_lor_3_lpi_1_dfm_3_cse
      | (~ inp_lookup_1_FpMul_6U_10U_else_2_if_acc_itm_6_1)) & or_11_cse;
  assign and_3286_cse = (chn_inp_in_crt_sva_8_739_736_1[0]) & main_stage_v_8;
  assign mux_660_nl = MUX_s_1_2_2(and_3113_cse, and_3286_cse, or_11_cse);
  assign cfg_precision_and_32_cse = core_wen & (~ and_dcpl_78) & (mux_660_nl);
  assign IsNaN_6U_10U_2_aelse_and_1_cse = core_wen & (~ and_dcpl_78) & (~ mux_666_itm);
  assign and_1364_rgt = (inp_lookup_2_FpMul_6U_10U_oelse_1_acc_itm_7_1 | reg_FpMul_6U_10U_lor_4_lpi_1_dfm_3_cse
      | (~ inp_lookup_2_FpMul_6U_10U_else_2_if_acc_itm_6_1)) & or_11_cse;
  assign and_3285_cse = (chn_inp_in_crt_sva_8_739_736_1[1]) & main_stage_v_8;
  assign mux_667_nl = MUX_s_1_2_2(and_3111_cse, and_3285_cse, or_11_cse);
  assign cfg_precision_and_33_cse = core_wen & (~ and_dcpl_78) & (mux_667_nl);
  assign IsNaN_6U_10U_2_aelse_and_2_cse = core_wen & (~ and_dcpl_78) & (~ mux_673_itm);
  assign and_1368_rgt = (inp_lookup_3_FpMul_6U_10U_oelse_1_acc_itm_7_1 | reg_FpMul_6U_10U_lor_5_lpi_1_dfm_3_cse
      | (~ inp_lookup_3_FpMul_6U_10U_else_2_if_acc_itm_6_1)) & or_11_cse;
  assign and_3283_cse = (chn_inp_in_crt_sva_8_739_736_1[2]) & main_stage_v_8;
  assign mux_674_nl = MUX_s_1_2_2(and_3110_cse, and_3283_cse, or_11_cse);
  assign cfg_precision_and_34_cse = core_wen & (~ and_dcpl_78) & (mux_674_nl);
  assign IsNaN_6U_10U_2_aelse_and_3_cse = core_wen & (~ and_dcpl_78) & (~ mux_680_itm);
  assign and_1372_rgt = (inp_lookup_4_FpMul_6U_10U_oelse_1_acc_itm_7_1 | reg_FpMul_6U_10U_lor_lpi_1_dfm_3_cse
      | (~ inp_lookup_4_FpMul_6U_10U_else_2_if_acc_itm_6_1)) & or_11_cse;
  assign and_3281_cse = (chn_inp_in_crt_sva_8_739_736_1[3]) & main_stage_v_8;
  assign mux_681_nl = MUX_s_1_2_2(and_3112_cse, and_3281_cse, or_11_cse);
  assign cfg_precision_and_35_cse = core_wen & (~ and_dcpl_78) & (mux_681_nl);
  assign mux_682_nl = MUX_s_1_2_2(main_stage_v_9, main_stage_v_8, or_11_cse);
  assign chn_inp_in_flow_and_32_cse = core_wen & (~ and_dcpl_78) & (mux_682_nl);
  assign nand_653_cse = ~(main_stage_v_10 & (cfg_precision_1_sva_st_87[1]));
  assign and_4178_cse = main_stage_v_9 & (chn_inp_in_crt_sva_9_739_736_1[0]) & (cfg_precision_1_sva_st_86==2'b10);
  assign and_4207_nl = main_stage_v_10 & (chn_inp_in_crt_sva_10_739_736_1[0]) & (cfg_precision_1_sva_st_87==2'b10);
  assign mux_685_nl = MUX_s_1_2_2((and_4207_nl), and_4178_cse, or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_5_cse = core_wen & (~ and_dcpl_78)
      & (mux_685_nl);
  assign nor_1435_nl = ~((cfg_precision_1_sva_st_87[0]) | (~((chn_inp_in_crt_sva_10_739_736_1[0])
      & main_stage_v_10 & (cfg_precision_1_sva_st_87[1]))));
  assign mux_690_nl = MUX_s_1_2_2((nor_1435_nl), and_4178_cse, or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_cse = core_wen & (~ and_dcpl_78)
      & (mux_690_nl);
  assign nand_776_nl = ~(main_stage_v_10 & (chn_inp_in_crt_sva_10_739_736_1[0]) &
      (cfg_precision_1_sva_st_87==2'b10));
  assign mux_698_nl = MUX_s_1_2_2((nand_776_nl), or_tmp_1389, or_11_cse);
  assign FpMul_6U_10U_o_expo_and_8_cse = core_wen & (~ and_dcpl_78) & (~ (mux_698_nl));
  assign mux_699_nl = MUX_s_1_2_2(or_tmp_1502, or_tmp_1389, or_11_cse);
  assign FpAdd_6U_10U_is_a_greater_and_cse = core_wen & (~ and_dcpl_78) & (~ (mux_699_nl));
  assign nand_652_cse = ~(main_stage_v_10 & (cfg_precision_1_sva_st_101[1]));
  assign and_4177_cse = main_stage_v_9 & (chn_inp_in_crt_sva_9_739_736_1[1]) & (cfg_precision_1_sva_st_100==2'b10);
  assign and_4206_nl = main_stage_v_10 & (chn_inp_in_crt_sva_10_739_736_1[1]) & (cfg_precision_1_sva_st_101==2'b10);
  assign mux_703_nl = MUX_s_1_2_2((and_4206_nl), and_4177_cse, or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_6_cse = core_wen & (~ and_dcpl_78)
      & (mux_703_nl);
  assign nor_1430_nl = ~((~ (chn_inp_in_crt_sva_10_739_736_1[1])) | (cfg_precision_1_sva_st_101[0])
      | nand_652_cse);
  assign mux_708_nl = MUX_s_1_2_2((nor_1430_nl), and_4177_cse, or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_13_cse = core_wen & (~ and_dcpl_78)
      & (mux_708_nl);
  assign nand_775_nl = ~(main_stage_v_10 & (chn_inp_in_crt_sva_10_739_736_1[1]) &
      (cfg_precision_1_sva_st_101==2'b10));
  assign mux_716_nl = MUX_s_1_2_2((nand_775_nl), or_tmp_1418, or_11_cse);
  assign FpMul_6U_10U_o_expo_and_10_cse = core_wen & (~ and_dcpl_78) & (~ (mux_716_nl));
  assign mux_717_nl = MUX_s_1_2_2(or_tmp_1537, or_tmp_1418, or_11_cse);
  assign FpAdd_6U_10U_is_a_greater_and_2_cse = core_wen & (~ and_dcpl_78) & (~ (mux_717_nl));
  assign and_4176_cse = main_stage_v_9 & (chn_inp_in_crt_sva_9_739_736_1[2]) & (cfg_precision_1_sva_st_112==2'b10);
  assign and_4205_nl = main_stage_v_10 & (chn_inp_in_crt_sva_10_739_736_1[2]) & (cfg_precision_1_sva_st_113==2'b10);
  assign mux_721_nl = MUX_s_1_2_2((and_4205_nl), and_4176_cse, or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_7_cse = core_wen & (~ and_dcpl_78)
      & (mux_721_nl);
  assign nor_1425_nl = ~((~ (chn_inp_in_crt_sva_10_739_736_1[2])) | (cfg_precision_1_sva_st_113[0])
      | (~(main_stage_v_10 & (cfg_precision_1_sva_st_113[1]))));
  assign mux_726_nl = MUX_s_1_2_2((nor_1425_nl), and_4176_cse, or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_15_cse = core_wen & (~ and_dcpl_78)
      & (mux_726_nl);
  assign nand_774_cse = ~(main_stage_v_10 & (chn_inp_in_crt_sva_10_739_736_1[2])
      & (cfg_precision_1_sva_st_113==2'b10));
  assign mux_734_nl = MUX_s_1_2_2(nand_774_cse, or_tmp_1444, or_11_cse);
  assign FpMul_6U_10U_o_expo_and_12_cse = core_wen & (~ and_dcpl_78) & (~ (mux_734_nl));
  assign and_4175_cse = main_stage_v_9 & (chn_inp_in_crt_sva_9_739_736_1[3]) & (cfg_precision_1_sva_st_124==2'b10);
  assign and_4204_nl = main_stage_v_10 & (chn_inp_in_crt_sva_10_739_736_1[3]) & (cfg_precision_1_sva_st_125==2'b10);
  assign mux_739_nl = MUX_s_1_2_2((and_4204_nl), and_4175_cse, or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_8_cse = core_wen & (~ and_dcpl_78)
      & (mux_739_nl);
  assign nor_1420_nl = ~((~ (chn_inp_in_crt_sva_10_739_736_1[3])) | (cfg_precision_1_sva_st_125[0])
      | (~(main_stage_v_10 & (cfg_precision_1_sva_st_125[1]))));
  assign mux_744_nl = MUX_s_1_2_2((nor_1420_nl), and_4175_cse, or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_17_cse = core_wen & (~ and_dcpl_78)
      & (mux_744_nl);
  assign nand_773_cse = ~(main_stage_v_10 & (chn_inp_in_crt_sva_10_739_736_1[3])
      & (cfg_precision_1_sva_st_125==2'b10));
  assign mux_752_nl = MUX_s_1_2_2(nand_773_cse, or_tmp_1467, or_11_cse);
  assign FpMul_6U_10U_o_expo_and_14_cse = core_wen & (~ and_dcpl_78) & (~ (mux_752_nl));
  assign mux_755_nl = MUX_s_1_2_2(main_stage_v_10, main_stage_v_9, or_11_cse);
  assign chn_inp_in_flow_and_36_cse = core_wen & (~ and_dcpl_78) & (mux_755_nl);
  assign mux_756_nl = MUX_s_1_2_2(or_1621_cse, or_tmp_1502, or_11_cse);
  assign FpAdd_6U_10U_is_addition_and_cse = core_wen & (~ and_dcpl_78) & (~ (mux_756_nl));
  assign or_1621_cse = (~ (chn_inp_in_crt_sva_11_739_736_1[0])) | (cfg_precision_1_sva_st_88[0])
      | not_tmp_698;
  assign mux_761_nl = MUX_s_1_2_2(or_1632_cse, or_tmp_1537, or_11_cse);
  assign FpAdd_6U_10U_is_addition_and_2_cse = core_wen & (~ and_dcpl_78) & (~ (mux_761_nl));
  assign or_1632_cse = (~ (chn_inp_in_crt_sva_11_739_736_1[1])) | (cfg_precision_1_sva_st_102[0])
      | not_tmp_703;
  assign mux_766_nl = MUX_s_1_2_2(or_1645_cse, nand_774_cse, or_11_cse);
  assign FpAdd_6U_10U_is_addition_and_4_cse = core_wen & (~ and_dcpl_78) & (~ (mux_766_nl));
  assign or_1645_cse = (~ (chn_inp_in_crt_sva_11_739_736_1[2])) | (cfg_precision_1_sva_st_114[0])
      | not_tmp_708;
  assign mux_771_nl = MUX_s_1_2_2(or_1658_cse, nand_773_cse, or_11_cse);
  assign FpAdd_6U_10U_is_addition_and_6_cse = core_wen & (~ and_dcpl_78) & (~ (mux_771_nl));
  assign or_1658_cse = (~ (chn_inp_in_crt_sva_11_739_736_1[3])) | (cfg_precision_1_sva_st_126[0])
      | not_tmp_711;
  assign chn_inp_in_flow_and_40_cse = core_wen & (~ and_dcpl_78) & mux_tmp_698;
  assign IsInf_6U_23U_aelse_and_cse = core_wen & (~(or_dcpl_264 | (~ main_stage_v_12)
      | and_dcpl_78 | (~ (chn_inp_in_crt_sva_12_739_736_1[0]))));
  assign nand_491_nl = ~((~((~(FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_1_sva_st_2
      & inp_lookup_1_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2)) & FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_1_sva_2))
      & main_stage_v_12 & (chn_inp_in_crt_sva_12_739_736_1[0]) & (cfg_precision_1_sva_st_89==2'b10));
  assign mux_777_nl = MUX_s_1_2_2((nand_491_nl), or_tmp_1661, or_11_cse);
  assign or_5699_nl = nor_1896_cse | or_tmp_1661;
  assign mux_778_nl = MUX_s_1_2_2(or_tmp_1665, or_tmp_1661, or_11_cse);
  assign mux_779_nl = MUX_s_1_2_2((mux_778_nl), (or_5699_nl), reg_FpNormalize_6U_23U_lor_1_lpi_1_dfm_4_cse);
  assign mux_780_nl = MUX_s_1_2_2((mux_779_nl), (mux_777_nl), FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_4[23]);
  assign FpAdd_6U_10U_and_43_cse = core_wen & (~ and_dcpl_78) & (~ (mux_780_nl));
  assign and_1386_rgt = or_11_cse & (~ reg_inp_lookup_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse);
  assign IsNaN_6U_10U_3_aelse_and_cse = core_wen & (~ and_dcpl_78) & (~ mux_782_itm);
  assign mux_789_nl = MUX_s_1_2_2(or_tmp_1690, or_tmp_1671, IsNaN_6U_10U_3_land_1_lpi_1_dfm_8);
  assign mux_790_nl = MUX_s_1_2_2((mux_789_nl), or_tmp_1687, or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_19_cse = core_wen & (~ and_dcpl_78)
      & (~ (mux_790_nl));
  assign IsInf_6U_23U_aelse_and_1_cse = core_wen & (~(or_dcpl_269 | or_dcpl_4));
  assign or_1697_nl = (~(FpAdd_6U_10U_mux_18_tmp_23 | (~ FpNormalize_6U_23U_if_FpNormalize_6U_23U_if_nand_1_tmp)))
      | (~ (chn_inp_in_crt_sva_11_739_736_1[1])) | (cfg_precision_1_sva_st_102[0])
      | not_tmp_703;
  assign mux_792_nl = MUX_s_1_2_2(or_tmp_1699, or_tmp_1697, FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_4[23]);
  assign mux_794_nl = MUX_s_1_2_2(mux_tmp_715, (mux_792_nl), FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_2_sva_2);
  assign or_1705_nl = (FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_4[23]) | inp_lookup_2_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2
      | (~ main_stage_v_12) | reg_FpNormalize_6U_23U_lor_2_lpi_1_dfm_4_cse | (~ (chn_inp_in_crt_sva_12_739_736_1[1]))
      | (cfg_precision_1_sva_st_103!=2'b10);
  assign mux_795_nl = MUX_s_1_2_2(mux_tmp_715, (or_1705_nl), FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_2_sva_2);
  assign mux_796_nl = MUX_s_1_2_2((mux_795_nl), (mux_794_nl), FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_2_sva_st_2);
  assign mux_797_nl = MUX_s_1_2_2((mux_796_nl), (or_1697_nl), or_11_cse);
  assign FpAdd_6U_10U_and_45_cse = core_wen & (~ and_dcpl_78) & (~ (mux_797_nl));
  assign and_1388_rgt = or_11_cse & (~ reg_inp_lookup_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse);
  assign IsNaN_6U_10U_3_aelse_and_1_cse = core_wen & (~ and_dcpl_78) & (~ mux_799_itm);
  assign nor_1407_cse = ~((~ main_stage_v_11) | (~ (chn_inp_in_crt_sva_11_739_736_1[1]))
      | (cfg_precision_1_sva_st_102[0]) | (~((cfg_precision_1_sva_st_102[1]) & ((~(IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_23
      | (~ IsNaN_6U_10U_3_land_2_lpi_1_dfm_7))) | IsNaN_6U_10U_2_land_2_lpi_1_dfm_25))));
  assign mux_803_nl = MUX_s_1_2_2(or_tmp_1728, or_1632_cse, or_11_cse);
  assign or_1732_nl = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | or_tmp_1728;
  assign mux_804_nl = MUX_s_1_2_2((or_1732_nl), (mux_803_nl), or_tmp_1724);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_21_cse = core_wen & (~ and_dcpl_78)
      & (~ (mux_804_nl));
  assign IsInf_6U_23U_aelse_and_2_cse = core_wen & (~((~ main_stage_v_12) | (~ (chn_inp_in_crt_sva_12_739_736_1[2]))
      | (~ (cfg_precision_1_sva_st_115[1])) | and_dcpl_78 | (cfg_precision_1_sva_st_115[0])));
  assign nand_88_nl = ~((FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_4[23]) & (~ or_tmp_1736));
  assign or_1740_nl = (~ (FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_4[23])) | FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_3_sva_2
      | (cfg_precision_1_sva_st_115[0]) | not_tmp_733;
  assign mux_806_nl = MUX_s_1_2_2((or_1740_nl), (nand_88_nl), FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_3_sva_st_2);
  assign mux_807_nl = MUX_s_1_2_2((mux_806_nl), or_tmp_1734, or_11_cse);
  assign mux_808_nl = MUX_s_1_2_2(or_tmp_1741, or_tmp_1736, FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_4[23]);
  assign or_1745_nl = FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_3_sva_2
      | (cfg_precision_1_sva_st_115[0]) | not_tmp_733;
  assign mux_810_nl = MUX_s_1_2_2(or_tmp_1741, (or_1745_nl), FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_4[23]);
  assign mux_812_nl = MUX_s_1_2_2((mux_810_nl), (mux_808_nl), FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_3_sva_st_2);
  assign mux_813_nl = MUX_s_1_2_2((mux_812_nl), or_tmp_1734, or_11_cse);
  assign mux_814_nl = MUX_s_1_2_2((mux_813_nl), (mux_807_nl), FpNormalize_6U_23U_lor_3_lpi_1_dfm_5);
  assign FpAdd_6U_10U_and_47_cse = core_wen & (~ and_dcpl_78) & (~ (mux_814_nl));
  assign and_1390_rgt = or_11_cse & (~ reg_inp_lookup_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse);
  assign IsNaN_6U_10U_3_aelse_and_2_cse = core_wen & (~ and_dcpl_78) & (~ mux_816_itm);
  assign nor_1397_cse = ~((~ main_stage_v_11) | (~ (chn_inp_in_crt_sva_11_739_736_1[2]))
      | (cfg_precision_1_sva_st_114[0]) | (~((cfg_precision_1_sva_st_114[1]) & ((~(IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_23
      | (~ IsNaN_6U_10U_3_land_3_lpi_1_dfm_7))) | IsNaN_6U_10U_2_land_3_lpi_1_dfm_25))));
  assign mux_821_nl = MUX_s_1_2_2(or_tmp_1774, or_1645_cse, or_11_cse);
  assign or_1778_nl = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | or_tmp_1774;
  assign mux_822_nl = MUX_s_1_2_2((or_1778_nl), (mux_821_nl), or_tmp_1770);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_23_cse = core_wen & (~ and_dcpl_78)
      & (~ (mux_822_nl));
  assign IsInf_6U_23U_aelse_and_3_cse = core_wen & (~(or_dcpl_278 | or_dcpl_4));
  assign or_1782_nl = (~(FpAdd_6U_10U_mux_50_tmp_23 | (~ FpNormalize_6U_23U_if_FpNormalize_6U_23U_if_nand_3_tmp)))
      | (~ (chn_inp_in_crt_sva_11_739_736_1[3])) | (cfg_precision_1_sva_st_126[0])
      | not_tmp_711;
  assign nand_667_nl = ~(inp_lookup_4_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2
      & FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_sva_st_2 & main_stage_v_12
      & (chn_inp_in_crt_sva_12_739_736_1[3]) & (cfg_precision_1_sva_st_127==2'b10));
  assign mux_824_nl = MUX_s_1_2_2(or_tmp_1784, (nand_667_nl), FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_4[23]);
  assign mux_825_nl = MUX_s_1_2_2(or_tmp_1784, or_tmp_1786, FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_4[23]);
  assign mux_826_nl = MUX_s_1_2_2((mux_825_nl), (mux_824_nl), FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_sva_2);
  assign mux_827_nl = MUX_s_1_2_2((mux_826_nl), (or_1782_nl), or_11_cse);
  assign FpAdd_6U_10U_and_49_cse = core_wen & (~ and_dcpl_78) & (~ (mux_827_nl));
  assign and_1392_rgt = or_11_cse & (~ reg_inp_lookup_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse);
  assign IsNaN_6U_10U_3_aelse_and_3_cse = core_wen & (~ and_dcpl_78) & (~ mux_829_itm);
  assign nand_664_nl = ~(FpAdd_6U_10U_or_19_cse & main_stage_v_12 & (chn_inp_in_crt_sva_12_739_736_1[3])
      & (cfg_precision_1_sva_st_127==2'b10));
  assign mux_834_nl = MUX_s_1_2_2((nand_664_nl), or_tmp_1806, or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_25_cse = core_wen & (~ and_dcpl_78)
      & (~ (mux_834_nl));
  assign mux_836_nl = MUX_s_1_2_2(main_stage_v_12, main_stage_v_11, or_11_cse);
  assign inp_lookup_and_cse = core_wen & (~ and_dcpl_78) & (mux_836_nl);
  assign or_1826_nl = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (chn_inp_in_crt_sva_12_739_736_1[3]) | inp_lookup_else_unequal_tmp_38 | (~
      main_stage_v_12);
  assign or_1830_nl = (chn_inp_in_crt_sva_12_739_736_1[3]) | inp_lookup_else_unequal_tmp_38
      | (~ main_stage_v_12);
  assign mux_840_nl = MUX_s_1_2_2((or_1830_nl), or_tmp_1826, or_11_cse);
  assign mux_841_nl = MUX_s_1_2_2((mux_840_nl), (or_1826_nl), inp_lookup_else_unequal_tmp_37);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_and_cse = core_wen & (~ and_dcpl_78)
      & (~ (mux_841_nl));
  assign or_1837_nl = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | inp_lookup_else_unequal_tmp_38 | (chn_inp_in_crt_sva_12_739_736_1[0]) | (~
      main_stage_v_12);
  assign or_1840_nl = inp_lookup_else_unequal_tmp_38 | (chn_inp_in_crt_sva_12_739_736_1[0])
      | (~ main_stage_v_12);
  assign mux_845_nl = MUX_s_1_2_2((or_1840_nl), or_tmp_1818, or_11_cse);
  assign mux_846_nl = MUX_s_1_2_2((mux_845_nl), (or_1837_nl), inp_lookup_else_unequal_tmp_37);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_cse = core_wen & (~ and_dcpl_78) &
      (~ (mux_846_nl));
  assign or_1849_nl = (chn_inp_in_crt_sva_12_739_736_1[2]) | inp_lookup_else_unequal_tmp_38
      | (~ main_stage_v_12);
  assign mux_849_nl = MUX_s_1_2_2((or_1849_nl), or_tmp_1845, or_11_cse);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_and_6_cse = core_wen & (~ and_dcpl_78)
      & (~ (mux_849_nl));
  assign or_1860_nl = inp_lookup_else_unequal_tmp_38 | (chn_inp_in_crt_sva_12_739_736_1[1])
      | (~ main_stage_v_12);
  assign mux_853_nl = MUX_s_1_2_2((or_1860_nl), or_tmp_1856, or_11_cse);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_2_cse = core_wen & (~ and_dcpl_78)
      & (~ (mux_853_nl));
  assign FpAdd_6U_10U_and_51_cse = core_wen & (and_dcpl_930 | and_dcpl_935 | and_dcpl_936)
      & mux_tmp_698;
  assign FpAdd_6U_10U_and_53_cse = core_wen & (and_dcpl_940 | and_dcpl_944 | and_dcpl_945)
      & mux_tmp_698;
  assign FpAdd_6U_10U_and_55_cse = core_wen & (and_dcpl_949 | and_dcpl_954 | and_dcpl_955)
      & mux_tmp_698;
  assign FpAdd_6U_10U_and_57_cse = core_wen & (and_dcpl_959 | and_dcpl_961 | and_dcpl_962)
      & mux_tmp_698;
  assign mux_854_cse = MUX_s_1_2_2(or_tmp_1182, or_tmp_959, or_11_cse);
  assign IsNaN_6U_10U_8_aelse_and_3_cse = core_wen & FpNormalize_6U_23U_1_if_FpNormalize_6U_23U_1_if_or_3_cse
      & (~ mux_854_cse);
  assign nor_1380_cse = ~((~ main_stage_v_1) | (cfg_precision_1_sva_st_90!=2'b10)
      | (chn_inp_in_crt_sva_1_739_395_1[341]));
  assign nor_257_cse = ~((chn_inp_in_crt_sva_2_739_736_1[0]) | (cfg_precision_1_sva_st_91!=2'b10));
  assign and_1468_rgt = and_dcpl_423 & (~((chn_inp_in_crt_sva_2_739_736_1[0]) | IsNaN_6U_10U_7_land_1_lpi_1_dfm_5))
      & and_dcpl_419;
  assign and_1471_rgt = and_dcpl_423 & (~ (chn_inp_in_crt_sva_2_739_736_1[0])) &
      IsNaN_6U_10U_7_land_1_lpi_1_dfm_5 & and_dcpl_419;
  assign or_1889_nl = nor_35_cse | (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_7_1_1
      & FpAdd_8U_23U_o_sign_1_lpi_1_dfm_7 & inp_lookup_1_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_tmp
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_9==4'b1111) & (IsNaN_6U_10U_4_nor_tmp
      | (~(inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_5_1 & (inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_4_0_1==5'b11111)
      & IsNaN_8U_23U_land_1_lpi_1_dfm_st_4))));
  assign mux_866_nl = MUX_s_1_2_2(and_tmp_111, (or_1889_nl), or_11_cse);
  assign mux_867_nl = MUX_s_1_2_2(nand_tmp_91, (mux_866_nl), nor_257_cse);
  assign nor_1372_nl = ~((~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ and_tmp_111));
  assign mux_868_nl = MUX_s_1_2_2((nor_1372_nl), nand_tmp_91, or_683_cse);
  assign nor_1373_nl = ~((~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (main_stage_v_3 & (~ or_tmp_1891)));
  assign mux_869_nl = MUX_s_1_2_2((nor_1373_nl), nand_tmp_91, or_471_cse);
  assign mux_870_nl = MUX_s_1_2_2((mux_869_nl), (mux_868_nl), main_stage_v_1);
  assign mux_871_nl = MUX_s_1_2_2((mux_870_nl), (mux_867_nl), main_stage_v_2);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_31_cse = FpAdd_8U_23U_o_expo_and_cse
      & FpMul_6U_10U_2_else_2_else_if_FpMul_6U_10U_2_else_2_else_if_or_3_cse & (mux_871_nl);
  assign or_1927_nl = nor_584_cse | (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_7_1_1
      & FpAdd_8U_23U_o_sign_2_lpi_1_dfm_7 & inp_lookup_2_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_tmp
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_9==4'b1111) & (IsNaN_6U_10U_4_nor_1_tmp
      | (~(inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_6_5_1 & (inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_6_4_0_1==5'b11111)
      & IsNaN_8U_23U_land_2_lpi_1_dfm_st_4))));
  assign mux_883_nl = MUX_s_1_2_2(and_tmp_116, (or_1927_nl), or_11_cse);
  assign mux_884_nl = MUX_s_1_2_2(nand_tmp_95, (mux_883_nl), nor_266_cse);
  assign nor_1359_nl = ~((~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ and_tmp_116));
  assign mux_885_nl = MUX_s_1_2_2((nor_1359_nl), nand_tmp_95, or_740_cse);
  assign nor_1360_nl = ~((~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (main_stage_v_3 & (~ or_tmp_1929)));
  assign mux_886_nl = MUX_s_1_2_2((nor_1360_nl), nand_tmp_95, or_763_cse);
  assign mux_887_nl = MUX_s_1_2_2((mux_886_nl), (mux_885_nl), main_stage_v_1);
  assign mux_888_nl = MUX_s_1_2_2((mux_887_nl), (mux_884_nl), main_stage_v_2);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_33_cse = FpAdd_8U_23U_o_expo_and_cse
      & FpMul_6U_10U_2_else_2_else_if_FpMul_6U_10U_2_else_2_else_if_or_2_cse & (mux_888_nl);
  assign nor_1354_cse = ~((~ main_stage_v_1) | (cfg_precision_1_sva_st_90!=2'b10)
      | (chn_inp_in_crt_sva_1_739_395_1[343]));
  assign nor_275_cse = ~((chn_inp_in_crt_sva_2_739_736_1[2]) | (cfg_precision_1_sva_st_91!=2'b10));
  assign and_1474_rgt = and_dcpl_423 & (~ IsNaN_6U_10U_7_land_3_lpi_1_dfm_5) & main_stage_v_2
      & and_dcpl_524;
  assign and_1477_rgt = and_dcpl_423 & IsNaN_6U_10U_7_land_3_lpi_1_dfm_5 & main_stage_v_2
      & and_dcpl_524;
  assign or_1965_nl = nor_586_cse | (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_7_1_1
      & FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_7_0_1 & inp_lookup_4_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_tmp
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_9==4'b1111) & (IsNaN_6U_10U_4_nor_3_tmp
      | (~(inp_lookup_else_if_a0_15_10_lpi_1_dfm_6_5_1 & (inp_lookup_else_if_a0_15_10_lpi_1_dfm_6_4_0_1==5'b11111)
      & IsNaN_8U_23U_land_lpi_1_dfm_st_4))));
  assign mux_900_nl = MUX_s_1_2_2(and_tmp_121, (or_1965_nl), or_11_cse);
  assign nor_279_nl = ~((chn_inp_in_crt_sva_2_739_736_1[3]) | (cfg_precision_1_sva_st_91!=2'b10));
  assign mux_901_nl = MUX_s_1_2_2(nand_tmp_99, (mux_900_nl), nor_279_nl);
  assign nor_1346_nl = ~((~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ and_tmp_121));
  assign mux_902_nl = MUX_s_1_2_2((nor_1346_nl), nand_tmp_99, or_1970_cse);
  assign nor_1347_nl = ~((~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (main_stage_v_3 & (~ or_tmp_1967)));
  assign mux_903_nl = MUX_s_1_2_2((nor_1347_nl), nand_tmp_99, or_114_cse);
  assign mux_904_nl = MUX_s_1_2_2((mux_903_nl), (mux_902_nl), main_stage_v_1);
  assign mux_905_nl = MUX_s_1_2_2((mux_904_nl), (mux_901_nl), main_stage_v_2);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_37_cse = FpAdd_8U_23U_o_expo_and_cse
      & (and_dcpl_1009 | and_dcpl_1007) & (mux_905_nl);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_asn_FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_conc_10_cgspt_7_mux_nl
      = MUX_v_8_2_2((chn_inp_in_crt_sva_1_739_395_1[179:172]), (chn_inp_in_crt_sva_1_739_395_1[307:300]),
      and_dcpl_406);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_mux1h_4_itm = MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_8,
      ({2'b0 , (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_asn_FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_conc_10_cgspt_7_mux_nl)}),
      mux_tmp_1845);
  assign and_1537_rgt = and_dcpl_1060 & (cfg_precision_rsci_d[1]) & (~ (chn_inp_in_rsci_d_mxwt[736]))
      & (chn_inp_in_rsci_d_mxwt[342]) & (chn_inp_in_rsci_d_mxwt[343]) & (chn_inp_in_rsci_d_mxwt[344])
      & (chn_inp_in_rsci_d_mxwt[345]) & (chn_inp_in_rsci_d_mxwt[346]) & IsDenorm_5U_10U_3_or_tmp;
  assign and_1538_rgt = or_dcpl_499 & and_dcpl_144;
  assign and_1588_rgt = and_dcpl_1060 & (cfg_precision_rsci_d[1]) & (~ (chn_inp_in_rsci_d_mxwt[737]))
      & (chn_inp_in_rsci_d_mxwt[358]) & (chn_inp_in_rsci_d_mxwt[359]) & (chn_inp_in_rsci_d_mxwt[360])
      & (chn_inp_in_rsci_d_mxwt[361]) & (chn_inp_in_rsci_d_mxwt[362]) & IsDenorm_5U_10U_3_or_1_tmp;
  assign and_1589_rgt = or_dcpl_542 & and_dcpl_214;
  assign and_1639_rgt = and_dcpl_1060 & (cfg_precision_rsci_d[1]) & (~ (chn_inp_in_rsci_d_mxwt[738]))
      & (chn_inp_in_rsci_d_mxwt[374]) & (chn_inp_in_rsci_d_mxwt[375]) & (chn_inp_in_rsci_d_mxwt[376])
      & (chn_inp_in_rsci_d_mxwt[377]) & (chn_inp_in_rsci_d_mxwt[378]) & IsDenorm_5U_10U_3_or_2_tmp;
  assign and_1640_rgt = or_dcpl_585 & and_dcpl_284;
  assign and_1690_rgt = and_dcpl_1060 & (cfg_precision_rsci_d[1]) & (~ (chn_inp_in_rsci_d_mxwt[739]))
      & (chn_inp_in_rsci_d_mxwt[390]) & (chn_inp_in_rsci_d_mxwt[391]) & (chn_inp_in_rsci_d_mxwt[392])
      & (chn_inp_in_rsci_d_mxwt[393]) & (chn_inp_in_rsci_d_mxwt[394]) & IsDenorm_5U_10U_3_or_3_tmp;
  assign and_1691_rgt = or_dcpl_628 & and_dcpl_354;
  assign IntLeadZero_35U_1_leading_sign_35_0_rtn_and_cse = core_wen & (~(and_dcpl_173
      | or_dcpl_631 | (fsm_output[0])));
  assign IntLeadZero_35U_1_leading_sign_35_0_rtn_and_1_cse = core_wen & (~(and_dcpl_243
      | or_dcpl_634 | (fsm_output[0])));
  assign IntLeadZero_35U_1_leading_sign_35_0_rtn_and_2_cse = core_wen & (~(and_dcpl_313
      | or_dcpl_637 | (fsm_output[0])));
  assign IntLeadZero_35U_1_leading_sign_35_0_rtn_and_3_cse = core_wen & (~(and_dcpl_383
      | or_dcpl_640 | (fsm_output[0])));
  assign mux_918_nl = MUX_s_1_2_2(or_tmp_213, nand_728_cse_1, or_11_cse);
  assign FpAdd_8U_23U_is_addition_and_9_cse = core_wen & (~ and_dcpl_78) & (~ (mux_918_nl));
  assign mux_919_nl = MUX_s_1_2_2(nand_693_cse, nand_598_cse, or_11_cse);
  assign FpAdd_8U_23U_is_addition_and_10_cse = core_wen & (~ and_dcpl_78) & (~ (mux_919_nl));
  assign mux_920_nl = MUX_s_1_2_2(or_tmp_347, or_tmp_621, or_11_cse);
  assign FpAdd_8U_23U_is_addition_and_11_cse = core_wen & (~ and_dcpl_78) & (~ (mux_920_nl));
  assign mux_921_nl = MUX_s_1_2_2(nand_tmp_3, nand_602_cse_1, or_11_cse);
  assign IsZero_8U_23U_1_and_cse = core_wen & (~ and_dcpl_78) & (~ (mux_921_nl));
  assign mux_923_nl = MUX_s_1_2_2(nand_tmp_8, nand_598_cse, or_11_cse);
  assign IsZero_8U_23U_1_and_1_cse = core_wen & (~ and_dcpl_78) & (~ (mux_923_nl));
  assign nor_1336_cse_1 = ~((cfg_precision_1_sva_st_90!=2'b10));
  assign nor_1340_cse = ~((cfg_precision_1_sva_st_91!=2'b10));
  assign or_2010_cse = (cfg_precision_1_sva_st_90!=2'b10);
  assign or_5695_itm = IsNaN_8U_23U_land_lpi_1_dfm_4 | IsNaN_8U_23U_1_land_lpi_1_dfm_4;
  assign and_1693_nl = and_dcpl_1217 & or_11_cse;
  assign and_1695_nl = and_dcpl_1219 & or_11_cse;
  assign mux_1924_nl = MUX_s_1_2_2((~ (chn_inp_in_crt_sva_2_739_736_1[3])), or_2010_cse,
      or_11_cse);
  assign mux1h_34_itm = MUX1HOT_v_31_3_2((chn_inp_in_crt_sva_1_739_395_1[211:181]),
      (chn_inp_in_crt_sva_1_739_395_1[339:309]), ({12'b0 , (inp_lookup_else_else_o_acc_psp_sva[52:34])}),
      {(and_1693_nl) , (and_1695_nl) , (mux_1924_nl)});
  assign or_5694_itm = IsNaN_8U_23U_land_3_lpi_1_dfm_4 | IsNaN_8U_23U_1_land_3_lpi_1_dfm_4;
  assign mux1h_36_itm = MUX1HOT_v_31_3_2((chn_inp_in_crt_sva_1_739_395_1[179:149]),
      (chn_inp_in_crt_sva_1_739_395_1[307:277]), ({12'b0 , (inp_lookup_else_else_o_acc_psp_3_sva[52:34])}),
      {and_dcpl_1224 , and_dcpl_1226 , (~ mux_tmp_1845)});
  assign mux_1925_nl = MUX_s_1_2_2(and_dcpl_423, (chn_inp_in_crt_sva_1_739_395_1[341]),
      or_11_cse);
  assign mux1h_38_itm = MUX1HOT_v_31_3_2((chn_inp_in_crt_sva_1_739_395_1[115:85]),
      (chn_inp_in_crt_sva_1_739_395_1[243:213]), ({12'b0 , (inp_lookup_else_else_o_acc_psp_1_sva[52:34])}),
      {and_dcpl_1230 , and_dcpl_1232 , (~ (mux_1925_nl))});
  assign nor_1869_cse = ~(IsNaN_8U_23U_1_IsNaN_8U_23U_1_nand_itm_2 | IsNaN_8U_23U_1_nor_itm_2);
  assign or_6042_cse = IsNaN_8U_23U_land_1_lpi_1_dfm_st_3 | nor_1869_cse;
  assign and_4210_cse = (cfg_precision_1_sva_st_90==2'b10);
  assign or_5693_itm = IsNaN_8U_23U_land_2_lpi_1_dfm_4 | IsNaN_8U_23U_1_land_2_lpi_1_dfm_4;
  assign and_1711_nl = IsNaN_8U_23U_land_2_lpi_1_dfm_4 & (cfg_precision_1_sva_st_90==2'b10)
      & or_11_cse;
  assign and_1714_nl = (~ IsNaN_8U_23U_land_2_lpi_1_dfm_4) & (cfg_precision_1_sva_st_90==2'b10)
      & or_11_cse;
  assign mux_1926_nl = MUX_s_1_2_2((~ (chn_inp_in_crt_sva_2_739_736_1[1])), or_2010_cse,
      or_11_cse);
  assign mux1h_40_itm = MUX1HOT_v_31_3_2((chn_inp_in_crt_sva_1_739_395_1[147:117]),
      (chn_inp_in_crt_sva_1_739_395_1[275:245]), ({12'b0 , (inp_lookup_else_else_o_acc_psp_2_sva[52:34])}),
      {(and_1711_nl) , (and_1714_nl) , (mux_1926_nl)});
  assign nor_1310_nl = ~((cfg_precision_1_sva_st_90!=2'b10) | (chn_inp_in_crt_sva_1_739_395_1[341])
      | (~(main_stage_v_1 & (nor_5_cse | (or_5882_cse & FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_6_1_1
      & FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_6_0_1 & (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_9==4'b1111)
      & or_178_cse)))));
  assign and_3251_nl = (~((~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[0])
      | (cfg_precision_1_sva_st_91!=2'b10))) & (~(((~ IsNaN_6U_10U_7_land_1_lpi_1_dfm_5)
      | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_14) & (FpMul_6U_10U_2_lor_6_lpi_1_dfm_st_3
      | (~ inp_lookup_1_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs))));
  assign mux_940_nl = MUX_s_1_2_2((and_3251_nl), (nor_1310_nl), or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_24_cse = core_wen & (~ and_dcpl_78)
      & (mux_940_nl);
  assign nor_1318_cse = ~((~ main_stage_v_1) | (cfg_precision_1_sva_st_90!=2'b10));
  assign nor_1697_cse = ~((~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10));
  assign nor_1309_nl = ~((cfg_precision_1_sva_st_90!=2'b10) | (chn_inp_in_crt_sva_1_739_395_1[342])
      | (~(main_stage_v_1 & (nor_13_cse | (or_5889_cse & FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_6_1_1
      & FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_6_0_1 & (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_9==4'b1111)
      & (~((FpFractionToFloat_35U_6U_10U_1_mux_40_tmp==5'b11111) & (IntLeadZero_35U_1_leading_sign_35_0_rtn_2_sva_2[5])
      & inp_lookup_2_FpMantRNE_36U_11U_1_else_and_svs_2 & (~ IsNaN_6U_10U_6_nor_1_tmp)
      & FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_st_2)))))));
  assign and_3250_nl = (~((~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[1])
      | (cfg_precision_1_sva_st_91!=2'b10))) & (~(((~ IsNaN_6U_10U_7_land_2_lpi_1_dfm_5)
      | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_14) & (FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_3
      | (~ inp_lookup_2_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs))));
  assign mux_942_nl = MUX_s_1_2_2((and_3250_nl), (nor_1309_nl), or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_27_cse = core_wen & (~ and_dcpl_78)
      & (mux_942_nl);
  assign and_3249_cse = inp_lookup_3_IsNaN_6U_10U_7_aif_IsNaN_6U_10U_7_aelse_IsNaN_6U_10U_7_aelse_or_tmp
      & FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_6_1_1 & FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_6_0_1
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_3_lpi_1_dfm_9==4'b1111);
  assign nor_301_cse = ~(FpMul_6U_10U_2_if_2_FpMul_6U_10U_2_if_2_or_5_tmp | (~ inp_lookup_3_FpMul_6U_10U_2_else_2_if_acc_itm_6_1));
  assign nor_1304_nl = ~((cfg_precision_1_sva_st_90!=2'b10) | (chn_inp_in_crt_sva_1_739_395_1[344])
      | (~(main_stage_v_1 & (nor_29_cse | (or_5904_cse & FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_6_1_1
      & FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_6_0_1 & (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_9==4'b1111)
      & (~((FpFractionToFloat_35U_6U_10U_1_mux_42_tmp==5'b11111) & (IntLeadZero_35U_1_leading_sign_35_0_rtn_sva_2[5])
      & inp_lookup_4_FpMantRNE_36U_11U_1_else_and_svs_2 & (~ IsNaN_6U_10U_6_nor_3_tmp)
      & FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2)))))));
  assign and_3248_nl = nor_74_cse & (~(((~ IsNaN_6U_10U_7_land_lpi_1_dfm_5) | IsNaN_6U_10U_2_land_lpi_1_dfm_st_14)
      & (FpMul_6U_10U_2_lor_1_lpi_1_dfm_st_3 | (~ inp_lookup_4_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs))));
  assign mux_948_nl = MUX_s_1_2_2((and_3248_nl), (nor_1304_nl), or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_33_cse = core_wen & (~ and_dcpl_78)
      & (mux_948_nl);
  assign and_3246_cse = FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_7_1_1
      & FpAdd_8U_23U_o_sign_1_lpi_1_dfm_7 & inp_lookup_1_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_tmp
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_9==4'b1111);
  assign and_1717_rgt = ((~((inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_4_0_1[4])
      & (inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_4_0_1[0]))) | (~((inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_4_0_1[2:1]==2'b11)))
      | (~((inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_4_0_1[3]) & inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_5_1))
      | IsNaN_6U_10U_4_nor_tmp | (~ IsNaN_8U_23U_land_1_lpi_1_dfm_st_4)) & and_dcpl_459;
  assign and_1725_rgt = and_dcpl_459 & and_dcpl_1247 & (inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_4_0_1[3:1]==3'b111)
      & inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_5_1 & and_dcpl_1243;
  assign and_3244_cse = FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_7_1_1
      & FpAdd_8U_23U_o_sign_2_lpi_1_dfm_7 & inp_lookup_2_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_tmp
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_9==4'b1111);
  assign and_1726_rgt = ((inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_6_4_0_1[3:0]!=4'b1111)
      | (~(IsNaN_8U_23U_land_2_lpi_1_dfm_st_4 & (inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_6_4_0_1[4])))
      | (~ inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_6_5_1) | IsNaN_6U_10U_4_nor_1_tmp)
      & and_dcpl_488;
  assign and_1734_rgt = and_dcpl_488 & and_dcpl_1256 & (inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_6_4_0_1[3:2]==2'b11)
      & IsNaN_8U_23U_land_2_lpi_1_dfm_st_4 & (inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_6_4_0_1[4])
      & and_dcpl_1252;
  assign and_3242_cse = FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_7_1_1
      & FpAdd_8U_23U_o_sign_3_lpi_1_dfm_7 & inp_lookup_3_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_tmp
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_9==4'b1111);
  assign and_1735_rgt = ((inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_6_4_0_1[3:0]!=4'b1111)
      | (~(IsNaN_8U_23U_land_3_lpi_1_dfm_st_4 & (inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_6_4_0_1[4])))
      | (~ inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_6_5_1) | IsNaN_6U_10U_4_nor_2_tmp)
      & and_dcpl_524;
  assign and_1743_rgt = and_dcpl_524 & and_dcpl_1265 & (inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_6_4_0_1[3:2]==2'b11)
      & IsNaN_8U_23U_land_3_lpi_1_dfm_st_4 & (inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_6_4_0_1[4])
      & and_dcpl_1261;
  assign and_3240_cse = FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_7_1_1
      & FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_7_0_1 & inp_lookup_4_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_tmp
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_9==4'b1111);
  assign and_1744_rgt = ((inp_lookup_else_if_a0_15_10_lpi_1_dfm_6_4_0_1[3:0]!=4'b1111)
      | (~(IsNaN_8U_23U_land_lpi_1_dfm_st_4 & (inp_lookup_else_if_a0_15_10_lpi_1_dfm_6_4_0_1[4])))
      | (~ inp_lookup_else_if_a0_15_10_lpi_1_dfm_6_5_1) | IsNaN_6U_10U_4_nor_3_tmp)
      & and_dcpl_559;
  assign and_1752_rgt = and_dcpl_559 & and_dcpl_1274 & (inp_lookup_else_if_a0_15_10_lpi_1_dfm_6_4_0_1[3:2]==2'b11)
      & IsNaN_8U_23U_land_lpi_1_dfm_st_4 & (inp_lookup_else_if_a0_15_10_lpi_1_dfm_6_4_0_1[4])
      & and_dcpl_1270;
  assign and_1754_rgt = and_dcpl_459 & (~(FpMul_6U_10U_1_if_2_FpMul_6U_10U_1_if_2_or_tmp
      | inp_lookup_1_FpMul_6U_10U_1_oelse_1_acc_itm_7_1));
  assign and_1755_rgt = and_dcpl_459 & or_457_cse;
  assign and_1757_rgt = and_dcpl_488 & (~(FpMul_6U_10U_1_if_2_FpMul_6U_10U_1_if_2_or_2_tmp
      | inp_lookup_2_FpMul_6U_10U_1_oelse_1_acc_itm_7_1));
  assign and_1758_rgt = and_dcpl_488 & or_519_cse;
  assign and_1760_rgt = and_dcpl_524 & (~(FpMul_6U_10U_1_if_2_FpMul_6U_10U_1_if_2_or_4_tmp
      | inp_lookup_3_FpMul_6U_10U_1_oelse_1_acc_itm_7_1));
  assign and_1761_rgt = and_dcpl_524 & or_593_cse;
  assign nor_1274_cse = ~(FpMul_6U_10U_2_lor_6_lpi_1_dfm_6 | FpMul_6U_10U_2_FpMul_6U_10U_2_and_itm_2);
  assign or_2176_cse = (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10);
  assign nor_1273_cse = ~(nor_1274_cse | FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_2);
  assign IsNaN_6U_10U_7_aelse_and_4_cse = core_wen & (~ and_dcpl_78) & (~ mux_197_itm);
  assign or_2197_nl = IsNaN_6U_10U_7_land_1_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_14
      | (cfg_precision_1_sva_st_91!=2'b10);
  assign mux_973_nl = MUX_s_1_2_2((or_2197_nl), or_tmp_439, chn_inp_in_crt_sva_2_739_736_1[0]);
  assign and_3230_nl = main_stage_v_2 & (~ (mux_973_nl));
  assign or_2198_nl = (cfg_precision_1_sva_st_80!=2'b10) | IsNaN_6U_10U_7_land_1_lpi_1_dfm_6
      | IsNaN_6U_10U_6_land_1_lpi_1_dfm_5;
  assign mux_974_nl = MUX_s_1_2_2((or_2198_nl), or_tmp_440, chn_inp_in_crt_sva_3_739_736_1[0]);
  assign and_3231_nl = main_stage_v_3 & (~ (mux_974_nl));
  assign mux_975_nl = MUX_s_1_2_2((and_3231_nl), (and_3230_nl), or_11_cse);
  assign FpMul_6U_10U_2_oelse_1_and_8_cse = core_wen & FpMul_6U_10U_2_oelse_1_FpMul_6U_10U_2_oelse_1_or_11_cse
      & (mux_975_nl);
  assign nor_1790_cse = ~(FpMul_6U_10U_2_lor_7_lpi_1_dfm_6 | FpMul_6U_10U_2_FpMul_6U_10U_2_and_16_itm_2);
  assign nor_1264_cse = ~(nor_1790_cse | FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_2);
  assign or_2232_nl = (cfg_precision_1_sva_st_91!=2'b10) | IsNaN_6U_10U_7_land_2_lpi_1_dfm_5
      | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_14;
  assign mux_983_nl = MUX_s_1_2_2((or_2232_nl), or_tmp_439, chn_inp_in_crt_sva_2_739_736_1[1]);
  assign and_3228_nl = main_stage_v_2 & (~ (mux_983_nl));
  assign or_2233_nl = IsNaN_6U_10U_6_land_2_lpi_1_dfm_5 | IsNaN_6U_10U_7_land_2_lpi_1_dfm_6
      | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_984_nl = MUX_s_1_2_2((or_2233_nl), or_tmp_440, chn_inp_in_crt_sva_3_739_736_1[1]);
  assign and_3229_nl = main_stage_v_3 & (~ (mux_984_nl));
  assign mux_985_nl = MUX_s_1_2_2((and_3229_nl), (and_3228_nl), or_11_cse);
  assign FpMul_6U_10U_2_oelse_1_and_9_cse = core_wen & IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_2_cse
      & (mux_985_nl);
  assign nor_1789_cse = ~(FpMul_6U_10U_2_lor_8_lpi_1_dfm_6 | FpMul_6U_10U_2_FpMul_6U_10U_2_and_17_itm_2);
  assign nor_1251_cse = ~(nor_1789_cse | FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_2);
  assign or_2269_nl = (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10) | IsNaN_6U_10U_7_land_3_lpi_1_dfm_5
      | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_14;
  assign mux_993_nl = MUX_s_1_2_2((or_2269_nl), or_2176_cse, chn_inp_in_crt_sva_2_739_736_1[2]);
  assign or_2270_nl = IsNaN_6U_10U_7_land_3_lpi_1_dfm_6 | IsNaN_6U_10U_6_land_3_lpi_1_dfm_5
      | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_994_nl = MUX_s_1_2_2((or_2270_nl), or_tmp_440, chn_inp_in_crt_sva_3_739_736_1[2]);
  assign nand_116_nl = ~(main_stage_v_3 & (~ (mux_994_nl)));
  assign mux_995_nl = MUX_s_1_2_2((nand_116_nl), (mux_993_nl), or_11_cse);
  assign FpMul_6U_10U_2_oelse_1_and_10_cse = core_wen & IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_1_cse
      & (~ (mux_995_nl));
  assign nand_661_cse = ~((chn_inp_in_crt_sva_3_739_736_1[3]) & main_stage_v_3 &
      (cfg_precision_1_sva_st_80==2'b10));
  assign nor_1238_cse = ~(FpMul_6U_10U_2_lor_1_lpi_1_dfm_6 | FpMul_6U_10U_2_FpMul_6U_10U_2_and_18_itm_2);
  assign or_2282_cse = (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10);
  assign nor_1237_cse = ~(nor_1238_cse | FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_sva_2);
  assign or_2296_nl = (cfg_precision_1_sva_st_91!=2'b10) | IsNaN_6U_10U_7_land_lpi_1_dfm_5
      | IsNaN_6U_10U_2_land_lpi_1_dfm_st_14;
  assign mux_1004_nl = MUX_s_1_2_2((or_2296_nl), or_tmp_439, chn_inp_in_crt_sva_2_739_736_1[3]);
  assign and_3226_nl = main_stage_v_2 & (~ (mux_1004_nl));
  assign and_3227_nl = main_stage_v_3 & (~((~(FpMul_6U_10U_2_FpMul_6U_10U_2_nor_3_ssc
      | (chn_inp_in_crt_sva_3_739_736_1[3]))) | (cfg_precision_1_sva_st_80!=2'b10)));
  assign mux_1005_nl = MUX_s_1_2_2((and_3227_nl), (and_3226_nl), or_11_cse);
  assign FpMul_6U_10U_2_oelse_1_and_11_cse = core_wen & IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_cse
      & (mux_1005_nl);
  assign and_1764_rgt = or_11_cse & or_648_cse;
  assign mux_1927_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_4_739_736_1[0]), (chn_inp_in_crt_sva_3_739_736_1[0]),
      or_11_cse);
  assign FpAdd_8U_23U_o_expo_FpAdd_8U_23U_o_expo_mux_rgt = MUX_v_8_2_2(({2'b0 , FpMul_6U_10U_1_else_2_else_ac_int_cctor_1_sva_mx0w0}),
      FpAdd_8U_23U_o_expo_1_lpi_1_dfm_7_mx1w1, mux_1927_nl);
  assign nor_1221_cse = ~((~ main_stage_v_4) | (cfg_precision_1_sva_st_81!=2'b10));
  assign nor_1217_cse = ~((~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10));
  assign nor_1225_cse = ~(FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_1_st_2 | FpMul_6U_10U_1_lor_6_lpi_1_dfm_6);
  assign nor_1224_cse = ~(nor_1225_cse | FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_9_1);
  assign mux_1015_cse = MUX_s_1_2_2((~ inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4),
      inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4,
      inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4);
  assign and_1768_rgt = or_11_cse & (~ IsNaN_6U_10U_6_land_1_lpi_1_dfm_5);
  assign nor_1210_cse = ~(FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_3 | (~ inp_lookup_1_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs));
  assign mux_1928_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_4_739_736_1[1]), (chn_inp_in_crt_sva_3_739_736_1[1]),
      or_11_cse);
  assign FpAdd_8U_23U_o_expo_FpAdd_8U_23U_o_expo_mux_1_rgt = MUX_v_8_2_2(({2'b0 ,
      FpMul_6U_10U_1_else_2_else_ac_int_cctor_2_sva_mx0w0}), FpAdd_8U_23U_o_expo_2_lpi_1_dfm_7_mx1w1,
      mux_1928_nl);
  assign nor_1208_cse = ~(FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_1_st_2 | FpMul_6U_10U_1_lor_7_lpi_1_dfm_6);
  assign nor_1207_cse = ~(nor_1208_cse | FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_9_1);
  assign mux_1031_cse = MUX_s_1_2_2((~ inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4),
      inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4,
      inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4);
  assign and_1772_rgt = or_11_cse & (~ IsNaN_6U_10U_6_land_2_lpi_1_dfm_5);
  assign nor_1193_cse = ~(FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_3 | (~ inp_lookup_2_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs));
  assign mux_1929_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_4_739_736_1[2]), (chn_inp_in_crt_sva_3_739_736_1[2]),
      or_11_cse);
  assign FpAdd_8U_23U_o_expo_FpAdd_8U_23U_o_expo_mux_2_rgt = MUX_v_8_2_2(({2'b0 ,
      FpMul_6U_10U_1_else_2_else_ac_int_cctor_3_sva_mx0w0}), FpAdd_8U_23U_o_expo_3_lpi_1_dfm_7_mx1w1,
      mux_1929_nl);
  assign nor_1191_cse = ~(FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_1_st_2 | FpMul_6U_10U_1_lor_8_lpi_1_dfm_6);
  assign nor_1190_cse = ~(nor_1191_cse | FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_9_1);
  assign and_1776_rgt = or_11_cse & (~ IsNaN_6U_10U_6_land_3_lpi_1_dfm_5);
  assign mux_1930_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_4_739_736_1[3]), (chn_inp_in_crt_sva_3_739_736_1[3]),
      or_11_cse);
  assign FpAdd_8U_23U_o_expo_FpAdd_8U_23U_o_expo_mux_3_rgt = MUX_v_8_2_2(({2'b0 ,
      FpMul_6U_10U_1_else_2_else_ac_int_cctor_sva_mx0w0}), FpAdd_8U_23U_o_expo_lpi_1_dfm_7_mx1w1,
      mux_1930_nl);
  assign or_5689_cse = (~ (inp_lookup_4_FpMul_6U_10U_1_p_mant_p1_mul_tmp[21])) |
      inp_lookup_4_FpMul_6U_10U_1_else_2_else_if_if_acc_1_itm_5_1;
  assign nor_1180_cse = ~(FpMul_6U_10U_1_lor_1_lpi_1_dfm_6 | FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_1_st_2);
  assign nand_432_nl = ~(main_stage_v_3 & inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4
      & (chn_inp_in_crt_sva_3_739_736_1[3]) & (cfg_precision_1_sva_st_80==2'b10));
  assign mux_1058_nl = MUX_s_1_2_2(nand_tmp_126, (nand_432_nl), or_11_cse);
  assign or_2433_nl = (~ main_stage_v_3) | inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4
      | (~ (chn_inp_in_crt_sva_3_739_736_1[3])) | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_1059_nl = MUX_s_1_2_2(nand_tmp_126, (or_2433_nl), or_11_cse);
  assign mux_1060_nl = MUX_s_1_2_2((mux_1059_nl), (mux_1058_nl), FpMul_6U_10U_2_else_2_else_if_if_slc_FpMul_6U_10U_2_else_2_else_if_if_acc_1_5_mdf_sva_st_2);
  assign IsZero_8U_23U_3_and_3_cse = core_wen & (~ and_dcpl_78) & (~ (mux_1060_nl));
  assign mux_1061_cse = MUX_s_1_2_2(inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4,
      (~ inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4),
      FpMul_6U_10U_2_else_2_else_if_if_slc_FpMul_6U_10U_2_else_2_else_if_if_acc_1_5_mdf_sva_st_2);
  assign and_1780_rgt = or_11_cse & (~ IsNaN_6U_10U_6_land_lpi_1_dfm_5);
  assign or_2444_cse = (~ IsNaN_8U_23U_2_land_lpi_1_dfm_st_7) | (cfg_precision_1_sva_st_81!=2'b10);
  assign or_2445_cse = IsNaN_8U_23U_2_land_lpi_1_dfm_st_7 | (cfg_precision_1_sva_st_81!=2'b10);
  assign mux_1064_nl = MUX_s_1_2_2(or_2445_cse, or_2444_cse, or_tmp_2441);
  assign nor_1171_nl = ~((~ main_stage_v_4) | (~ (chn_inp_in_crt_sva_4_739_736_1[3]))
      | FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_4 | (mux_1064_nl));
  assign nor_1172_nl = ~((~ (chn_inp_in_crt_sva_5_739_736_1[3])) | IsNaN_8U_23U_2_land_lpi_1_dfm_9
      | (~ IsNaN_8U_23U_3_land_lpi_1_dfm_5) | (cfg_precision_1_sva_st_82[0]) | not_tmp_374);
  assign mux_1065_nl = MUX_s_1_2_2((nor_1172_nl), (nor_1171_nl), or_11_cse);
  assign FpAdd_8U_23U_o_expo_and_12_ssc = core_wen & (~ and_dcpl_78) & (mux_1065_nl);
  assign IsNaN_8U_23U_3_aelse_and_4_cse = core_wen & IsNaN_8U_23U_2_aelse_IsNaN_8U_23U_2_aelse_or_cse
      & (~ mux_1066_itm);
  assign IsNaN_8U_23U_3_aelse_and_5_cse = core_wen & FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_1_cse
      & (~ mux_1067_itm);
  assign nor_1169_nl = ~((~ main_stage_v_4) | IsNaN_6U_10U_5_land_2_lpi_1_dfm_6 |
      (~ (chn_inp_in_crt_sva_4_739_736_1[1])) | (~ FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_4)
      | (cfg_precision_1_sva_st_81!=2'b10));
  assign nor_1170_nl = ~((~ (chn_inp_in_crt_sva_5_739_736_1[1])) | (~ IsNaN_8U_23U_3_land_2_lpi_1_dfm_6)
      | IsNaN_8U_23U_2_land_2_lpi_1_dfm_9 | (cfg_precision_1_sva_st_82!=2'b10) |
      (~ main_stage_v_5));
  assign mux_1068_nl = MUX_s_1_2_2((nor_1170_nl), (nor_1169_nl), or_11_cse);
  assign FpAdd_8U_23U_o_expo_and_13_ssc = core_wen & (~ and_dcpl_78) & (mux_1068_nl);
  assign IsNaN_8U_23U_3_aelse_and_6_cse = core_wen & FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_2_cse
      & (~ mux_1067_itm);
  assign nor_1167_nl = ~((~ main_stage_v_4) | IsNaN_6U_10U_5_land_1_lpi_1_dfm_6 |
      (~ FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_4) | (~ (chn_inp_in_crt_sva_4_739_736_1[0]))
      | (cfg_precision_1_sva_st_81!=2'b10));
  assign nor_1168_nl = ~((~ (chn_inp_in_crt_sva_5_739_736_1[0])) | IsNaN_8U_23U_2_land_1_lpi_1_dfm_9
      | (~ IsNaN_8U_23U_3_land_1_lpi_1_dfm_6) | (cfg_precision_1_sva_st_82[0]) |
      not_tmp_374);
  assign mux_1070_nl = MUX_s_1_2_2((nor_1168_nl), (nor_1167_nl), or_11_cse);
  assign FpAdd_8U_23U_o_expo_and_14_ssc = core_wen & (~ and_dcpl_78) & (mux_1070_nl);
  assign IsNaN_8U_23U_3_aelse_and_7_cse = core_wen & FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_3_cse
      & (~ mux_1066_itm);
  assign mux_1931_nl = MUX_s_1_2_2(IsNaN_8U_23U_2_land_1_lpi_1_dfm_9, IsNaN_6U_10U_5_land_1_lpi_1_dfm_6,
      or_11_cse);
  assign mux1h_47_itm = MUX_v_31_2_2(({8'b0 , FpAdd_8U_23U_o_mant_1_lpi_1_dfm_6}),
      (chn_inp_in_crt_sva_4_127_0_1[30:0]), mux_1931_nl);
  assign mux_1932_nl = MUX_s_1_2_2(IsNaN_8U_23U_2_land_2_lpi_1_dfm_9, IsNaN_6U_10U_5_land_2_lpi_1_dfm_6,
      or_11_cse);
  assign mux1h_49_itm = MUX_v_31_2_2(({8'b0 , FpAdd_8U_23U_o_mant_2_lpi_1_dfm_6}),
      (chn_inp_in_crt_sva_4_127_0_1[62:32]), mux_1932_nl);
  assign mux_1933_nl = MUX_s_1_2_2(IsNaN_8U_23U_2_land_3_lpi_1_dfm_9, IsNaN_6U_10U_5_land_3_lpi_1_dfm_6,
      or_11_cse);
  assign mux1h_51_itm = MUX_v_31_2_2(({8'b0 , FpAdd_8U_23U_o_mant_3_lpi_1_dfm_6}),
      (chn_inp_in_crt_sva_4_127_0_1[94:64]), mux_1933_nl);
  assign mux_1934_nl = MUX_s_1_2_2(IsNaN_8U_23U_2_land_lpi_1_dfm_9, FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_4,
      or_11_cse);
  assign mux1h_53_itm = MUX_v_31_2_2(({8'b0 , FpAdd_8U_23U_o_mant_lpi_1_dfm_6}),
      (chn_inp_in_crt_sva_4_127_0_1[126:96]), mux_1934_nl);
  assign and_1794_rgt = (~(FpAdd_6U_10U_1_is_a_greater_acc_itm_6 | (chn_inp_in_crt_sva_4_739_736_1[0])))
      & or_11_cse;
  assign and_1796_rgt = FpAdd_6U_10U_1_is_a_greater_acc_itm_6 & (~ (chn_inp_in_crt_sva_4_739_736_1[0]))
      & or_11_cse;
  assign or_2486_nl = (~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[0]) |
      (cfg_precision_1_sva_st_81!=2'b10);
  assign mux_1081_nl = MUX_s_1_2_2(or_tmp_2486, (or_2486_nl), or_11_cse);
  assign FpAdd_6U_10U_1_is_addition_and_cse = core_wen & (~ and_dcpl_78) & (~ (mux_1081_nl));
  assign and_1798_rgt = (~(FpAdd_6U_10U_1_is_a_greater_acc_1_itm_6 | (chn_inp_in_crt_sva_4_739_736_1[1])))
      & or_11_cse;
  assign and_1800_rgt = FpAdd_6U_10U_1_is_a_greater_acc_1_itm_6 & (~ (chn_inp_in_crt_sva_4_739_736_1[1]))
      & or_11_cse;
  assign or_2490_nl = (~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[1]) |
      (cfg_precision_1_sva_st_81!=2'b10);
  assign mux_1082_nl = MUX_s_1_2_2(or_tmp_2490, (or_2490_nl), or_11_cse);
  assign FpAdd_6U_10U_1_is_addition_and_1_cse = core_wen & (~ and_dcpl_78) & (~ (mux_1082_nl));
  assign and_1802_rgt = (~(FpAdd_6U_10U_1_is_a_greater_acc_2_itm_6 | (chn_inp_in_crt_sva_4_739_736_1[2])))
      & or_11_cse;
  assign and_1804_rgt = FpAdd_6U_10U_1_is_a_greater_acc_2_itm_6 & (~ (chn_inp_in_crt_sva_4_739_736_1[2]))
      & or_11_cse;
  assign or_2494_nl = (~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[2]) |
      (cfg_precision_1_sva_st_81!=2'b10);
  assign mux_1083_nl = MUX_s_1_2_2(or_tmp_2494, (or_2494_nl), or_11_cse);
  assign FpAdd_6U_10U_1_is_addition_and_2_cse = core_wen & (~ and_dcpl_78) & (~ (mux_1083_nl));
  assign and_1806_rgt = (~(FpAdd_6U_10U_1_is_a_greater_acc_3_itm_6_1 | (chn_inp_in_crt_sva_4_739_736_1[3])))
      & or_11_cse;
  assign and_1808_rgt = FpAdd_6U_10U_1_is_a_greater_acc_3_itm_6_1 & (~ (chn_inp_in_crt_sva_4_739_736_1[3]))
      & or_11_cse;
  assign or_2498_nl = (~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[3]) |
      (cfg_precision_1_sva_st_81!=2'b10);
  assign mux_1084_nl = MUX_s_1_2_2(or_tmp_2498, (or_2498_nl), or_11_cse);
  assign FpAdd_6U_10U_1_is_addition_and_3_cse = core_wen & (~ and_dcpl_78) & (~ (mux_1084_nl));
  assign mux_1092_nl = MUX_s_1_2_2(chn_inp_in_crt_sva_4_411_1, (~ chn_inp_in_crt_sva_4_411_1),
      inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5);
  assign or_2525_nl = (~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[0]) |
      (cfg_precision_1_sva_st_81[0]) | (~((cfg_precision_1_sva_st_81[1]) & (~((~((~
      IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_tmp) & (~ IsNaN_6U_10U_9_nor_tmp) & FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_5_1
      & FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_4_1 & (FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_3_0_1==4'b1111)))
      & FpAdd_6U_10U_1_is_a_greater_acc_itm_6 & (mux_1092_nl)))));
  assign or_2531_nl = (~ IsNaN_8U_23U_2_land_1_lpi_1_dfm_st_7) | chn_inp_in_crt_sva_5_411_1;
  assign mux_1094_nl = MUX_s_1_2_2(or_tmp_2531, mux_tmp_1015, or_2531_nl);
  assign mux_1095_nl = MUX_s_1_2_2(or_tmp_2531, (mux_1094_nl), IsNaN_8U_23U_2_land_1_lpi_1_dfm_9);
  assign mux_1096_nl = MUX_s_1_2_2((mux_1095_nl), mux_tmp_1015, IsNaN_8U_23U_3_land_1_lpi_1_dfm_6);
  assign or_860_nl = (~ IsNaN_6U_10U_9_land_1_lpi_1_dfm_6) | IsNaN_6U_10U_8_land_1_lpi_1_dfm_6;
  assign mux_1097_nl = MUX_s_1_2_2(or_tmp_2531, (mux_1096_nl), or_860_nl);
  assign mux_1098_nl = MUX_s_1_2_2((mux_1097_nl), (or_2525_nl), or_11_cse);
  assign FpMul_6U_10U_2_o_expo_and_12_cse = core_wen & (~ and_dcpl_78) & (~ (mux_1098_nl));
  assign mux_1101_nl = MUX_s_1_2_2(mux_tmp_444, nand_tmp_138, or_11_cse);
  assign IsZero_6U_10U_9_and_cse = core_wen & FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_3_cse
      & (~ (mux_1101_nl));
  assign mux_1109_nl = MUX_s_1_2_2(chn_inp_in_crt_sva_4_427_1, (~ chn_inp_in_crt_sva_4_427_1),
      inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5);
  assign or_2562_nl = (~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[1]) |
      (cfg_precision_1_sva_st_81[0]) | (~((cfg_precision_1_sva_st_81[1]) & (~((~((~
      IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_1_tmp) & (~ IsNaN_6U_10U_9_nor_1_tmp) & FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_5_1
      & FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_4_1 & (FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_3_0_1==4'b1111)))
      & FpAdd_6U_10U_1_is_a_greater_acc_1_itm_6 & (mux_1109_nl)))));
  assign or_2568_nl = (~ IsNaN_8U_23U_2_land_2_lpi_1_dfm_st_7) | chn_inp_in_crt_sva_5_427_1;
  assign mux_1111_nl = MUX_s_1_2_2(or_tmp_2490, mux_tmp_1032, or_2568_nl);
  assign mux_1112_nl = MUX_s_1_2_2(or_tmp_2490, (mux_1111_nl), IsNaN_8U_23U_2_land_2_lpi_1_dfm_9);
  assign mux_1113_nl = MUX_s_1_2_2((mux_1112_nl), mux_tmp_1032, IsNaN_8U_23U_3_land_2_lpi_1_dfm_6);
  assign or_889_nl = (~ IsNaN_6U_10U_9_land_2_lpi_1_dfm_6) | IsNaN_6U_10U_8_land_2_lpi_1_dfm_4;
  assign mux_1114_nl = MUX_s_1_2_2(or_tmp_2490, (mux_1113_nl), or_889_nl);
  assign mux_1115_nl = MUX_s_1_2_2((mux_1114_nl), (or_2562_nl), or_11_cse);
  assign FpMul_6U_10U_2_o_expo_and_15_cse = core_wen & (~ and_dcpl_78) & (~ (mux_1115_nl));
  assign mux_1118_nl = MUX_s_1_2_2(mux_tmp_457, nand_tmp_142, or_11_cse);
  assign IsZero_6U_10U_9_and_1_cse = core_wen & FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_2_cse
      & (~ (mux_1118_nl));
  assign mux_1126_nl = MUX_s_1_2_2(chn_inp_in_crt_sva_4_443_1, (~ chn_inp_in_crt_sva_4_443_1),
      inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5);
  assign or_2599_nl = (~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[2]) |
      (cfg_precision_1_sva_st_81[0]) | (~((cfg_precision_1_sva_st_81[1]) & (~((~((~
      IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_2_tmp) & (~ IsNaN_6U_10U_9_nor_2_tmp) & FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_5_1
      & FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_4_1 & (FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_3_0_1==4'b1111)))
      & FpAdd_6U_10U_1_is_a_greater_acc_2_itm_6 & (mux_1126_nl)))));
  assign or_2605_nl = (~ IsNaN_8U_23U_2_land_3_lpi_1_dfm_st_7) | chn_inp_in_crt_sva_5_443_1;
  assign mux_1128_nl = MUX_s_1_2_2(or_tmp_2494, mux_tmp_1049, or_2605_nl);
  assign mux_1129_nl = MUX_s_1_2_2(or_tmp_2494, (mux_1128_nl), IsNaN_8U_23U_2_land_3_lpi_1_dfm_9);
  assign mux_1130_nl = MUX_s_1_2_2((mux_1129_nl), mux_tmp_1049, IsNaN_8U_23U_3_land_3_lpi_1_dfm_6);
  assign or_926_nl = (~ IsNaN_6U_10U_9_land_3_lpi_1_dfm_6) | IsNaN_6U_10U_8_land_3_lpi_1_dfm_4;
  assign mux_1131_nl = MUX_s_1_2_2(or_tmp_2494, (mux_1130_nl), or_926_nl);
  assign mux_1132_nl = MUX_s_1_2_2((mux_1131_nl), (or_2599_nl), or_11_cse);
  assign FpMul_6U_10U_2_o_expo_and_18_cse = core_wen & (~ and_dcpl_78) & (~ (mux_1132_nl));
  assign mux_1135_nl = MUX_s_1_2_2(mux_tmp_467, nand_tmp_146, or_11_cse);
  assign IsZero_6U_10U_9_and_2_cse = core_wen & FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_1_cse
      & (~ (mux_1135_nl));
  assign mux_1140_cse = MUX_s_1_2_2((~ chn_inp_in_crt_sva_4_459_1), chn_inp_in_crt_sva_4_459_1,
      IsNaN_8U_23U_2_land_lpi_1_dfm_st_7);
  assign nor_1130_cse = ~((~ IsNaN_8U_23U_2_land_lpi_1_dfm_st_8) | chn_inp_in_crt_sva_5_459_1);
  assign mux_1144_nl = MUX_s_1_2_2(chn_inp_in_crt_sva_4_459_1, (~ chn_inp_in_crt_sva_4_459_1),
      IsNaN_8U_23U_2_land_lpi_1_dfm_st_7);
  assign or_2637_nl = (~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[3]) |
      (cfg_precision_1_sva_st_81[0]) | (~((cfg_precision_1_sva_st_81[1]) & (~((~((~
      IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_3_tmp) & (~ IsNaN_6U_10U_9_nor_3_tmp) & FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_5_1
      & FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_4_1 & (FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_3_0_1==4'b1111)))
      & FpAdd_6U_10U_1_is_a_greater_acc_3_itm_6_1 & (mux_1144_nl)))));
  assign or_2643_nl = (~ IsNaN_8U_23U_2_land_lpi_1_dfm_st_8) | chn_inp_in_crt_sva_5_459_1;
  assign mux_1146_nl = MUX_s_1_2_2(or_tmp_2643, mux_tmp_1067, or_2643_nl);
  assign mux_1147_nl = MUX_s_1_2_2(or_tmp_2643, (mux_1146_nl), IsNaN_8U_23U_2_land_lpi_1_dfm_9);
  assign mux_1148_nl = MUX_s_1_2_2((mux_1147_nl), mux_tmp_1067, IsNaN_8U_23U_3_land_lpi_1_dfm_5);
  assign or_2638_nl = (~ IsNaN_6U_10U_9_land_lpi_1_dfm_6) | IsNaN_6U_10U_8_land_lpi_1_dfm_4;
  assign mux_1149_nl = MUX_s_1_2_2(or_tmp_2643, (mux_1148_nl), or_2638_nl);
  assign mux_1150_nl = MUX_s_1_2_2((mux_1149_nl), (or_2637_nl), or_11_cse);
  assign FpMul_6U_10U_2_o_expo_and_21_cse = core_wen & (~ and_dcpl_78) & (~ (mux_1150_nl));
  assign mux_1153_nl = MUX_s_1_2_2(mux_tmp_478, nand_tmp_148, or_11_cse);
  assign IsZero_6U_10U_9_and_3_cse = core_wen & IsNaN_8U_23U_2_aelse_IsNaN_8U_23U_2_aelse_or_cse
      & (~ (mux_1153_nl));
  assign nor_1124_cse = ~((chn_inp_in_crt_sva_5_739_736_1[0]) | (cfg_precision_1_sva_st_82[0])
      | not_tmp_374);
  assign and_1816_rgt = (~(IsNaN_8U_23U_3_land_1_lpi_1_dfm_6 | IsNaN_8U_23U_2_land_1_lpi_1_dfm_9))
      & (chn_inp_in_crt_sva_5_739_736_1[0]) & or_11_cse;
  assign and_1821_rgt = or_dcpl_727 & and_dcpl_688;
  assign or_2663_cse = (~ inp_lookup_2_FpMantRNE_49U_24U_1_else_and_tmp) | inp_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_1_itm_7_1;
  assign and_1829_rgt = (~(IsNaN_8U_23U_3_land_2_lpi_1_dfm_6 | IsNaN_8U_23U_2_land_2_lpi_1_dfm_9))
      & (chn_inp_in_crt_sva_5_739_736_1[1]) & or_11_cse;
  assign and_1834_rgt = or_dcpl_732 & and_dcpl_699;
  assign and_1842_rgt = (~(IsNaN_8U_23U_3_land_3_lpi_1_dfm_6 | IsNaN_8U_23U_2_land_3_lpi_1_dfm_9))
      & (chn_inp_in_crt_sva_5_739_736_1[2]) & or_11_cse;
  assign or_2676_cse = (~ inp_lookup_3_FpMantRNE_49U_24U_1_else_and_tmp) | inp_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_1_itm_7;
  assign and_1847_rgt = or_dcpl_737 & or_11_cse & (~ IsNaN_8U_23U_3_land_3_lpi_1_dfm_6);
  assign nor_1113_cse = ~((chn_inp_in_crt_sva_5_739_736_1[3]) | (cfg_precision_1_sva_st_82[0])
      | not_tmp_374);
  assign and_1855_rgt = (~(IsNaN_8U_23U_3_land_lpi_1_dfm_5 | IsNaN_8U_23U_2_land_lpi_1_dfm_9))
      & (chn_inp_in_crt_sva_5_739_736_1[3]) & or_11_cse;
  assign and_1860_rgt = or_dcpl_742 & and_dcpl_717;
  assign and_3875_ssc = core_wen & (cfg_precision_1_sva_st_83==2'b10) & or_tmp_2703
      & main_stage_v_6 & (~ (chn_inp_in_crt_sva_6_739_736_1[2])) & or_11_cse;
  assign nor_1913_cse = ~((chn_inp_in_crt_sva_6_739_736_1[2]) | IsNaN_6U_10U_9_land_3_lpi_1_dfm_7
      | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_18);
  assign mux_2117_nl = MUX_s_1_2_2(or_tmp_4737, nor_1913_cse, inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8);
  assign or_6073_nl = inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8
      | inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7;
  assign mux_2118_nl = MUX_s_1_2_2((mux_2117_nl), or_tmp_4737, or_6073_nl);
  assign and_3880_cse = (~ (mux_2118_nl)) & core_wen & (cfg_precision_1_sva_st_83==2'b10)
      & or_11_cse & main_stage_v_6;
  assign mux_1941_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_7_739_736_1[0]), (chn_inp_in_crt_sva_6_739_736_1[0]),
      or_11_cse);
  assign FpMul_6U_10U_1_o_expo_mux1h_23_itm = MUX_v_4_2_2(FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_7_3_0_1,
      ({1'b0 , FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_2_sva_mx0w0}),
      mux_1941_nl);
  assign or_5680_cse = IsNaN_6U_10U_9_land_2_lpi_1_dfm_8 | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_19;
  assign mux_1942_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_7_739_736_1[1]), (chn_inp_in_crt_sva_6_739_736_1[1]),
      or_11_cse);
  assign FpMul_6U_10U_1_o_expo_mux1h_29_itm = MUX_v_4_2_2(FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_7_3_0_1,
      ({1'b0 , FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_3_sva_mx0w0}),
      mux_1942_nl);
  assign FpMul_6U_10U_1_o_expo_mux1h_35_itm = MUX_v_4_2_2(FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_7_3_0_1,
      ({1'b0 , FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_4_sva_mx0w0}),
      mux_tmp_1862);
  assign mux_1943_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_7_739_736_1[3]), (chn_inp_in_crt_sva_6_739_736_1[3]),
      or_11_cse);
  assign FpMul_6U_10U_1_o_expo_mux1h_41_itm = MUX_v_4_2_2(FpMul_6U_10U_1_o_expo_lpi_1_dfm_7_3_0_1,
      ({1'b0 , FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_1_sva_mx0w0}),
      mux_1943_nl);
  assign IsNaN_6U_10U_2_aelse_and_12_cse = core_wen & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_or_15_cse
      & (~ mux_623_itm);
  assign IsNaN_6U_10U_2_aelse_and_13_cse = core_wen & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_or_14_cse
      & (~ mux_632_itm);
  assign IsNaN_6U_10U_2_aelse_and_14_cse = core_wen & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_or_13_cse
      & (~ mux_623_itm);
  assign IsNaN_6U_10U_2_aelse_and_15_cse = core_wen & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_or_12_cse
      & (~ mux_623_itm);
  assign nor_1727_cse = ~(IsNaN_6U_10U_8_land_1_lpi_1_dfm_7 | IsNaN_6U_10U_9_land_1_lpi_1_dfm_8);
  assign and_1871_rgt = or_11_cse & FpAdd_6U_10U_1_or_12_cse;
  assign or_2797_cse = (~ IsNaN_6U_10U_1_land_1_lpi_1_dfm_5) | IsNaN_6U_10U_land_1_lpi_1_dfm_5;
  assign and_1873_rgt = or_11_cse & (~ IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_5);
  assign and_3374_cse = main_stage_v_8 & (chn_inp_in_crt_sva_8_739_736_1[1]) & (cfg_precision_1_sva_st_85==2'b10);
  assign or_2810_cse = (~ IsNaN_6U_10U_1_land_2_lpi_1_dfm_5) | IsNaN_6U_10U_land_2_lpi_1_dfm_5;
  assign and_1875_rgt = or_11_cse & (~ IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_5);
  assign and_1877_rgt = or_11_cse & (~ IsNaN_6U_10U_8_land_lpi_1_dfm_st_5);
  assign or_2822_cse = (~ IsNaN_6U_10U_1_land_lpi_1_dfm_5) | IsNaN_6U_10U_land_lpi_1_dfm_5;
  assign nor_1076_nl = ~((~ (chn_inp_in_crt_sva_8_739_736_1[0])) | (cfg_precision_1_sva_st_85!=2'b10)
      | (~ IsNaN_6U_10U_1_land_1_lpi_1_dfm_5) | IsNaN_6U_10U_land_1_lpi_1_dfm_5 |
      (~ main_stage_v_8));
  assign nor_1077_nl = ~((~ (chn_inp_in_crt_sva_9_739_736_1[0])) | IsNaN_6U_10U_land_1_lpi_1_dfm_6
      | (~ IsNaN_6U_10U_1_land_1_lpi_1_dfm_6) | (~ main_stage_v_9) | (cfg_precision_1_sva_st_86!=2'b10));
  assign mux_1221_nl = MUX_s_1_2_2((nor_1077_nl), (nor_1076_nl), or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_28_cse = core_wen & (~ and_dcpl_78)
      & (mux_1221_nl);
  assign or_5020_cse = inp_lookup_1_FpMul_6U_10U_oelse_1_acc_itm_7_1 | reg_FpMul_6U_10U_lor_3_lpi_1_dfm_3_cse;
  assign and_1881_rgt = (~ IsNaN_6U_10U_land_1_lpi_1_dfm_5) & IsNaN_6U_10U_1_land_1_lpi_1_dfm_5
      & or_11_cse;
  assign nor_1765_rgt = ~(inp_lookup_1_FpMul_6U_10U_oelse_1_acc_itm_7_1 | IsNaN_6U_10U_land_1_lpi_1_dfm_5
      | IsNaN_6U_10U_1_land_1_lpi_1_dfm_5 | reg_FpMul_6U_10U_lor_3_lpi_1_dfm_3_cse
      | (~ or_11_cse));
  assign and_1888_rgt = or_5020_cse & (~ IsNaN_6U_10U_land_1_lpi_1_dfm_5) & (~ IsNaN_6U_10U_1_land_1_lpi_1_dfm_5)
      & or_11_cse;
  assign nor_1070_nl = ~((cfg_precision_1_sva_st_85!=2'b10) | (~ (chn_inp_in_crt_sva_8_739_736_1[1]))
      | (~ IsNaN_6U_10U_1_land_2_lpi_1_dfm_5) | IsNaN_6U_10U_land_2_lpi_1_dfm_5 |
      (~ main_stage_v_8));
  assign nor_1071_nl = ~((~ (chn_inp_in_crt_sva_9_739_736_1[1])) | IsNaN_6U_10U_land_2_lpi_1_dfm_6
      | (~ IsNaN_6U_10U_1_land_2_lpi_1_dfm_6) | (~ main_stage_v_9) | (cfg_precision_1_sva_st_100!=2'b10));
  assign mux_1225_nl = MUX_s_1_2_2((nor_1071_nl), (nor_1070_nl), or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_31_cse = core_wen & (~ and_dcpl_78)
      & (mux_1225_nl);
  assign or_5021_cse = inp_lookup_2_FpMul_6U_10U_oelse_1_acc_itm_7_1 | reg_FpMul_6U_10U_lor_4_lpi_1_dfm_3_cse;
  assign and_1892_rgt = (~ IsNaN_6U_10U_land_2_lpi_1_dfm_5) & IsNaN_6U_10U_1_land_2_lpi_1_dfm_5
      & or_11_cse;
  assign nor_1764_rgt = ~(inp_lookup_2_FpMul_6U_10U_oelse_1_acc_itm_7_1 | IsNaN_6U_10U_land_2_lpi_1_dfm_5
      | IsNaN_6U_10U_1_land_2_lpi_1_dfm_5 | reg_FpMul_6U_10U_lor_4_lpi_1_dfm_3_cse
      | (~ or_11_cse));
  assign and_1899_rgt = or_5021_cse & (~ IsNaN_6U_10U_land_2_lpi_1_dfm_5) & (~ IsNaN_6U_10U_1_land_2_lpi_1_dfm_5)
      & or_11_cse;
  assign nor_1065_nl = ~((~ (chn_inp_in_crt_sva_8_739_736_1[2])) | (~ IsNaN_6U_10U_1_land_3_lpi_1_dfm_5)
      | IsNaN_6U_10U_land_3_lpi_1_dfm_5 | (cfg_precision_1_sva_st_85!=2'b10) | (~
      main_stage_v_8));
  assign nor_1066_nl = ~((~ (chn_inp_in_crt_sva_9_739_736_1[2])) | IsNaN_6U_10U_land_3_lpi_1_dfm_6
      | (~ IsNaN_6U_10U_1_land_3_lpi_1_dfm_6) | (~ main_stage_v_9) | (cfg_precision_1_sva_st_112!=2'b10));
  assign mux_1229_nl = MUX_s_1_2_2((nor_1066_nl), (nor_1065_nl), or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_34_cse = core_wen & (~ and_dcpl_78)
      & (mux_1229_nl);
  assign or_5022_cse = inp_lookup_3_FpMul_6U_10U_oelse_1_acc_itm_7_1 | reg_FpMul_6U_10U_lor_5_lpi_1_dfm_3_cse;
  assign and_1903_rgt = (~ IsNaN_6U_10U_land_3_lpi_1_dfm_5) & IsNaN_6U_10U_1_land_3_lpi_1_dfm_5
      & or_11_cse;
  assign nor_1763_rgt = ~(inp_lookup_3_FpMul_6U_10U_oelse_1_acc_itm_7_1 | IsNaN_6U_10U_land_3_lpi_1_dfm_5
      | IsNaN_6U_10U_1_land_3_lpi_1_dfm_5 | reg_FpMul_6U_10U_lor_5_lpi_1_dfm_3_cse
      | (~ or_11_cse));
  assign and_1910_rgt = or_5022_cse & (~ IsNaN_6U_10U_land_3_lpi_1_dfm_5) & (~ IsNaN_6U_10U_1_land_3_lpi_1_dfm_5)
      & or_11_cse;
  assign nor_1061_nl = ~((~ (chn_inp_in_crt_sva_8_739_736_1[3])) | (~ IsNaN_6U_10U_1_land_lpi_1_dfm_5)
      | IsNaN_6U_10U_land_lpi_1_dfm_5 | (cfg_precision_1_sva_st_85!=2'b10) | (~ main_stage_v_8));
  assign nor_1062_nl = ~((~ (chn_inp_in_crt_sva_9_739_736_1[3])) | IsNaN_6U_10U_land_lpi_1_dfm_6
      | (~ IsNaN_6U_10U_1_land_lpi_1_dfm_6) | (~ main_stage_v_9) | (cfg_precision_1_sva_st_124!=2'b10));
  assign mux_1233_nl = MUX_s_1_2_2((nor_1062_nl), (nor_1061_nl), or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_37_cse = core_wen & (~ and_dcpl_78)
      & (mux_1233_nl);
  assign or_5023_cse = inp_lookup_4_FpMul_6U_10U_oelse_1_acc_itm_7_1 | reg_FpMul_6U_10U_lor_lpi_1_dfm_3_cse;
  assign and_1914_rgt = (~ IsNaN_6U_10U_land_lpi_1_dfm_5) & IsNaN_6U_10U_1_land_lpi_1_dfm_5
      & or_11_cse;
  assign nor_1762_rgt = ~(inp_lookup_4_FpMul_6U_10U_oelse_1_acc_itm_7_1 | IsNaN_6U_10U_land_lpi_1_dfm_5
      | IsNaN_6U_10U_1_land_lpi_1_dfm_5 | reg_FpMul_6U_10U_lor_lpi_1_dfm_3_cse |
      (~ or_11_cse));
  assign and_1921_rgt = or_5023_cse & (~ IsNaN_6U_10U_land_lpi_1_dfm_5) & (~ IsNaN_6U_10U_1_land_lpi_1_dfm_5)
      & or_11_cse;
  assign mux_1237_nl = MUX_s_1_2_2(or_tmp_1502, nand_tmp_162, or_11_cse);
  assign IsZero_6U_10U_3_and_cse = core_wen & (~ and_dcpl_78) & (~ (mux_1237_nl));
  assign mux_1239_nl = MUX_s_1_2_2(or_tmp_1537, nand_tmp_163, or_11_cse);
  assign IsZero_6U_10U_3_and_1_cse = core_wen & (~ and_dcpl_78) & (~ (mux_1239_nl));
  assign mux_1241_nl = MUX_s_1_2_2(nand_774_cse, nand_tmp_164, or_11_cse);
  assign IsZero_6U_10U_3_and_2_cse = core_wen & (~ and_dcpl_78) & (~ (mux_1241_nl));
  assign mux_1243_nl = MUX_s_1_2_2(nand_773_cse, nand_tmp_165, or_11_cse);
  assign IsZero_6U_10U_3_and_3_cse = core_wen & (~ and_dcpl_78) & (~ (mux_1243_nl));
  assign or_2923_nl = nor_1896_cse | (chn_inp_in_crt_sva_10_739_736_1[3]) | inp_lookup_else_unequal_tmp_36
      | (~ main_stage_v_10);
  assign mux_1244_nl = MUX_s_1_2_2(or_tmp_1826, or_tmp_2924, or_11_cse);
  assign mux_1245_nl = MUX_s_1_2_2((mux_1244_nl), (or_2923_nl), inp_lookup_else_unequal_tmp_37);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_4_cse = core_wen & (~ and_dcpl_78)
      & (~ (mux_1245_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_9_cse
      = (or_11_cse & IsNaN_6U_10U_2_land_lpi_1_dfm_24) | and_dcpl_1448;
  assign or_2934_nl = (~ (chn_inp_in_crt_sva_10_739_736_1[3])) | (cfg_precision_1_sva_st_125!=2'b10)
      | (~((IsNaN_6U_10U_3_land_lpi_1_dfm_6 | IsNaN_6U_10U_2_land_lpi_1_dfm_24) &
      main_stage_v_10));
  assign mux_1247_nl = MUX_s_1_2_2(or_tmp_1806, (or_2934_nl), or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_39_cse = core_wen & FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_9_cse
      & (~ (mux_1247_nl));
  assign mux_1248_nl = MUX_s_1_2_2(or_tmp_1845, or_tmp_2935, or_11_cse);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_5_cse = core_wen & (~ and_dcpl_78)
      & (~ (mux_1248_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_8_cse
      = (or_11_cse & IsNaN_6U_10U_2_land_3_lpi_1_dfm_24) | and_dcpl_1450;
  assign or_2949_nl = (~ (chn_inp_in_crt_sva_10_739_736_1[2])) | (cfg_precision_1_sva_st_113!=2'b10)
      | not_tmp_1202;
  assign mux_1250_nl = MUX_s_1_2_2(or_1645_cse, (or_2949_nl), or_11_cse);
  assign or_2952_nl = nor_1896_cse | (~ (chn_inp_in_crt_sva_10_739_736_1[2])) | (cfg_precision_1_sva_st_113!=2'b10)
      | not_tmp_1202;
  assign mux_1251_nl = MUX_s_1_2_2((or_2952_nl), (mux_1250_nl), or_tmp_1770);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_41_cse = core_wen & FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_8_cse
      & (~ (mux_1251_nl));
  assign mux_1252_nl = MUX_s_1_2_2(or_tmp_1856, or_tmp_2953, or_11_cse);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_6_cse = core_wen & (~ and_dcpl_78)
      & (~ (mux_1252_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_7_cse
      = (or_11_cse & IsNaN_6U_10U_2_land_2_lpi_1_dfm_24) | and_dcpl_1452;
  assign or_2967_nl = (~ (chn_inp_in_crt_sva_10_739_736_1[1])) | (cfg_precision_1_sva_st_101[0])
      | not_tmp_1208;
  assign mux_1254_nl = MUX_s_1_2_2(or_1632_cse, (or_2967_nl), or_11_cse);
  assign or_2970_nl = nor_1896_cse | (~ (chn_inp_in_crt_sva_10_739_736_1[1])) | (cfg_precision_1_sva_st_101[0])
      | not_tmp_1208;
  assign mux_1255_nl = MUX_s_1_2_2((or_2970_nl), (mux_1254_nl), or_tmp_1724);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_43_cse = core_wen & FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_7_cse
      & (~ (mux_1255_nl));
  assign or_2973_nl = nor_1896_cse | (chn_inp_in_crt_sva_10_739_736_1[0]) | inp_lookup_else_unequal_tmp_36
      | (~ main_stage_v_10);
  assign mux_1256_nl = MUX_s_1_2_2(or_tmp_1818, or_tmp_2974, or_11_cse);
  assign mux_1257_nl = MUX_s_1_2_2((mux_1256_nl), (or_2973_nl), inp_lookup_else_unequal_tmp_37);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_7_cse = core_wen & (~ and_dcpl_78)
      & (~ (mux_1257_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_6_cse
      = (or_11_cse & IsNaN_6U_10U_2_land_1_lpi_1_dfm_24) | and_dcpl_1454;
  assign or_2983_nl = (~ (chn_inp_in_crt_sva_10_739_736_1[0])) | (cfg_precision_1_sva_st_87[0])
      | not_tmp_1212;
  assign mux_1260_nl = MUX_s_1_2_2(or_tmp_1687, (or_2983_nl), or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_45_cse = core_wen & FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_6_cse
      & (~ (mux_1260_nl));
  assign inp_lookup_if_or_6_rgt = ((~ FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_1_mx0w0)
      & inp_lookup_if_and_m1c_11) | (IsNaN_6U_10U_3_land_lpi_1_dfm_6 & inp_lookup_if_and_m1c_10);
  assign inp_lookup_if_or_7_rgt = (FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_1_mx0w0
      & inp_lookup_if_and_m1c_11) | (IsNaN_6U_10U_2_land_lpi_1_dfm_24 & inp_lookup_if_and_m1c_9);
  assign inp_lookup_if_and_31_rgt = inp_lookup_if_unequal_tmp_1_mx0w0 & and_dcpl_1722;
  assign and_1941_rgt = or_11_cse & (~ (chn_inp_in_crt_sva_10_739_736_1[3]));
  assign inp_lookup_if_or_4_rgt = ((~ FpAdd_6U_10U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0)
      & inp_lookup_if_and_m1c_8) | (IsNaN_6U_10U_3_land_3_lpi_1_dfm_6 & inp_lookup_if_and_m1c_7);
  assign inp_lookup_if_or_5_rgt = (FpAdd_6U_10U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0
      & inp_lookup_if_and_m1c_8) | (IsNaN_6U_10U_2_land_3_lpi_1_dfm_24 & inp_lookup_if_and_m1c_6);
  assign inp_lookup_if_and_23_rgt = inp_lookup_if_unequal_tmp_1_mx0w0 & and_1942_m1c;
  assign and_1943_rgt = or_11_cse & (~ (chn_inp_in_crt_sva_10_739_736_1[2]));
  assign inp_lookup_if_or_2_rgt = ((~ FpAdd_6U_10U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0)
      & inp_lookup_if_and_m1c_5) | (IsNaN_6U_10U_3_land_2_lpi_1_dfm_6 & inp_lookup_if_and_m1c_4);
  assign inp_lookup_if_or_3_rgt = (FpAdd_6U_10U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0
      & inp_lookup_if_and_m1c_5) | (IsNaN_6U_10U_2_land_2_lpi_1_dfm_24 & inp_lookup_if_and_m1c_3);
  assign inp_lookup_if_and_15_rgt = inp_lookup_if_unequal_tmp_1_mx0w0 & and_1944_m1c;
  assign and_1945_rgt = or_11_cse & (~ (chn_inp_in_crt_sva_10_739_736_1[1]));
  assign inp_lookup_if_or_rgt = ((~ FpAdd_6U_10U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0)
      & inp_lookup_if_and_m1c_2) | (IsNaN_6U_10U_3_land_1_lpi_1_dfm_6 & inp_lookup_if_and_m1c_1);
  assign inp_lookup_if_or_1_rgt = (FpAdd_6U_10U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0
      & inp_lookup_if_and_m1c_2) | (IsNaN_6U_10U_2_land_1_lpi_1_dfm_24 & inp_lookup_if_and_m1c);
  assign inp_lookup_if_and_7_rgt = inp_lookup_if_unequal_tmp_1_mx0w0 & and_dcpl_1473;
  assign and_1947_rgt = or_11_cse & (~ (chn_inp_in_crt_sva_10_739_736_1[0]));
  assign FpAdd_6U_10U_and_35_cse = core_wen & ((or_dcpl_280 & main_stage_v_10 & (cfg_precision_1_sva_st_87==2'b10)
      & and_dcpl_1473) | and_dcpl_1481);
  assign FpAdd_6U_10U_and_37_cse = core_wen & ((or_dcpl_283 & and_dcpl_1484 & or_11_cse
      & (chn_inp_in_crt_sva_10_739_736_1[1])) | and_dcpl_1488);
  assign FpAdd_6U_10U_and_39_cse = core_wen & ((or_dcpl_286 & main_stage_v_10 & (cfg_precision_1_sva_st_113==2'b10)
      & or_11_cse & (chn_inp_in_crt_sva_10_739_736_1[2])) | and_dcpl_1497);
  assign nor_268_cse = ~(FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_3 | (~ inp_lookup_2_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs));
  assign nor_267_cse = ~(FpMul_6U_10U_2_lor_7_lpi_1_dfm_5 | (~ inp_lookup_2_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2));
  assign nor_266_cse = ~((chn_inp_in_crt_sva_2_739_736_1[1]) | (cfg_precision_1_sva_st_91!=2'b10));
  assign and_1975_rgt = and_dcpl_423 & (~(IsNaN_6U_10U_7_land_2_lpi_1_dfm_5 | (chn_inp_in_crt_sva_2_739_736_1[1])))
      & and_dcpl_419;
  assign and_1978_rgt = and_dcpl_423 & IsNaN_6U_10U_7_land_2_lpi_1_dfm_5 & (~ (chn_inp_in_crt_sva_2_739_736_1[1]))
      & and_dcpl_419;
  assign and_1982_rgt = (~ IsNaN_6U_10U_7_land_lpi_1_dfm_5) & (cfg_precision_1_sva_st_91[1])
      & and_dcpl_1504 & and_dcpl_419;
  assign and_1985_rgt = IsNaN_6U_10U_7_land_lpi_1_dfm_5 & (cfg_precision_1_sva_st_91[1])
      & and_dcpl_1504 & and_dcpl_419;
  assign and_2012_rgt = or_dcpl_818 & or_11_cse;
  assign and_3150_nl = (~((~ IsNaN_8U_23U_nor_tmp) & (chn_inp_in_rsci_d_mxwt[510:503]==8'b11111111)))
      & (chn_inp_in_rsci_d_mxwt[736]) & (cfg_precision_rsci_d==2'b10) & chn_inp_in_rsci_bawt;
  assign nor_1025_nl = ~((~ main_stage_v_1) | (~ (chn_inp_in_crt_sva_1_739_395_1[341]))
      | IsNaN_8U_23U_land_1_lpi_1_dfm_st_3 | (cfg_precision_1_sva_st_90!=2'b10));
  assign mux_1325_nl = MUX_s_1_2_2((nor_1025_nl), (and_3150_nl), or_11_cse);
  assign IsNaN_8U_23U_1_and_cse = core_wen & (~ and_dcpl_78) & (mux_1325_nl);
  assign and_3149_cse = or_5882_cse & FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_6_1_1
      & FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_6_0_1 & (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_9==4'b1111);
  assign and_2013_rgt = ((FpFractionToFloat_35U_6U_10U_1_mux_tmp!=5'b11111) | IsNaN_6U_10U_6_nor_tmp
      | (~ inp_lookup_1_FpMantRNE_36U_11U_1_else_and_svs_2) | (~((IntLeadZero_35U_1_leading_sign_35_0_rtn_1_sva_2[5])
      & FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_st_2))) & and_dcpl_393;
  assign and_2022_rgt = and_dcpl_393 & and_dcpl_1545 & and_dcpl_1541 & (~ IsNaN_6U_10U_6_nor_tmp)
      & inp_lookup_1_FpMantRNE_36U_11U_1_else_and_svs_2 & (IntLeadZero_35U_1_leading_sign_35_0_rtn_1_sva_2[5])
      & FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_st_2;
  assign and_2023_rgt = ((FpFractionToFloat_35U_6U_10U_1_mux_40_tmp!=5'b11111) |
      IsNaN_6U_10U_6_nor_1_tmp | (~ (IntLeadZero_35U_1_leading_sign_35_0_rtn_2_sva_2[5]))
      | (~(inp_lookup_2_FpMantRNE_36U_11U_1_else_and_svs_2 & FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_st_2)))
      & and_dcpl_401;
  assign and_2033_rgt = and_dcpl_1556 & or_11_cse & (FpFractionToFloat_35U_6U_10U_1_mux_40_tmp[4:3]==2'b11)
      & (~ IsNaN_6U_10U_6_nor_1_tmp) & (IntLeadZero_35U_1_leading_sign_35_0_rtn_2_sva_2[5])
      & inp_lookup_2_FpMantRNE_36U_11U_1_else_and_svs_2 & (~ (chn_inp_in_crt_sva_1_739_395_1[342]))
      & FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_st_2;
  assign nor_1017_cse = ~(IsNaN_6U_10U_7_land_3_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_14);
  assign and_2034_rgt = ((~((FpFractionToFloat_35U_6U_10U_1_mux_41_tmp[4]) & (FpFractionToFloat_35U_6U_10U_1_mux_41_tmp[2])
      & (FpFractionToFloat_35U_6U_10U_1_mux_41_tmp[0]))) | (~(inp_lookup_3_FpMantRNE_36U_11U_1_else_and_svs_2
      & FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_st_2)) | (~((IntLeadZero_35U_1_leading_sign_35_0_rtn_3_sva_2[5])
      & (FpFractionToFloat_35U_6U_10U_1_mux_41_tmp[1]))) | (~ (FpFractionToFloat_35U_6U_10U_1_mux_41_tmp[3]))
      | IsNaN_6U_10U_6_nor_2_tmp) & and_dcpl_409;
  assign and_2043_rgt = and_dcpl_409 & and_dcpl_1566 & FpFractionToFloat_35U_6U_10U_1_and_2_cse
      & (IntLeadZero_35U_1_leading_sign_35_0_rtn_3_sva_2[5]) & (FpFractionToFloat_35U_6U_10U_1_mux_41_tmp[1])
      & (FpFractionToFloat_35U_6U_10U_1_mux_41_tmp[3]) & (~ IsNaN_6U_10U_6_nor_2_tmp);
  assign and_2044_rgt = ((FpFractionToFloat_35U_6U_10U_1_mux_42_tmp!=5'b11111) |
      IsNaN_6U_10U_6_nor_3_tmp | (~ inp_lookup_4_FpMantRNE_36U_11U_1_else_and_svs_2)
      | (~((IntLeadZero_35U_1_leading_sign_35_0_rtn_sva_2[5]) & FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2)))
      & and_dcpl_415;
  assign and_2054_rgt = and_dcpl_1577 & or_11_cse & (FpFractionToFloat_35U_6U_10U_1_mux_42_tmp[4:3]==2'b11)
      & (~ IsNaN_6U_10U_6_nor_3_tmp) & (~ (chn_inp_in_crt_sva_1_739_395_1[344]))
      & inp_lookup_4_FpMantRNE_36U_11U_1_else_and_svs_2 & (IntLeadZero_35U_1_leading_sign_35_0_rtn_sva_2[5])
      & FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2;
  assign and_2058_nl = and_dcpl_423 & and_dcpl_428 & IsNaN_6U_10U_7_land_1_lpi_1_dfm_5
      & main_stage_v_2 & or_11_cse;
  assign and_2060_nl = and_dcpl_423 & and_dcpl_433 & and_dcpl_419;
  assign or_5132_nl = (~ main_stage_v_2) | IsNaN_6U_10U_7_land_1_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_14
      | (chn_inp_in_crt_sva_2_739_736_1[0]) | (cfg_precision_1_sva_st_91!=2'b10);
  assign mux_1948_nl = MUX_s_1_2_2(or_tmp_4282, (or_5132_nl), or_11_cse);
  assign or_5136_nl = IsNaN_6U_10U_7_land_1_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_14
      | (chn_inp_in_crt_sva_2_739_736_1[0]) | (cfg_precision_1_sva_st_91!=2'b10);
  assign mux_1949_nl = MUX_s_1_2_2(or_tmp_4282, (or_5136_nl), or_11_cse);
  assign or_5554_nl = ((~ (mux_1948_nl)) & (fsm_output[1])) | ((~ (mux_1949_nl))
      & main_stage_v_2);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_mux1h_11_rgt = MUX1HOT_v_10_4_2(({reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_7_itm
      , reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_7_1_itm}), FpFractionToFloat_35U_6U_10U_1_o_mant_1_lpi_1_dfm_8,
      FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_3_mx0w0, ({4'b0 , FpMul_6U_10U_2_else_2_else_ac_int_cctor_1_sva_mx0w0}),
      {(and_2058_nl) , (and_2060_nl) , and_dcpl_458 , (or_5554_nl)});
  assign or_5800_cse = (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10) |
      (chn_inp_in_crt_sva_2_739_736_1[0]);
  assign and_2065_rgt = and_dcpl_423 & and_dcpl_468 & and_dcpl_1588;
  assign and_2067_rgt = and_dcpl_423 & and_dcpl_471 & and_dcpl_419;
  assign and_2069_rgt = and_dcpl_423 & and_dcpl_465 & and_dcpl_1588;
  assign and_2073_rgt = and_dcpl_423 & and_dcpl_504 & and_dcpl_1596;
  assign and_2076_rgt = and_dcpl_423 & IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_14 & main_stage_v_2
      & and_dcpl_524;
  assign and_2078_rgt = and_dcpl_423 & nor_1017_cse & and_dcpl_1596;
  assign and_2082_nl = and_dcpl_539 & and_dcpl_423 & (~ (chn_inp_in_crt_sva_2_739_736_1[3]))
      & main_stage_v_2 & or_11_cse;
  assign and_2085_nl = IsNaN_6U_10U_2_land_lpi_1_dfm_st_14 & (cfg_precision_1_sva_st_91[1])
      & and_dcpl_1504 & and_dcpl_419;
  assign nor_nl = ~((~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[3]) | (cfg_precision_1_sva_st_91!=2'b10)
      | IsNaN_6U_10U_7_land_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_lpi_1_dfm_st_14);
  assign nor_1787_nl = ~((~ main_stage_v_3) | IsNaN_6U_10U_7_land_lpi_1_dfm_6 | IsNaN_6U_10U_6_land_lpi_1_dfm_5
      | (chn_inp_in_crt_sva_3_739_736_1[3]) | (cfg_precision_1_sva_st_80!=2'b10));
  assign mux_1953_nl = MUX_s_1_2_2((nor_1787_nl), (nor_nl), or_11_cse);
  assign or_5558_nl = ((mux_1953_nl) & (fsm_output[1])) | (and_dcpl_633 & (~ IsNaN_6U_10U_6_land_lpi_1_dfm_5)
      & (~ IsNaN_6U_10U_7_land_lpi_1_dfm_6) & (cfg_precision_1_sva_st_91[0]) & main_stage_v_3
      & and_dcpl_78);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_mux1h_16_rgt = MUX1HOT_v_10_4_2(({reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_7_itm
      , reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_7_1_itm}), FpFractionToFloat_35U_6U_10U_1_o_mant_lpi_1_dfm_8,
      FpMul_6U_10U_2_o_mant_lpi_1_dfm_3_mx0w0, ({4'b0 , FpMul_6U_10U_2_else_2_else_ac_int_cctor_sva_mx0w0}),
      {(and_2082_nl) , (and_2085_nl) , and_dcpl_1007 , (or_5558_nl)});
  assign nor_1800_cse = ~((cfg_precision_1_sva_st_80!=2'b10) | (chn_inp_in_crt_sva_3_739_736_1[3])
      | (~ main_stage_v_3));
  assign or_5809_cse = (~ (cfg_precision_1_sva_st_91[1])) | (chn_inp_in_crt_sva_2_739_736_1[3])
      | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91[0]);
  assign FpMul_6U_10U_1_o_expo_FpMul_6U_10U_1_o_expo_or_7_cse = and_dcpl_1617 | and_dcpl_1619
      | and_dcpl_719;
  assign and_2097_rgt = or_11_cse & (~ IsNaN_6U_10U_8_land_lpi_1_dfm_4);
  assign or_5152_cse = IsNaN_6U_10U_8_land_lpi_1_dfm_4 | (chn_inp_in_crt_sva_5_739_736_1[3]);
  assign FpMul_6U_10U_1_o_expo_FpMul_6U_10U_1_o_expo_or_5_cse = and_dcpl_1624 | and_dcpl_1626
      | and_dcpl_712;
  assign and_2104_rgt = or_11_cse & (~ IsNaN_6U_10U_8_land_3_lpi_1_dfm_4);
  assign or_3167_cse = (cfg_precision_1_sva_st_82!=2'b10) | (~ main_stage_v_5);
  assign and_1185_tmp = or_11_cse & IsNaN_8U_23U_3_land_3_lpi_1_dfm_6;
  assign mux_1958_m1c = MUX_s_1_2_2((chn_inp_in_crt_sva_6_739_736_1[2]), (chn_inp_in_crt_sva_5_739_736_1[2]),
      or_11_cse);
  assign FpMul_6U_10U_1_o_expo_FpMul_6U_10U_1_o_expo_or_3_cse = and_dcpl_1632 | and_dcpl_1634
      | and_dcpl_701;
  assign and_2112_rgt = or_11_cse & (~ IsNaN_6U_10U_8_land_2_lpi_1_dfm_4);
  assign or_5154_cse = IsNaN_6U_10U_8_land_2_lpi_1_dfm_4 | (chn_inp_in_crt_sva_5_739_736_1[1]);
  assign FpMul_6U_10U_1_o_expo_FpMul_6U_10U_1_o_expo_or_1_cse = and_dcpl_1639 | and_dcpl_1641
      | and_dcpl_690;
  assign and_2119_rgt = or_11_cse & (~ IsNaN_6U_10U_8_land_1_lpi_1_dfm_6);
  assign or_5155_cse = IsNaN_6U_10U_8_land_1_lpi_1_dfm_6 | (chn_inp_in_crt_sva_5_739_736_1[0]);
  assign IsNaN_6U_10U_2_aelse_and_30_cse = core_wen & (~ and_dcpl_78) & (~ mux_854_cse);
  assign mux_1372_nl = MUX_s_1_2_2(or_tmp_2924, or_tmp_3224, or_11_cse);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_8_cse = core_wen & (~ and_dcpl_78)
      & (~ (mux_1372_nl));
  assign mux_1373_nl = MUX_s_1_2_2(or_tmp_2935, or_tmp_3227, or_11_cse);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_9_cse = core_wen & (~ and_dcpl_78)
      & (~ (mux_1373_nl));
  assign mux_1374_nl = MUX_s_1_2_2(or_tmp_2953, or_tmp_3230, or_11_cse);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_10_cse = core_wen & (~ and_dcpl_78)
      & (~ (mux_1374_nl));
  assign mux_1375_nl = MUX_s_1_2_2(or_tmp_2974, or_tmp_3233, or_11_cse);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_11_cse = core_wen & (~ and_dcpl_78)
      & (~ (mux_1375_nl));
  assign and_2125_rgt = or_11_cse & (chn_inp_in_crt_sva_9_739_736_1[3]);
  assign and_2130_rgt = or_11_cse & (chn_inp_in_crt_sva_9_739_736_1[2]);
  assign and_2135_rgt = or_11_cse & (chn_inp_in_crt_sva_9_739_736_1[1]);
  assign and_2140_rgt = or_11_cse & (chn_inp_in_crt_sva_9_739_736_1[0]);
  assign mux_1376_nl = MUX_s_1_2_2(or_tmp_2986, or_tmp_3235, or_11_cse);
  assign inp_lookup_else_and_20_cse = core_wen & (~ and_dcpl_78) & (~ (mux_1376_nl));
  assign mux_1385_nl = MUX_s_1_2_2(or_tmp_2990, or_tmp_3246, or_11_cse);
  assign inp_lookup_else_and_21_cse = core_wen & (~ and_dcpl_78) & (~ (mux_1385_nl));
  assign mux_1394_nl = MUX_s_1_2_2(or_tmp_2993, or_tmp_3257, or_11_cse);
  assign inp_lookup_else_and_22_cse = core_wen & (~ and_dcpl_78) & (~ (mux_1394_nl));
  assign mux_1403_nl = MUX_s_1_2_2(or_tmp_2997, or_tmp_3268, or_11_cse);
  assign inp_lookup_else_and_23_cse = core_wen & (~ and_dcpl_78) & (~ (mux_1403_nl));
  assign or_3291_cse = (cfg_precision_1_sva_20!=2'b10);
  assign nand_358_cse = ~(main_stage_v_2 & (chn_inp_in_crt_sva_2_739_736_1[1]) &
      (cfg_precision_1_sva_st_91==2'b10));
  assign or_3384_cse = (cfg_precision_1_sva_st_82!=2'b10);
  assign or_3379_cse = (cfg_precision_1_sva_st_81!=2'b10);
  assign nor_959_cse = ~((chn_inp_in_crt_sva_4_739_736_1[3]) | (cfg_precision_1_sva_st_81[0])
      | not_tmp_1425);
  assign nor_960_cse = ~((cfg_precision_1_sva_st_81[0]) | not_tmp_1425);
  assign nor_962_itm = ~((cfg_precision_1_sva_st_82[0]) | not_tmp_374);
  assign mux_2206_nl = MUX_s_1_2_2(main_stage_v_5, nor_962_itm, or_3384_cse);
  assign mux_1480_cse = MUX_s_1_2_2((mux_2206_nl), main_stage_v_5, chn_inp_in_crt_sva_5_739_736_1[3]);
  assign mux_1476_cse = MUX_s_1_2_2(main_stage_v_4, nor_960_cse, or_3379_cse);
  assign nor_956_cse = ~((cfg_precision_1_sva_st_81!=2'b10));
  assign mux_1483_cse = MUX_s_1_2_2(nor_960_cse, main_stage_v_4, nor_956_cse);
  assign nor_950_cse = ~((chn_inp_in_crt_sva_4_739_736_1[2]) | (cfg_precision_1_sva_st_81[0])
      | not_tmp_1425);
  assign nor_952_cse = ~((chn_inp_in_crt_sva_5_739_736_1[2]) | (cfg_precision_1_sva_st_82[0])
      | not_tmp_374);
  assign mux_2207_nl = MUX_s_1_2_2(main_stage_v_5, nor_962_itm, or_3384_cse);
  assign mux_1493_cse = MUX_s_1_2_2((mux_2207_nl), main_stage_v_5, chn_inp_in_crt_sva_5_739_736_1[2]);
  assign nor_941_cse = ~((chn_inp_in_crt_sva_4_739_736_1[1]) | (cfg_precision_1_sva_st_81[0])
      | not_tmp_1425);
  assign nor_943_cse = ~((chn_inp_in_crt_sva_5_739_736_1[1]) | (cfg_precision_1_sva_st_82[0])
      | not_tmp_374);
  assign mux_2208_nl = MUX_s_1_2_2(main_stage_v_5, nor_962_itm, or_3384_cse);
  assign mux_1506_cse = MUX_s_1_2_2((mux_2208_nl), main_stage_v_5, chn_inp_in_crt_sva_5_739_736_1[1]);
  assign nor_932_cse = ~((chn_inp_in_crt_sva_4_739_736_1[0]) | (cfg_precision_1_sva_st_81[0])
      | not_tmp_1425);
  assign mux_1479_nl = MUX_s_1_2_2(main_stage_v_5, nor_962_itm, or_3384_cse);
  assign mux_1519_cse = MUX_s_1_2_2((mux_1479_nl), main_stage_v_5, chn_inp_in_crt_sva_5_739_736_1[0]);
  assign and_3588_cse = ((FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_22_13_lpi_1_dfm_mx0w1!=10'b0000000000)
      | (FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_9_0_lpi_1_dfm!=10'b0000000000))
      & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_13_1_1;
  assign or_3482_nl = (chn_inp_in_crt_sva_8_739_736_1[3]) | (~ main_stage_v_8) |
      inp_lookup_else_unequal_tmp_55;
  assign mux_1540_nl = MUX_s_1_2_2(or_tmp_3224, (or_3482_nl), or_11_cse);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_12_cse = core_wen & (~ and_dcpl_78)
      & (~ (mux_1540_nl));
  assign or_3484_cse = (cfg_precision_1_sva_18!=2'b10);
  assign or_3489_cse = (cfg_precision_1_sva_19!=2'b10);
  assign nor_1756_nl = ~((cfg_precision_1_sva_st_85[0]) | nand_544_cse);
  assign mux_1541_cse = MUX_s_1_2_2(main_stage_v_8, (nor_1756_nl), or_3484_cse);
  assign and_3587_cse = ((FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_22_13_3_lpi_1_dfm_mx0w1!=10'b0000000000)
      | (FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_9_0_3_lpi_1_dfm!=10'b0000000000))
      & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_13_1_1;
  assign or_3495_nl = (chn_inp_in_crt_sva_8_739_736_1[2]) | (~ main_stage_v_8) |
      inp_lookup_else_unequal_tmp_55;
  assign mux_1548_nl = MUX_s_1_2_2(or_tmp_3227, (or_3495_nl), or_11_cse);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_13_cse = core_wen & (~ and_dcpl_78)
      & (~ (mux_1548_nl));
  assign and_3586_cse = ((FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_22_13_2_lpi_1_dfm_mx0w1!=10'b0000000000)
      | (FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_9_0_2_lpi_1_dfm!=10'b0000000000))
      & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_13_1_1;
  assign or_3508_nl = (chn_inp_in_crt_sva_8_739_736_1[1]) | (~ main_stage_v_8) |
      inp_lookup_else_unequal_tmp_55;
  assign mux_1556_nl = MUX_s_1_2_2(or_tmp_3230, (or_3508_nl), or_11_cse);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_14_cse = core_wen & (~ and_dcpl_78)
      & (~ (mux_1556_nl));
  assign and_3585_cse = ((FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_22_13_1_lpi_1_dfm_mx0w1!=10'b0000000000)
      | (FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_9_0_1_lpi_1_dfm!=10'b0000000000))
      & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_13_1_1;
  assign or_3510_nl = (chn_inp_in_crt_sva_8_739_736_1[0]) | (~ main_stage_v_8) |
      inp_lookup_else_unequal_tmp_55;
  assign mux_1557_nl = MUX_s_1_2_2(or_tmp_3233, (or_3510_nl), or_11_cse);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_15_cse = core_wen & (~ and_dcpl_78)
      & (~ (mux_1557_nl));
  assign mux_1963_cse = MUX_s_1_2_2(inp_lookup_else_unequal_tmp_35, inp_lookup_else_unequal_tmp_55,
      or_11_cse);
  assign IntShiftRight_69U_6U_32U_obits_fixed_mux1h_25_itm = MUX_v_17_2_2(({8'b0
      , (FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_9_0_lpi_1_dfm_2_mx0[9:1])}), (IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_12[17:1]),
      mux_1963_cse);
  assign IntShiftRight_69U_6U_32U_obits_fixed_mux1h_27_itm = MUX_v_17_2_2(({8'b0
      , (FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_9_0_3_lpi_1_dfm_2_mx0[9:1])}), (IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_12[17:1]),
      mux_1963_cse);
  assign IntShiftRight_69U_6U_32U_obits_fixed_mux1h_29_itm = MUX_v_17_2_2(({8'b0
      , (FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_9_0_2_lpi_1_dfm_2_mx0[9:1])}), (IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_12[17:1]),
      mux_1963_cse);
  assign IntShiftRight_69U_6U_32U_obits_fixed_mux1h_31_itm = MUX_v_17_2_2(({8'b0
      , (FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_9_0_1_lpi_1_dfm_2_mx0[9:1])}), (IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_12[17:1]),
      mux_1963_cse);
  assign and_307_cse = (chn_inp_in_crt_sva_8_739_736_1[1]) & main_stage_v_8 & or_3484_cse;
  assign and_2194_rgt = or_11_cse & (~ inp_lookup_else_unequal_tmp_55);
  assign IntShiftRight_69U_6U_32U_obits_fixed_inp_lookup_else_or_7_cse = (or_11_cse
      & inp_lookup_else_unequal_tmp_55) | and_2194_rgt;
  assign and_3113_cse = (chn_inp_in_crt_sva_9_739_736_1[0]) & main_stage_v_9;
  assign and_3112_cse = (chn_inp_in_crt_sva_9_739_736_1[3]) & main_stage_v_9;
  assign and_3111_cse = (chn_inp_in_crt_sva_9_739_736_1[1]) & main_stage_v_9;
  assign and_3110_cse = (chn_inp_in_crt_sva_9_739_736_1[2]) & main_stage_v_9;
  assign FpAdd_6U_10U_and_41_cse = core_wen & ((or_dcpl_289 & main_stage_v_10 & (cfg_precision_1_sva_st_125==2'b10)
      & and_dcpl_1722) | and_dcpl_1731);
  assign nand_332_cse = ~(main_stage_v_8 & inp_lookup_else_unequal_tmp_55);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_cse = core_wen & (~(or_dcpl_631
      | (fsm_output[0])));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_3_cse = core_wen & (~(or_dcpl_634
      | (fsm_output[0])));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_6_cse = core_wen & (~(or_dcpl_637
      | (fsm_output[0])));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_9_cse = core_wen & (~(or_dcpl_640
      | (fsm_output[0])));
  assign or_3558_cse = (cfg_precision_1_sva_17!=2'b10);
  assign and_312_cse = main_stage_v_7 & (chn_inp_in_crt_sva_7_739_736_1[1]) & or_3558_cse;
  assign IsZero_6U_10U_1_and_12_cse = core_wen & (~ and_dcpl_78) & (~ mux_115_itm);
  assign nor_905_cse = ~((~ (inp_lookup_1_FpMul_6U_10U_1_p_mant_p1_mul_tmp[21]))
      | inp_lookup_1_FpMul_6U_10U_1_else_2_else_if_if_acc_1_itm_5_1);
  assign nor_908_cse = ~((~ FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_9_1)
      | inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5);
  assign and_2284_rgt = (((~ IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_15) & IsNaN_6U_10U_5_land_1_lpi_1_dfm_5)
      | (chn_inp_in_crt_sva_3_739_736_1[0])) & or_11_cse;
  assign and_2287_rgt = (~(IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_15 | IsNaN_6U_10U_5_land_1_lpi_1_dfm_5
      | (chn_inp_in_crt_sva_3_739_736_1[0]))) & or_11_cse;
  assign and_2289_rgt = IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_15 & (~ (chn_inp_in_crt_sva_3_739_736_1[0]))
      & or_11_cse;
  assign nor_898_cse = ~((~ (inp_lookup_2_FpMul_6U_10U_1_p_mant_p1_mul_tmp[21]))
      | inp_lookup_2_FpMul_6U_10U_1_else_2_else_if_if_acc_1_itm_5_1);
  assign nor_901_cse = ~((~ FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_9_1)
      | inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5);
  assign and_2291_rgt = (((~ IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_15) & IsNaN_6U_10U_5_land_2_lpi_1_dfm_5)
      | (chn_inp_in_crt_sva_3_739_736_1[1])) & or_11_cse;
  assign and_2294_rgt = (~(IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_15 | IsNaN_6U_10U_5_land_2_lpi_1_dfm_5
      | (chn_inp_in_crt_sva_3_739_736_1[1]))) & or_11_cse;
  assign and_2296_rgt = IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_15 & (~ (chn_inp_in_crt_sva_3_739_736_1[1]))
      & or_11_cse;
  assign nor_894_cse = ~((~ FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_9_1)
      | inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4);
  assign nor_572_cse = ~(FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_3 | (~ inp_lookup_4_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs));
  assign and_2298_rgt = (((~ IsNaN_6U_10U_2_land_lpi_1_dfm_st_15) & IsNaN_6U_10U_5_land_lpi_1_dfm_5)
      | (chn_inp_in_crt_sva_3_739_736_1[3])) & or_11_cse;
  assign and_2301_rgt = (~((chn_inp_in_crt_sva_3_739_736_1[3]) | IsNaN_6U_10U_2_land_lpi_1_dfm_st_15
      | IsNaN_6U_10U_5_land_lpi_1_dfm_5)) & or_11_cse;
  assign and_2303_rgt = (~ (chn_inp_in_crt_sva_3_739_736_1[3])) & IsNaN_6U_10U_2_land_lpi_1_dfm_st_15
      & or_11_cse;
  assign or_5766_rgt = ((chn_inp_in_crt_sva_4_739_736_1[0]) & IsNaN_6U_10U_5_land_1_lpi_1_dfm_6
      & or_11_cse) | (FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5 & and_m1c_3);
  assign or_5767_rgt = ((~ FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5) & and_m1c_3)
      | (FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_4 & and_2307_m1c);
  assign or_5764_rgt = (IsNaN_6U_10U_5_land_2_lpi_1_dfm_6 & (chn_inp_in_crt_sva_4_739_736_1[1])
      & or_11_cse) | (FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5 & and_m1c_2);
  assign or_5765_rgt = ((~ FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5) & and_m1c_2)
      | (FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_4 & and_2311_m1c);
  assign or_5762_rgt = ((chn_inp_in_crt_sva_4_739_736_1[2]) & IsNaN_6U_10U_5_land_3_lpi_1_dfm_6
      & or_11_cse) | (FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5 & and_m1c_1);
  assign or_5763_rgt = ((~ FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5) & and_m1c_1)
      | (FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_4 & and_2315_m1c);
  assign or_5760_rgt = ((chn_inp_in_crt_sva_4_739_736_1[3]) & FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_4
      & or_11_cse) | (FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5 & and_m1c);
  assign or_5761_rgt = ((~ FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5) & and_m1c)
      | (IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0 & and_2319_m1c);
  assign and_2320_cse = or_3384_cse & or_11_cse;
  assign or_3716_cse = (chn_inp_in_crt_sva_5_739_736_1[3]) | (~ main_stage_v_5);
  assign IntShiftRight_69U_6U_32U_obits_fixed_or_6_rgt = ((~ FpAdd_6U_10U_1_is_a_greater_lor_lpi_1_dfm_1_mx0w0)
      & IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_7) | (IsNaN_6U_10U_9_land_lpi_1_dfm_6
      & IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_6);
  assign IntShiftRight_69U_6U_32U_obits_fixed_or_7_rgt = (FpAdd_6U_10U_1_is_a_greater_lor_lpi_1_dfm_1_mx0w0
      & IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_7) | (IsNaN_6U_10U_8_land_lpi_1_dfm_4
      & and_2321_m1c);
  assign or_3718_cse = (chn_inp_in_crt_sva_5_739_736_1[2]) | (~ main_stage_v_5);
  assign IntShiftRight_69U_6U_32U_obits_fixed_or_4_rgt = ((~ FpAdd_6U_10U_1_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0)
      & IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_5) | (IsNaN_6U_10U_9_land_3_lpi_1_dfm_6
      & IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_4);
  assign IntShiftRight_69U_6U_32U_obits_fixed_or_5_rgt = (FpAdd_6U_10U_1_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0
      & IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_5) | (IsNaN_6U_10U_8_land_3_lpi_1_dfm_4
      & and_2321_m1c);
  assign or_3720_cse = (chn_inp_in_crt_sva_5_739_736_1[1]) | (~ main_stage_v_5);
  assign IntShiftRight_69U_6U_32U_obits_fixed_or_2_rgt = ((~ FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0)
      & IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_3) | (IsNaN_6U_10U_9_land_2_lpi_1_dfm_6
      & IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_2);
  assign IntShiftRight_69U_6U_32U_obits_fixed_or_3_rgt = (FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0
      & IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_3) | (IsNaN_6U_10U_8_land_2_lpi_1_dfm_4
      & and_2321_m1c);
  assign or_3722_cse = (chn_inp_in_crt_sva_5_739_736_1[0]) | (~ main_stage_v_5);
  assign IntShiftRight_69U_6U_32U_obits_fixed_or_rgt = ((~ FpAdd_6U_10U_1_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0)
      & IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_1) | (IsNaN_6U_10U_9_land_1_lpi_1_dfm_6
      & IntShiftRight_69U_6U_32U_obits_fixed_and_m1c);
  assign IntShiftRight_69U_6U_32U_obits_fixed_or_1_rgt = (FpAdd_6U_10U_1_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0
      & IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_1) | (IsNaN_6U_10U_8_land_1_lpi_1_dfm_6
      & and_2321_m1c);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_100_cse = core_wen & (and_dcpl_1853
      | and_dcpl_1854) & mux_tmp_6;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_103_cse = core_wen & (and_dcpl_1856
      | and_dcpl_1857) & mux_tmp_6;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_106_cse = core_wen & (and_dcpl_1859
      | and_dcpl_1860) & mux_tmp_6;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_109_cse = core_wen & (and_dcpl_1862
      | and_dcpl_1863) & mux_tmp_6;
  assign nor_884_cse = ~((~ IsNaN_6U_10U_5_land_1_lpi_1_dfm_5) | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_15);
  assign nor_880_cse = ~((~ IsNaN_6U_10U_5_land_2_lpi_1_dfm_5) | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_15);
  assign nor_584_cse = ~(inp_lookup_2_FpMul_6U_10U_1_oelse_1_acc_itm_7_1 | FpMul_6U_10U_1_if_2_FpMul_6U_10U_1_if_2_or_2_tmp
      | (~ inp_lookup_2_FpMul_6U_10U_1_else_2_if_acc_itm_6_1));
  assign nor_875_cse = ~((~ IsNaN_6U_10U_5_land_lpi_1_dfm_5) | IsNaN_6U_10U_2_land_lpi_1_dfm_st_15);
  assign nor_586_cse = ~(inp_lookup_4_FpMul_6U_10U_1_oelse_1_acc_itm_7_1 | FpMul_6U_10U_1_if_2_FpMul_6U_10U_1_if_2_or_6_tmp
      | (~ inp_lookup_4_FpMul_6U_10U_1_else_2_if_acc_itm_6_1));
  assign or_3779_cse = (~ inp_lookup_4_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs)
      | FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_3;
  assign and_2342_rgt = (~ IsNaN_6U_10U_5_land_1_lpi_1_dfm_5) & (~ (chn_inp_in_crt_sva_3_739_736_1[0]))
      & or_11_cse;
  assign and_2345_rgt = and_dcpl_597 & or_11_cse;
  assign and_2348_rgt = and_dcpl_627 & or_11_cse;
  assign nor_605_cse = ~((~ inp_lookup_4_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp)
      | FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_3_itm_23_1);
  assign or_3850_cse = (~ main_stage_v_4) | (cfg_precision_1_sva_st_81!=2'b10);
  assign and_2350_rgt = and_dcpl_642 & or_11_cse;
  assign and_2351_rgt = and_dcpl_645 & or_11_cse;
  assign or_3885_cse = (~ IsNaN_6U_10U_8_land_1_lpi_1_dfm_6) | (~ main_stage_v_5)
      | (chn_inp_in_crt_sva_5_739_736_1[0]);
  assign nor_623_cse = ~((cfg_precision_1_sva_st_82!=2'b10));
  assign or_3913_cse = (~ IsNaN_6U_10U_8_land_2_lpi_1_dfm_4) | (~ main_stage_v_5)
      | (chn_inp_in_crt_sva_5_739_736_1[1]);
  assign or_3941_cse = (~ IsNaN_6U_10U_8_land_3_lpi_1_dfm_4) | (~ main_stage_v_5)
      | (chn_inp_in_crt_sva_5_739_736_1[2]);
  assign or_3969_cse = (~ IsNaN_6U_10U_8_land_lpi_1_dfm_4) | (~ main_stage_v_5) |
      (chn_inp_in_crt_sva_5_739_736_1[3]);
  assign FpAdd_8U_23U_o_sign_and_cse = core_wen & (~ and_dcpl_78);
  assign and_348_cse = FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_7_1_1
      & FpAdd_8U_23U_o_sign_3_lpi_1_dfm_7 & inp_lookup_3_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_tmp
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_9==4'b1111) & (IsNaN_6U_10U_4_nor_2_tmp
      | (~(inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_6_5_1 & (inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_6_4_0_1==5'b11111)
      & IsNaN_8U_23U_land_3_lpi_1_dfm_st_4)));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_cse = core_wen & (~(or_dcpl_630
      | and_dcpl_78 | (~ (chn_inp_in_rsci_d_mxwt[737])) | (fsm_output[0])));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_3_cse = core_wen & (~(or_dcpl_630
      | and_dcpl_78 | (~ (chn_inp_in_rsci_d_mxwt[739])) | (fsm_output[0])));
  assign and_2358_rgt = and_dcpl_1852 & or_11_cse & IsDenorm_5U_10U_or_tmp & (chn_inp_in_rsci_d_mxwt[410:406]==5'b11111);
  assign and_2359_rgt = or_dcpl_985 & and_dcpl_1853;
  assign and_2367_rgt = and_dcpl_1060 & (cfg_precision_rsci_d[1]) & (chn_inp_in_rsci_d_mxwt[737])
      & (chn_inp_in_rsci_d_mxwt[422]) & (chn_inp_in_rsci_d_mxwt[423]) & (chn_inp_in_rsci_d_mxwt[424])
      & (chn_inp_in_rsci_d_mxwt[425]) & (chn_inp_in_rsci_d_mxwt[426]) & IsDenorm_5U_10U_or_1_tmp;
  assign and_2368_rgt = or_dcpl_990 & and_dcpl_1856;
  assign and_2375_rgt = and_dcpl_1858 & or_11_cse & (chn_inp_in_rsci_d_mxwt[442])
      & (chn_inp_in_rsci_d_mxwt[441]) & (chn_inp_in_rsci_d_mxwt[438]) & (chn_inp_in_rsci_d_mxwt[440])
      & IsDenorm_5U_10U_or_2_tmp & (chn_inp_in_rsci_d_mxwt[439]);
  assign and_2376_rgt = or_dcpl_995 & and_dcpl_1859;
  assign and_2384_rgt = and_dcpl_1060 & (cfg_precision_rsci_d[1]) & (chn_inp_in_rsci_d_mxwt[739])
      & (chn_inp_in_rsci_d_mxwt[454]) & (chn_inp_in_rsci_d_mxwt[455]) & (chn_inp_in_rsci_d_mxwt[456])
      & (chn_inp_in_rsci_d_mxwt[457]) & (chn_inp_in_rsci_d_mxwt[458]) & IsDenorm_5U_10U_or_3_tmp;
  assign and_2385_rgt = or_dcpl_1000 & and_dcpl_1862;
  assign IntSaturation_51U_32U_o_IntSaturation_51U_32U_o_nor_rgt = ~(inp_lookup_4_IntSaturation_51U_32U_else_if_acc_itm_2_1
      | inp_lookup_4_IntSaturation_51U_32U_if_acc_itm_2_1 | and_dcpl_78);
  assign IntSaturation_51U_32U_and_7_rgt = inp_lookup_4_IntSaturation_51U_32U_else_if_acc_itm_2_1
      & (~ inp_lookup_4_IntSaturation_51U_32U_if_acc_itm_2_1) & (~ and_dcpl_78);
  assign IntSaturation_51U_32U_o_and_7_rgt = inp_lookup_4_IntSaturation_51U_32U_if_acc_itm_2_1
      & (~ and_dcpl_78);
  assign IntSaturation_51U_32U_o_IntSaturation_51U_32U_o_nor_1_rgt = ~(inp_lookup_3_IntSaturation_51U_32U_else_if_acc_itm_2_1
      | inp_lookup_3_IntSaturation_51U_32U_if_acc_itm_2_1 | and_dcpl_78);
  assign IntSaturation_51U_32U_and_5_rgt = inp_lookup_3_IntSaturation_51U_32U_else_if_acc_itm_2_1
      & (~ inp_lookup_3_IntSaturation_51U_32U_if_acc_itm_2_1) & (~ and_dcpl_78);
  assign IntSaturation_51U_32U_o_and_5_rgt = inp_lookup_3_IntSaturation_51U_32U_if_acc_itm_2_1
      & (~ and_dcpl_78);
  assign IntSaturation_51U_32U_o_IntSaturation_51U_32U_o_nor_2_rgt = ~(inp_lookup_2_IntSaturation_51U_32U_else_if_acc_itm_2_1
      | inp_lookup_2_IntSaturation_51U_32U_if_acc_itm_2_1 | and_dcpl_78);
  assign IntSaturation_51U_32U_and_3_rgt = inp_lookup_2_IntSaturation_51U_32U_else_if_acc_itm_2_1
      & (~ inp_lookup_2_IntSaturation_51U_32U_if_acc_itm_2_1) & (~ and_dcpl_78);
  assign IntSaturation_51U_32U_o_and_3_rgt = inp_lookup_2_IntSaturation_51U_32U_if_acc_itm_2_1
      & (~ and_dcpl_78);
  assign IntSaturation_51U_32U_o_IntSaturation_51U_32U_o_nor_3_rgt = ~(inp_lookup_1_IntSaturation_51U_32U_else_if_acc_itm_2_1
      | inp_lookup_1_IntSaturation_51U_32U_if_acc_itm_2_1 | and_dcpl_78);
  assign IntSaturation_51U_32U_and_1_rgt = inp_lookup_1_IntSaturation_51U_32U_else_if_acc_itm_2_1
      & (~ inp_lookup_1_IntSaturation_51U_32U_if_acc_itm_2_1) & (~ and_dcpl_78);
  assign IntSaturation_51U_32U_o_and_1_rgt = inp_lookup_1_IntSaturation_51U_32U_if_acc_itm_2_1
      & (~ and_dcpl_78);
  assign and_2392_rgt = or_dcpl_1005 & or_11_cse;
  assign and_2399_rgt = or_dcpl_1010 & or_11_cse;
  assign and_2404_rgt = and_dcpl_1927 & and_dcpl_1859;
  assign and_2405_rgt = or_dcpl_818 & and_dcpl_1859;
  assign and_2412_rgt = or_dcpl_1015 & or_11_cse;
  assign and_2414_rgt = IsNaN_8U_23U_land_2_lpi_1_dfm_4 & (chn_inp_in_crt_sva_1_739_395_1[342])
      & or_11_cse;
  assign and_2416_rgt = (~ IsNaN_8U_23U_land_2_lpi_1_dfm_4) & (chn_inp_in_crt_sva_1_739_395_1[342])
      & or_11_cse;
  assign and_2417_rgt = and_dcpl_1217 & and_dcpl_416;
  assign and_2418_rgt = and_dcpl_1219 & and_dcpl_416;
  assign and_2419_rgt = (or_2010_cse | (~ (chn_inp_in_crt_sva_1_739_395_1[344])))
      & or_11_cse;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_6_cse = core_wen & (~(or_dcpl_630
      | and_dcpl_78 | (~ (chn_inp_in_rsci_d_mxwt[736])) | (fsm_output[0])));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_9_cse = core_wen & (~(or_dcpl_630
      | and_dcpl_78 | (~ (chn_inp_in_rsci_d_mxwt[738])) | (fsm_output[0])));
  assign and_2497_rgt = or_2010_cse & (~ (chn_inp_in_crt_sva_1_739_395_1[341])) &
      or_11_cse;
  assign and_2499_rgt = and_4210_cse & (~ or_5873_cse) & and_dcpl_393;
  assign and_2501_rgt = and_4210_cse & or_5873_cse & and_dcpl_393;
  assign and_2503_rgt = or_2010_cse & (~ (chn_inp_in_crt_sva_1_739_395_1[342])) &
      or_11_cse;
  assign and_2505_rgt = and_4210_cse & (~ or_5890_cse) & and_dcpl_401;
  assign and_2507_rgt = and_4210_cse & or_5890_cse & and_dcpl_401;
  assign and_2509_rgt = or_2010_cse & (~ (chn_inp_in_crt_sva_1_739_395_1[343])) &
      or_11_cse;
  assign and_2511_rgt = and_4210_cse & (~ FpMul_6U_10U_2_if_2_FpMul_6U_10U_2_if_2_or_5_tmp)
      & and_dcpl_409;
  assign and_2513_rgt = and_4210_cse & FpMul_6U_10U_2_if_2_FpMul_6U_10U_2_if_2_or_5_tmp
      & and_dcpl_409;
  assign and_2515_rgt = or_2010_cse & (~ (chn_inp_in_crt_sva_1_739_395_1[344])) &
      or_11_cse;
  assign and_2517_rgt = and_4210_cse & (~ FpMul_6U_10U_2_if_2_FpMul_6U_10U_2_if_2_or_7_tmp)
      & and_dcpl_415;
  assign and_2519_rgt = and_4210_cse & FpMul_6U_10U_2_if_2_FpMul_6U_10U_2_if_2_or_7_tmp
      & and_dcpl_415;
  assign nl_inp_lookup_1_else_else_a0_acc_nl = ({1'b1 , (~ (chn_inp_in_rsci_d_mxwt[162:128]))})
      + 36'b100000000000000000000000000000000001;
  assign inp_lookup_1_else_else_a0_acc_nl = nl_inp_lookup_1_else_else_a0_acc_nl[35:0];
  assign nl_inp_lookup_if_else_ob_acc_8_nl = ({1'b1 , (~ (chn_inp_in_rsci_d_mxwt[639:609]))})
      + 32'b1;
  assign inp_lookup_if_else_ob_acc_8_nl = nl_inp_lookup_if_else_ob_acc_8_nl[31:0];
  assign nl_inp_lookup_if_else_ob_acc_nl = conv_s2s_32_33(chn_inp_in_rsci_d_mxwt[31:0])
      + conv_s2s_32_33(~ (chn_inp_in_rsci_d_mxwt[511:480]));
  assign inp_lookup_if_else_ob_acc_nl = nl_inp_lookup_if_else_ob_acc_nl[32:0];
  assign nl_inp_lookup_1_if_else_a_acc_nl = conv_s2u_33_34({(inp_lookup_if_else_ob_acc_8_nl)
      , (~ (chn_inp_in_rsci_d_mxwt[608]))}) + conv_s2u_33_34(inp_lookup_if_else_ob_acc_nl);
  assign inp_lookup_1_if_else_a_acc_nl = nl_inp_lookup_1_if_else_a_acc_nl[33:0];
  assign and_2521_nl = or_2_cse & (~ (chn_inp_in_rsci_d_mxwt[736])) & or_11_cse;
  assign mux_1972_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_1_739_395_1[341]), (chn_inp_in_rsci_d_mxwt[736]),
      or_11_cse);
  assign mux_1973_nl = MUX_s_1_2_2(or_dcpl_897, or_dcpl_44, or_11_cse);
  assign inp_lookup_else_else_a0_mux1h_rgt = MUX1HOT_v_36_3_2((inp_lookup_1_else_else_a0_acc_nl),
      ({2'b0 , (inp_lookup_1_if_else_a_acc_nl)}), ({1'b0 , inp_lookup_else_if_a0_frac_1_sva_mx0w0}),
      {(and_2521_nl) , (mux_1972_nl) , (~ (mux_1973_nl))});
  assign nor_1798_cse = ~((cfg_precision_rsci_d!=2'b10));
  assign nl_inp_lookup_2_else_else_a0_acc_nl = ({1'b1 , (~ (chn_inp_in_rsci_d_mxwt[197:163]))})
      + 36'b100000000000000000000000000000000001;
  assign inp_lookup_2_else_else_a0_acc_nl = nl_inp_lookup_2_else_else_a0_acc_nl[35:0];
  assign nl_inp_lookup_if_else_ob_acc_9_nl = ({1'b1 , (~ (chn_inp_in_rsci_d_mxwt[671:641]))})
      + 32'b1;
  assign inp_lookup_if_else_ob_acc_9_nl = nl_inp_lookup_if_else_ob_acc_9_nl[31:0];
  assign nl_inp_lookup_if_else_ob_acc_2_nl = conv_s2s_32_33(chn_inp_in_rsci_d_mxwt[63:32])
      + conv_s2s_32_33(~ (chn_inp_in_rsci_d_mxwt[543:512]));
  assign inp_lookup_if_else_ob_acc_2_nl = nl_inp_lookup_if_else_ob_acc_2_nl[32:0];
  assign nl_inp_lookup_2_if_else_a_acc_nl = conv_s2u_33_34({(inp_lookup_if_else_ob_acc_9_nl)
      , (~ (chn_inp_in_rsci_d_mxwt[640]))}) + conv_s2u_33_34(inp_lookup_if_else_ob_acc_2_nl);
  assign inp_lookup_2_if_else_a_acc_nl = nl_inp_lookup_2_if_else_a_acc_nl[33:0];
  assign and_2524_nl = or_2_cse & (~ (chn_inp_in_rsci_d_mxwt[737])) & or_11_cse;
  assign mux_1974_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_1_739_395_1[342]), (chn_inp_in_rsci_d_mxwt[737]),
      or_11_cse);
  assign mux_1975_nl = MUX_s_1_2_2(or_dcpl_903, or_dcpl_80, or_11_cse);
  assign inp_lookup_else_else_a0_mux1h_1_rgt = MUX1HOT_v_36_3_2((inp_lookup_2_else_else_a0_acc_nl),
      ({2'b0 , (inp_lookup_2_if_else_a_acc_nl)}), ({1'b0 , inp_lookup_else_if_a0_frac_2_sva_mx0w0}),
      {(and_2524_nl) , (mux_1974_nl) , (~ (mux_1975_nl))});
  assign nl_inp_lookup_3_else_else_a0_acc_nl = ({1'b1 , (~ (chn_inp_in_rsci_d_mxwt[232:198]))})
      + 36'b100000000000000000000000000000000001;
  assign inp_lookup_3_else_else_a0_acc_nl = nl_inp_lookup_3_else_else_a0_acc_nl[35:0];
  assign nl_inp_lookup_if_else_ob_acc_10_nl = ({1'b1 , (~ (chn_inp_in_rsci_d_mxwt[703:673]))})
      + 32'b1;
  assign inp_lookup_if_else_ob_acc_10_nl = nl_inp_lookup_if_else_ob_acc_10_nl[31:0];
  assign nl_inp_lookup_if_else_ob_acc_4_nl = conv_s2s_32_33(chn_inp_in_rsci_d_mxwt[95:64])
      + conv_s2s_32_33(~ (chn_inp_in_rsci_d_mxwt[575:544]));
  assign inp_lookup_if_else_ob_acc_4_nl = nl_inp_lookup_if_else_ob_acc_4_nl[32:0];
  assign nl_inp_lookup_3_if_else_a_acc_nl = conv_s2u_33_34({(inp_lookup_if_else_ob_acc_10_nl)
      , (~ (chn_inp_in_rsci_d_mxwt[672]))}) + conv_s2u_33_34(inp_lookup_if_else_ob_acc_4_nl);
  assign inp_lookup_3_if_else_a_acc_nl = nl_inp_lookup_3_if_else_a_acc_nl[33:0];
  assign and_2527_nl = or_2_cse & (~ (chn_inp_in_rsci_d_mxwt[738])) & or_11_cse;
  assign mux_1976_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_1_739_395_1[343]), (chn_inp_in_rsci_d_mxwt[738]),
      or_11_cse);
  assign mux_1977_nl = MUX_s_1_2_2(or_801_cse, or_dcpl_116, or_11_cse);
  assign inp_lookup_else_else_a0_mux1h_2_rgt = MUX1HOT_v_36_3_2((inp_lookup_3_else_else_a0_acc_nl),
      ({2'b0 , (inp_lookup_3_if_else_a_acc_nl)}), ({1'b0 , inp_lookup_else_if_a0_frac_3_sva_mx0w0}),
      {(and_2527_nl) , (mux_1976_nl) , (~ (mux_1977_nl))});
  assign nor_758_cse = ~((chn_inp_in_crt_sva_1_739_395_1[343]) | nor_1336_cse_1);
  assign nl_inp_lookup_4_else_else_a0_acc_nl = ({1'b1 , (~ (chn_inp_in_rsci_d_mxwt[267:233]))})
      + 36'b100000000000000000000000000000000001;
  assign inp_lookup_4_else_else_a0_acc_nl = nl_inp_lookup_4_else_else_a0_acc_nl[35:0];
  assign nl_inp_lookup_if_else_ob_acc_11_nl = ({1'b1 , (~ (chn_inp_in_rsci_d_mxwt[735:705]))})
      + 32'b1;
  assign inp_lookup_if_else_ob_acc_11_nl = nl_inp_lookup_if_else_ob_acc_11_nl[31:0];
  assign nl_inp_lookup_if_else_ob_acc_6_nl = conv_s2s_32_33(chn_inp_in_rsci_d_mxwt[127:96])
      + conv_s2s_32_33(~ (chn_inp_in_rsci_d_mxwt[607:576]));
  assign inp_lookup_if_else_ob_acc_6_nl = nl_inp_lookup_if_else_ob_acc_6_nl[32:0];
  assign nl_inp_lookup_4_if_else_a_acc_nl = conv_s2u_33_34({(inp_lookup_if_else_ob_acc_11_nl)
      , (~ (chn_inp_in_rsci_d_mxwt[704]))}) + conv_s2u_33_34(inp_lookup_if_else_ob_acc_6_nl);
  assign inp_lookup_4_if_else_a_acc_nl = nl_inp_lookup_4_if_else_a_acc_nl[33:0];
  assign and_2530_nl = or_2_cse & (~ (chn_inp_in_rsci_d_mxwt[739])) & or_11_cse;
  assign mux_1978_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_1_739_395_1[344]), (chn_inp_in_rsci_d_mxwt[739]),
      or_11_cse);
  assign mux_1979_nl = MUX_s_1_2_2(or_1970_cse, or_dcpl_152, or_11_cse);
  assign inp_lookup_else_else_a0_mux1h_3_rgt = MUX1HOT_v_36_3_2((inp_lookup_4_else_else_a0_acc_nl),
      ({2'b0 , (inp_lookup_4_if_else_a_acc_nl)}), ({1'b0 , inp_lookup_else_if_a0_frac_sva_mx0w0}),
      {(and_2530_nl) , (mux_1978_nl) , (~ (mux_1979_nl))});
  assign nor_756_cse = ~((chn_inp_in_crt_sva_1_739_395_1[344]) | nor_1336_cse_1);
  assign and_518_nl = and_dcpl_40 & and_dcpl_38 & (fsm_output[1]);
  assign inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_518_nl);
  assign and_522_nl = and_dcpl_40 & or_11_cse & (~ (chn_inp_in_rsci_d_mxwt[736]))
      & (fsm_output[1]);
  assign inp_lookup_1_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_522_nl);
  assign and_524_nl = and_dcpl_40 & and_dcpl_49 & (fsm_output[1]);
  assign inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_524_nl);
  assign and_528_nl = and_dcpl_40 & or_11_cse & (~ (chn_inp_in_rsci_d_mxwt[737]))
      & (fsm_output[1]);
  assign inp_lookup_2_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_528_nl);
  assign and_530_nl = and_dcpl_40 & and_dcpl_57 & (fsm_output[1]);
  assign inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_530_nl);
  assign and_534_nl = and_dcpl_40 & or_11_cse & (~ (chn_inp_in_rsci_d_mxwt[738]))
      & (fsm_output[1]);
  assign inp_lookup_3_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_534_nl);
  assign and_536_nl = and_dcpl_40 & and_dcpl_65 & (fsm_output[1]);
  assign inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_2_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_536_nl);
  assign and_540_nl = and_dcpl_40 & or_11_cse & (~ (chn_inp_in_rsci_d_mxwt[739]))
      & (fsm_output[1]);
  assign inp_lookup_4_NV_NVDLA_SDP_CORE_Y_inp_core_nvdla_float_h_ln433_assert_iExpoWidth_le_oExpoWidth_5_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_540_nl);
  assign IsNaN_8U_23U_nor_tmp = ~((chn_inp_in_rsci_d_mxwt[502:480]!=23'b00000000000000000000000));
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_nl = ({1'b1 , (chn_inp_in_rsci_d_mxwt[502:480])})
      + conv_u2u_23_24(~ (chn_inp_in_rsci_d_mxwt[630:608])) + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_nl[23:0];
  assign nl_FpAdd_8U_23U_is_a_greater_acc_nl = ({1'b1 , (chn_inp_in_rsci_d_mxwt[638:631])})
      + conv_u2u_8_9(~ (chn_inp_in_rsci_d_mxwt[510:503])) + 9'b1;
  assign FpAdd_8U_23U_is_a_greater_acc_nl = nl_FpAdd_8U_23U_is_a_greater_acc_nl[8:0];
  assign FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0 = (~((readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_nl)))
      | ((chn_inp_in_rsci_d_mxwt[510:503]) != (chn_inp_in_rsci_d_mxwt[638:631]))))
      | (readslicef_9_1_8((FpAdd_8U_23U_is_a_greater_acc_nl)));
  assign inp_lookup_else_if_unequal_tmp_mx0w1 = (chn_inp_in_rsci_d_mxwt[162:128]!=35'b00000000000000000000000000000000000);
  assign nl_inp_lookup_else_if_a0_frac_1_sva_mx0w0 = (~ (chn_inp_in_rsci_d_mxwt[162:128]))
      + 35'b1;
  assign inp_lookup_else_if_a0_frac_1_sva_mx0w0 = nl_inp_lookup_else_if_a0_frac_1_sva_mx0w0[34:0];
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_nl
      = ~((chn_inp_in_rsci_d_mxwt[346]) | IsZero_5U_10U_3_land_1_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_mux_2_nl = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_1_sva[4]), IsDenorm_5U_10U_3_land_1_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_3_0_mx0w0 = (FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_mux_2_nl)
      | IsInf_5U_10U_3_land_1_lpi_1_dfm | IsNaN_5U_10U_3_land_1_lpi_1_dfm;
  assign IsZero_5U_10U_3_aelse_not_27_nl = ~ IsZero_5U_10U_3_land_1_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_and_2_nl
      = MUX_v_4_2_2(4'b0000, (chn_inp_in_rsci_d_mxwt[345:342]), (IsZero_5U_10U_3_aelse_not_27_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_mux1h_nl
      = MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_and_2_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_1_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_cse
      , IsDenorm_5U_10U_3_land_1_lpi_1_dfm , IsInf_5U_10U_3_land_1_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_mux1h_nl),
      4'b1111, IsNaN_5U_10U_3_land_1_lpi_1_dfm);
  assign inp_lookup_1_FpMantRNE_36U_11U_1_else_and_tmp = FpMantRNE_36U_11U_1_else_carry_1_sva
      & (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[35:25]==11'b11111111111);
  assign nl_inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_nl =
      conv_u2u_5_6(libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_12[5:1])
      + 6'b110001;
  assign inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_nl = nl_inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_nl[5:0];
  assign inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_itm_5 =
      readslicef_6_1_5((inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_nl));
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_nl = ({1'b1 , (chn_inp_in_rsci_d_mxwt[534:512])})
      + conv_u2u_23_24(~ (chn_inp_in_rsci_d_mxwt[662:640])) + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_nl[23:0];
  assign nl_FpAdd_8U_23U_is_a_greater_acc_1_nl = ({1'b1 , (chn_inp_in_rsci_d_mxwt[670:663])})
      + conv_u2u_8_9(~ (chn_inp_in_rsci_d_mxwt[542:535])) + 9'b1;
  assign FpAdd_8U_23U_is_a_greater_acc_1_nl = nl_FpAdd_8U_23U_is_a_greater_acc_1_nl[8:0];
  assign FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0 = (~((readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_1_nl)))
      | ((chn_inp_in_rsci_d_mxwt[542:535]) != (chn_inp_in_rsci_d_mxwt[670:663]))))
      | (readslicef_9_1_8((FpAdd_8U_23U_is_a_greater_acc_1_nl)));
  assign inp_lookup_else_if_unequal_tmp_1_mx0w1 = (chn_inp_in_rsci_d_mxwt[197:163]!=35'b00000000000000000000000000000000000);
  assign nl_inp_lookup_else_if_a0_frac_2_sva_mx0w0 = (~ (chn_inp_in_rsci_d_mxwt[197:163]))
      + 35'b1;
  assign inp_lookup_else_if_a0_frac_2_sva_mx0w0 = nl_inp_lookup_else_if_a0_frac_2_sva_mx0w0[34:0];
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_1_nl
      = ~((chn_inp_in_rsci_d_mxwt[362]) | IsZero_5U_10U_3_land_2_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_mux_7_nl = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_1_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_2_sva[4]), IsDenorm_5U_10U_3_land_2_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_3_0_mx0w0 = (FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_mux_7_nl)
      | IsInf_5U_10U_3_land_2_lpi_1_dfm | IsNaN_5U_10U_3_land_2_lpi_1_dfm;
  assign IsZero_5U_10U_3_aelse_not_26_nl = ~ IsZero_5U_10U_3_land_2_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_and_5_nl
      = MUX_v_4_2_2(4'b0000, (chn_inp_in_rsci_d_mxwt[361:358]), (IsZero_5U_10U_3_aelse_not_26_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_mux1h_1_nl
      = MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_and_5_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_2_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_1_cse
      , IsDenorm_5U_10U_3_land_2_lpi_1_dfm , IsInf_5U_10U_3_land_2_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_mux1h_1_nl),
      4'b1111, IsNaN_5U_10U_3_land_2_lpi_1_dfm);
  assign inp_lookup_2_FpMantRNE_36U_11U_1_else_and_tmp = FpMantRNE_36U_11U_1_else_carry_2_sva
      & (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[35:25]==11'b11111111111);
  assign nl_inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_nl =
      conv_u2u_5_6(libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_13[5:1])
      + 6'b110001;
  assign inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_nl = nl_inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_nl[5:0];
  assign inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_itm_5 =
      readslicef_6_1_5((inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_nl));
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_nl = ({1'b1 , (chn_inp_in_rsci_d_mxwt[566:544])})
      + conv_u2u_23_24(~ (chn_inp_in_rsci_d_mxwt[694:672])) + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_nl[23:0];
  assign nl_FpAdd_8U_23U_is_a_greater_acc_2_nl = ({1'b1 , (chn_inp_in_rsci_d_mxwt[702:695])})
      + conv_u2u_8_9(~ (chn_inp_in_rsci_d_mxwt[574:567])) + 9'b1;
  assign FpAdd_8U_23U_is_a_greater_acc_2_nl = nl_FpAdd_8U_23U_is_a_greater_acc_2_nl[8:0];
  assign FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0 = (~((readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_2_nl)))
      | ((chn_inp_in_rsci_d_mxwt[574:567]) != (chn_inp_in_rsci_d_mxwt[702:695]))))
      | (readslicef_9_1_8((FpAdd_8U_23U_is_a_greater_acc_2_nl)));
  assign nl_inp_lookup_else_if_a0_frac_3_sva_mx0w0 = (~ (chn_inp_in_rsci_d_mxwt[232:198]))
      + 35'b1;
  assign inp_lookup_else_if_a0_frac_3_sva_mx0w0 = nl_inp_lookup_else_if_a0_frac_3_sva_mx0w0[34:0];
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_2_nl
      = ~((chn_inp_in_rsci_d_mxwt[378]) | IsZero_5U_10U_3_land_3_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_mux_12_nl = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_2_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_3_sva[4]), IsDenorm_5U_10U_3_land_3_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_3_0_mx0w0 = (FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_mux_12_nl)
      | IsInf_5U_10U_3_land_3_lpi_1_dfm | IsNaN_5U_10U_3_land_3_lpi_1_dfm;
  assign IsZero_5U_10U_3_aelse_not_25_nl = ~ IsZero_5U_10U_3_land_3_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_and_8_nl
      = MUX_v_4_2_2(4'b0000, (chn_inp_in_rsci_d_mxwt[377:374]), (IsZero_5U_10U_3_aelse_not_25_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_mux1h_2_nl
      = MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_and_8_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_3_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_2_cse
      , IsDenorm_5U_10U_3_land_3_lpi_1_dfm , IsInf_5U_10U_3_land_3_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_3_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_mux1h_2_nl),
      4'b1111, IsNaN_5U_10U_3_land_3_lpi_1_dfm);
  assign inp_lookup_3_FpMantRNE_36U_11U_1_else_and_tmp = FpMantRNE_36U_11U_1_else_carry_3_sva
      & (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[35:25]==11'b11111111111);
  assign nl_inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_nl =
      conv_u2u_5_6(libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_14[5:1])
      + 6'b110001;
  assign inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_nl = nl_inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_nl[5:0];
  assign inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_itm_5 =
      readslicef_6_1_5((inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_nl));
  assign inp_lookup_else_if_unequal_tmp_3_mx0w1 = (chn_inp_in_rsci_d_mxwt[267:233]!=35'b00000000000000000000000000000000000);
  assign nl_inp_lookup_else_if_a0_frac_sva_mx0w0 = (~ (chn_inp_in_rsci_d_mxwt[267:233]))
      + 35'b1;
  assign inp_lookup_else_if_a0_frac_sva_mx0w0 = nl_inp_lookup_else_if_a0_frac_sva_mx0w0[34:0];
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_3_nl
      = ~((chn_inp_in_rsci_d_mxwt[394]) | IsZero_5U_10U_3_land_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_mux_17_nl = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_3_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_sva[4]), IsDenorm_5U_10U_3_land_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_3_0_mx0w0 = (FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_mux_17_nl)
      | IsInf_5U_10U_3_land_lpi_1_dfm | IsNaN_5U_10U_3_land_lpi_1_dfm;
  assign IsZero_5U_10U_3_aelse_not_24_nl = ~ IsZero_5U_10U_3_land_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_and_11_nl
      = MUX_v_4_2_2(4'b0000, (chn_inp_in_rsci_d_mxwt[393:390]), (IsZero_5U_10U_3_aelse_not_24_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_mux1h_3_nl
      = MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_and_11_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_3_cse
      , IsDenorm_5U_10U_3_land_lpi_1_dfm , IsInf_5U_10U_3_land_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_mux1h_3_nl),
      4'b1111, IsNaN_5U_10U_3_land_lpi_1_dfm);
  assign inp_lookup_4_FpMantRNE_36U_11U_1_else_and_tmp = FpMantRNE_36U_11U_1_else_carry_sva
      & (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[35:25]==11'b11111111111);
  assign nl_inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_nl =
      conv_u2u_5_6(libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_15[5:1])
      + 6'b110001;
  assign inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_nl = nl_inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_nl[5:0];
  assign inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_itm_5 =
      readslicef_6_1_5((inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_nl));
  assign FpFractionToFloat_35U_6U_10U_is_zero_1_lpi_1_dfm_mx0w0 = ~(inp_lookup_1_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_itm_5_1
      | inp_lookup_1_FpMantRNE_36U_11U_else_and_tmp);
  assign mux_75_nl = MUX_s_1_2_2(FpAdd_8U_23U_else_6_mux_mx0w1, (chn_inp_in_crt_sva_1_739_395_1[116]),
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_3);
  assign inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_mx0w1
      = (chn_inp_in_crt_sva_1_127_0_1[31]) ^ (mux_75_nl);
  assign FpFractionToFloat_35U_6U_10U_1_o_mant_1_lpi_1_dfm_3_mx0w0 = FpFractionToFloat_35U_6U_10U_1_o_mant_1_lpi_1_dfm_6
      & ({{9{FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_st_2}}, FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_st_2})
      & (signext_10_1(~ FpFractionToFloat_35U_6U_10U_1_is_zero_1_lpi_1_dfm_1));
  assign nl_inp_lookup_1_FpMul_6U_10U_2_else_2_acc_1_nl = conv_u2u_6_7({FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_3_5_mx0w0
      , FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_3_4_0_mx0w0}) + conv_u2u_6_7({FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_6_1_1
      , FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_6_0_1 , FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_9});
  assign inp_lookup_1_FpMul_6U_10U_2_else_2_acc_1_nl = nl_inp_lookup_1_FpMul_6U_10U_2_else_2_acc_1_nl[6:0];
  assign nl_inp_lookup_1_FpMul_6U_10U_2_else_2_if_acc_nl = conv_u2u_6_7(readslicef_7_6_1((inp_lookup_1_FpMul_6U_10U_2_else_2_acc_1_nl)))
      + 7'b1010001;
  assign inp_lookup_1_FpMul_6U_10U_2_else_2_if_acc_nl = nl_inp_lookup_1_FpMul_6U_10U_2_else_2_if_acc_nl[6:0];
  assign inp_lookup_1_FpMul_6U_10U_2_else_2_if_acc_itm_6 = readslicef_7_1_6((inp_lookup_1_FpMul_6U_10U_2_else_2_if_acc_nl));
  assign nl_FpMul_6U_10U_2_oelse_1_acc_nl = conv_u2s_6_7({FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_6_1_1
      , FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_6_0_1 , FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_9})
      + 7'b1100001;
  assign FpMul_6U_10U_2_oelse_1_acc_nl = nl_FpMul_6U_10U_2_oelse_1_acc_nl[6:0];
  assign nl_inp_lookup_1_FpMul_6U_10U_2_oelse_1_acc_nl = conv_s2s_7_8(FpMul_6U_10U_2_oelse_1_acc_nl)
      + conv_u2s_6_8({FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_3_5_mx0w0
      , FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_3_4_0_mx0w0});
  assign inp_lookup_1_FpMul_6U_10U_2_oelse_1_acc_nl = nl_inp_lookup_1_FpMul_6U_10U_2_oelse_1_acc_nl[7:0];
  assign inp_lookup_1_FpMul_6U_10U_2_oelse_1_acc_itm_7 = readslicef_8_1_7((inp_lookup_1_FpMul_6U_10U_2_oelse_1_acc_nl));
  assign IsZero_6U_10U_6_IsZero_6U_10U_6_nor_tmp = ~((FpFractionToFloat_35U_6U_10U_1_o_mant_1_lpi_1_dfm_3_mx0w0!=10'b0000000000)
      | FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_3_5_mx0w0 | (FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_3_4_0_mx0w0!=5'b00000));
  assign FpFractionToFloat_35U_6U_10U_is_zero_2_lpi_1_dfm_mx0w0 = ~(inp_lookup_2_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_itm_5_1
      | inp_lookup_2_FpMantRNE_36U_11U_else_and_tmp);
  assign mux_76_nl = MUX_s_1_2_2(FpAdd_8U_23U_else_6_mux_3_mx0w1, (chn_inp_in_crt_sva_1_739_395_1[148]),
      IsNaN_8U_23U_land_2_lpi_1_dfm_4);
  assign inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_mx0w1
      = (chn_inp_in_crt_sva_1_127_0_1[63]) ^ (mux_76_nl);
  assign FpFractionToFloat_35U_6U_10U_1_o_mant_2_lpi_1_dfm_3_mx0w0 = FpFractionToFloat_35U_6U_10U_1_o_mant_2_lpi_1_dfm_6
      & ({{9{FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_st_2}}, FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_st_2})
      & (signext_10_1(~ FpFractionToFloat_35U_6U_10U_1_is_zero_2_lpi_1_dfm_1));
  assign nl_inp_lookup_2_FpMul_6U_10U_2_else_2_acc_1_nl = conv_u2u_6_7({FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_3_5_mx0w0
      , FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_3_4_0_mx0w0}) + conv_u2u_6_7({FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_6_1_1
      , FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_6_0_1 , FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_9});
  assign inp_lookup_2_FpMul_6U_10U_2_else_2_acc_1_nl = nl_inp_lookup_2_FpMul_6U_10U_2_else_2_acc_1_nl[6:0];
  assign nl_inp_lookup_2_FpMul_6U_10U_2_else_2_if_acc_nl = conv_u2u_6_7(readslicef_7_6_1((inp_lookup_2_FpMul_6U_10U_2_else_2_acc_1_nl)))
      + 7'b1010001;
  assign inp_lookup_2_FpMul_6U_10U_2_else_2_if_acc_nl = nl_inp_lookup_2_FpMul_6U_10U_2_else_2_if_acc_nl[6:0];
  assign inp_lookup_2_FpMul_6U_10U_2_else_2_if_acc_itm_6 = readslicef_7_1_6((inp_lookup_2_FpMul_6U_10U_2_else_2_if_acc_nl));
  assign nl_FpMul_6U_10U_2_oelse_1_acc_1_nl = conv_u2s_6_7({FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_6_1_1
      , FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_6_0_1 , FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_9})
      + 7'b1100001;
  assign FpMul_6U_10U_2_oelse_1_acc_1_nl = nl_FpMul_6U_10U_2_oelse_1_acc_1_nl[6:0];
  assign nl_inp_lookup_2_FpMul_6U_10U_2_oelse_1_acc_nl = conv_s2s_7_8(FpMul_6U_10U_2_oelse_1_acc_1_nl)
      + conv_u2s_6_8({FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_3_5_mx0w0
      , FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_3_4_0_mx0w0});
  assign inp_lookup_2_FpMul_6U_10U_2_oelse_1_acc_nl = nl_inp_lookup_2_FpMul_6U_10U_2_oelse_1_acc_nl[7:0];
  assign inp_lookup_2_FpMul_6U_10U_2_oelse_1_acc_itm_7 = readslicef_8_1_7((inp_lookup_2_FpMul_6U_10U_2_oelse_1_acc_nl));
  assign IsZero_6U_10U_6_IsZero_6U_10U_6_nor_1_tmp = ~((FpFractionToFloat_35U_6U_10U_1_o_mant_2_lpi_1_dfm_3_mx0w0!=10'b0000000000)
      | FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_3_5_mx0w0 | (FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_3_4_0_mx0w0!=5'b00000));
  assign FpFractionToFloat_35U_6U_10U_is_zero_3_lpi_1_dfm_mx0w0 = ~(inp_lookup_3_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_itm_5_1
      | inp_lookup_3_FpMantRNE_36U_11U_else_and_tmp);
  assign mux_77_nl = MUX_s_1_2_2(FpAdd_8U_23U_else_6_mux_6_mx0w1, (chn_inp_in_crt_sva_1_739_395_1[180]),
      IsNaN_8U_23U_land_3_lpi_1_dfm_4);
  assign inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_mx0w1
      = (chn_inp_in_crt_sva_1_127_0_1[95]) ^ (mux_77_nl);
  assign FpFractionToFloat_35U_6U_10U_1_o_mant_3_lpi_1_dfm_3_mx0w0 = FpFractionToFloat_35U_6U_10U_1_o_mant_3_lpi_1_dfm_6
      & ({{9{FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_st_2}}, FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_st_2})
      & (signext_10_1(~ FpFractionToFloat_35U_6U_10U_1_is_zero_3_lpi_1_dfm_1));
  assign nl_inp_lookup_3_FpMul_6U_10U_2_else_2_acc_1_nl = conv_u2u_6_7({FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_3_5_mx0w0
      , FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_3_4_0_mx0w0}) + conv_u2u_6_7({FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_6_1_1
      , FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_6_0_1 , FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_3_lpi_1_dfm_9});
  assign inp_lookup_3_FpMul_6U_10U_2_else_2_acc_1_nl = nl_inp_lookup_3_FpMul_6U_10U_2_else_2_acc_1_nl[6:0];
  assign nl_inp_lookup_3_FpMul_6U_10U_2_else_2_if_acc_nl = conv_u2u_6_7(readslicef_7_6_1((inp_lookup_3_FpMul_6U_10U_2_else_2_acc_1_nl)))
      + 7'b1010001;
  assign inp_lookup_3_FpMul_6U_10U_2_else_2_if_acc_nl = nl_inp_lookup_3_FpMul_6U_10U_2_else_2_if_acc_nl[6:0];
  assign inp_lookup_3_FpMul_6U_10U_2_else_2_if_acc_itm_6_1 = readslicef_7_1_6((inp_lookup_3_FpMul_6U_10U_2_else_2_if_acc_nl));
  assign nl_FpMul_6U_10U_2_oelse_1_acc_2_nl = conv_u2s_6_7({FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_6_1_1
      , FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_6_0_1 , FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_3_lpi_1_dfm_9})
      + 7'b1100001;
  assign FpMul_6U_10U_2_oelse_1_acc_2_nl = nl_FpMul_6U_10U_2_oelse_1_acc_2_nl[6:0];
  assign nl_inp_lookup_3_FpMul_6U_10U_2_oelse_1_acc_nl = conv_s2s_7_8(FpMul_6U_10U_2_oelse_1_acc_2_nl)
      + conv_u2s_6_8({FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_3_5_mx0w0
      , FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_3_4_0_mx0w0});
  assign inp_lookup_3_FpMul_6U_10U_2_oelse_1_acc_nl = nl_inp_lookup_3_FpMul_6U_10U_2_oelse_1_acc_nl[7:0];
  assign FpMul_6U_10U_2_if_2_FpMul_6U_10U_2_if_2_or_5_tmp = (readslicef_8_1_7((inp_lookup_3_FpMul_6U_10U_2_oelse_1_acc_nl)))
      | IsZero_6U_10U_7_IsZero_6U_10U_7_and_2_itm_2 | (~((FpFractionToFloat_35U_6U_10U_1_o_mant_3_lpi_1_dfm_3_mx0w0!=10'b0000000000)
      | FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_3_5_mx0w0 | (FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_3_4_0_mx0w0!=5'b00000)));
  assign FpFractionToFloat_35U_6U_10U_is_zero_lpi_1_dfm_mx0w0 = ~(inp_lookup_4_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_itm_5_1
      | inp_lookup_4_FpMantRNE_36U_11U_else_and_tmp);
  assign mux_69_nl = MUX_s_1_2_2(FpAdd_8U_23U_else_6_mux_9_mx0w1, (chn_inp_in_crt_sva_1_739_395_1[212]),
      IsNaN_8U_23U_land_lpi_1_dfm_4);
  assign inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_mx0w1
      = (chn_inp_in_crt_sva_1_127_0_1[127]) ^ (mux_69_nl);
  assign FpFractionToFloat_35U_6U_10U_1_o_mant_lpi_1_dfm_3_mx0w0 = FpFractionToFloat_35U_6U_10U_1_o_mant_lpi_1_dfm_6
      & ({{9{FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2}}, FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2})
      & (signext_10_1(~ FpFractionToFloat_35U_6U_10U_1_is_zero_lpi_1_dfm_1));
  assign nl_inp_lookup_4_FpMul_6U_10U_2_else_2_acc_1_nl = conv_u2u_6_7({FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_3_5_mx0w0
      , FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_3_4_0_mx0w0}) + conv_u2u_6_7({FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_6_1_1
      , FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_6_0_1 , FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_9});
  assign inp_lookup_4_FpMul_6U_10U_2_else_2_acc_1_nl = nl_inp_lookup_4_FpMul_6U_10U_2_else_2_acc_1_nl[6:0];
  assign nl_inp_lookup_4_FpMul_6U_10U_2_else_2_if_acc_nl = conv_u2u_6_7(readslicef_7_6_1((inp_lookup_4_FpMul_6U_10U_2_else_2_acc_1_nl)))
      + 7'b1010001;
  assign inp_lookup_4_FpMul_6U_10U_2_else_2_if_acc_nl = nl_inp_lookup_4_FpMul_6U_10U_2_else_2_if_acc_nl[6:0];
  assign inp_lookup_4_FpMul_6U_10U_2_else_2_if_acc_itm_6 = readslicef_7_1_6((inp_lookup_4_FpMul_6U_10U_2_else_2_if_acc_nl));
  assign nl_FpMul_6U_10U_2_oelse_1_acc_3_nl = conv_u2s_6_7({FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_6_1_1
      , FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_6_0_1 , FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_9})
      + 7'b1100001;
  assign FpMul_6U_10U_2_oelse_1_acc_3_nl = nl_FpMul_6U_10U_2_oelse_1_acc_3_nl[6:0];
  assign nl_inp_lookup_4_FpMul_6U_10U_2_oelse_1_acc_nl = conv_s2s_7_8(FpMul_6U_10U_2_oelse_1_acc_3_nl)
      + conv_u2s_6_8({FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_3_5_mx0w0 ,
      FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_3_4_0_mx0w0});
  assign inp_lookup_4_FpMul_6U_10U_2_oelse_1_acc_nl = nl_inp_lookup_4_FpMul_6U_10U_2_oelse_1_acc_nl[7:0];
  assign inp_lookup_4_FpMul_6U_10U_2_oelse_1_acc_itm_7 = readslicef_8_1_7((inp_lookup_4_FpMul_6U_10U_2_oelse_1_acc_nl));
  assign IsZero_6U_10U_6_IsZero_6U_10U_6_nor_3_tmp = ~((FpFractionToFloat_35U_6U_10U_1_o_mant_lpi_1_dfm_3_mx0w0!=10'b0000000000)
      | FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_3_5_mx0w0 | (FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_3_4_0_mx0w0!=5'b00000));
  assign FpMul_6U_10U_2_if_2_FpMul_6U_10U_2_if_2_or_7_tmp = inp_lookup_4_FpMul_6U_10U_2_oelse_1_acc_itm_7
      | IsZero_6U_10U_7_IsZero_6U_10U_7_and_3_itm_2 | IsZero_6U_10U_6_IsZero_6U_10U_6_nor_3_tmp;
  assign nl_inp_lookup_1_FpAdd_8U_23U_if_3_if_acc_1_nl = ({1'b1 , (reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_7_1_itm[7:1])})
      + 8'b1;
  assign inp_lookup_1_FpAdd_8U_23U_if_3_if_acc_1_nl = nl_inp_lookup_1_FpAdd_8U_23U_if_3_if_acc_1_nl[7:0];
  assign inp_lookup_1_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1 = readslicef_8_1_7((inp_lookup_1_FpAdd_8U_23U_if_3_if_acc_1_nl));
  assign inp_lookup_1_FpMantRNE_22U_11U_2_else_and_tmp = FpMantRNE_22U_11U_2_else_carry_1_sva_mx1w1
      & (FpMul_6U_10U_2_p_mant_20_1_1_lpi_1_dfm_3_mx0[19:10]==10'b1111111111);
  assign FpAdd_8U_23U_or_cse = FpMul_6U_10U_2_and_ssc | IsNaN_6U_10U_6_land_1_lpi_1_dfm_5;
  assign nl_inp_lookup_1_FpAdd_8U_23U_if_4_if_acc_nl = FpAdd_8U_23U_o_expo_1_lpi_1_dfm_10
      + 8'b1;
  assign inp_lookup_1_FpAdd_8U_23U_if_4_if_acc_nl = nl_inp_lookup_1_FpAdd_8U_23U_if_4_if_acc_nl[7:0];
  assign FpAdd_8U_23U_and_nl = (~(FpAdd_8U_23U_and_tmp | FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0))
      & FpMul_6U_10U_2_FpMul_6U_10U_2_nor_ssc;
  assign FpAdd_8U_23U_and_6_nl = FpAdd_8U_23U_and_tmp & (~ FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0)
      & FpMul_6U_10U_2_FpMul_6U_10U_2_nor_ssc;
  assign FpAdd_8U_23U_and_28_nl = FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0 & FpMul_6U_10U_2_FpMul_6U_10U_2_nor_ssc;
  assign FpAdd_8U_23U_o_expo_1_lpi_1_dfm_7_mx1w1 = MUX1HOT_v_8_4_2(FpAdd_8U_23U_o_expo_1_lpi_1_dfm_10,
      (inp_lookup_1_FpAdd_8U_23U_if_4_if_acc_nl), 8'b11111110, reg_chn_inp_in_crt_sva_3_510_480_reg,
      {(FpAdd_8U_23U_and_nl) , (FpAdd_8U_23U_and_6_nl) , (FpAdd_8U_23U_and_28_nl)
      , FpAdd_8U_23U_or_cse});
  assign inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_3_5_mx0w1 = inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_5_1
      & IsNaN_8U_23U_land_1_lpi_1_dfm_st_4;
  assign inp_lookup_else_if_a0_9_0_1_lpi_1_dfm_3_mx0w0 = FpFractionToFloat_35U_6U_10U_if_else_mux_2_itm_2
      & (signext_10_1(~ FpFractionToFloat_35U_6U_10U_is_zero_1_lpi_1_dfm_5)) & ({{9{IsNaN_8U_23U_land_1_lpi_1_dfm_st_4}},
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_4});
  assign nl_inp_lookup_1_FpMul_6U_10U_1_else_2_acc_1_nl = conv_u2u_6_7({inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_3_5_mx0w1
      , inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_3_4_0_mx0w0}) + conv_u2u_6_7({FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_7_1_1
      , FpAdd_8U_23U_o_sign_1_lpi_1_dfm_7 , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_9});
  assign inp_lookup_1_FpMul_6U_10U_1_else_2_acc_1_nl = nl_inp_lookup_1_FpMul_6U_10U_1_else_2_acc_1_nl[6:0];
  assign nl_inp_lookup_1_FpMul_6U_10U_1_else_2_if_acc_nl = conv_u2u_6_7(readslicef_7_6_1((inp_lookup_1_FpMul_6U_10U_1_else_2_acc_1_nl)))
      + 7'b1010001;
  assign inp_lookup_1_FpMul_6U_10U_1_else_2_if_acc_nl = nl_inp_lookup_1_FpMul_6U_10U_1_else_2_if_acc_nl[6:0];
  assign inp_lookup_1_FpMul_6U_10U_1_else_2_if_acc_itm_6_1 = readslicef_7_1_6((inp_lookup_1_FpMul_6U_10U_1_else_2_if_acc_nl));
  assign nl_inp_lookup_1_FpMul_6U_10U_2_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_6U_10U_2_else_2_else_ac_int_cctor_1_sva_mx0w0[5:1])})
      + 6'b1;
  assign inp_lookup_1_FpMul_6U_10U_2_else_2_else_if_if_acc_1_nl = nl_inp_lookup_1_FpMul_6U_10U_2_else_2_else_if_if_acc_1_nl[5:0];
  assign inp_lookup_1_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1 = readslicef_6_1_5((inp_lookup_1_FpMul_6U_10U_2_else_2_else_if_if_acc_1_nl));
  assign FpMul_6U_10U_2_FpMul_6U_10U_2_and_20_nl = (FpMul_6U_10U_2_o_expo_1_lpi_1_dfm[5])
      & (~ FpMul_6U_10U_2_lor_9_lpi_1_dfm);
  assign FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_3_5_mx1w1 = MUX1HOT_s_1_3_2(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_2,
      FpMantRNE_22U_11U_1_else_carry_1_sva_1, (FpMul_6U_10U_2_FpMul_6U_10U_2_and_20_nl),
      {IsNaN_6U_10U_6_land_1_lpi_1_dfm_5 , FpMul_6U_10U_2_and_ssc , FpMul_6U_10U_2_FpMul_6U_10U_2_nor_ssc});
  assign nl_inp_lookup_2_FpAdd_8U_23U_if_3_if_acc_1_nl = ({1'b1 , (reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_7_1_itm[7:1])})
      + 8'b1;
  assign inp_lookup_2_FpAdd_8U_23U_if_3_if_acc_1_nl = nl_inp_lookup_2_FpAdd_8U_23U_if_3_if_acc_1_nl[7:0];
  assign inp_lookup_2_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1 = readslicef_8_1_7((inp_lookup_2_FpAdd_8U_23U_if_3_if_acc_1_nl));
  assign inp_lookup_2_FpMantRNE_22U_11U_2_else_and_tmp = FpMantRNE_22U_11U_2_else_carry_2_sva_mx1w1
      & (FpMul_6U_10U_2_p_mant_20_1_2_lpi_1_dfm_3_mx0[19:10]==10'b1111111111);
  assign FpAdd_8U_23U_or_1_cse = FpMul_6U_10U_2_and_2_ssc | IsNaN_6U_10U_6_land_2_lpi_1_dfm_5;
  assign nl_inp_lookup_2_FpAdd_8U_23U_if_4_if_acc_nl = FpAdd_8U_23U_o_expo_2_lpi_1_dfm_10
      + 8'b1;
  assign inp_lookup_2_FpAdd_8U_23U_if_4_if_acc_nl = nl_inp_lookup_2_FpAdd_8U_23U_if_4_if_acc_nl[7:0];
  assign FpAdd_8U_23U_and_29_nl = (~(FpAdd_8U_23U_and_1_tmp | FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0))
      & FpMul_6U_10U_2_FpMul_6U_10U_2_nor_1_ssc;
  assign FpAdd_8U_23U_and_13_nl = FpAdd_8U_23U_and_1_tmp & (~ FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0)
      & FpMul_6U_10U_2_FpMul_6U_10U_2_nor_1_ssc;
  assign FpAdd_8U_23U_and_30_nl = FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0 & FpMul_6U_10U_2_FpMul_6U_10U_2_nor_1_ssc;
  assign FpAdd_8U_23U_o_expo_2_lpi_1_dfm_7_mx1w1 = MUX1HOT_v_8_4_2(FpAdd_8U_23U_o_expo_2_lpi_1_dfm_10,
      (inp_lookup_2_FpAdd_8U_23U_if_4_if_acc_nl), 8'b11111110, reg_chn_inp_in_crt_sva_3_542_512_reg,
      {(FpAdd_8U_23U_and_29_nl) , (FpAdd_8U_23U_and_13_nl) , (FpAdd_8U_23U_and_30_nl)
      , FpAdd_8U_23U_or_1_cse});
  assign inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_3_5_mx0w1 = inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_6_5_1
      & IsNaN_8U_23U_land_2_lpi_1_dfm_st_4;
  assign inp_lookup_else_if_a0_9_0_2_lpi_1_dfm_3_mx0w0 = FpFractionToFloat_35U_6U_10U_if_else_mux_6_itm_2
      & (signext_10_1(~ FpFractionToFloat_35U_6U_10U_is_zero_2_lpi_1_dfm_5)) & ({{9{IsNaN_8U_23U_land_2_lpi_1_dfm_st_4}},
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_4});
  assign nl_inp_lookup_2_FpMul_6U_10U_1_else_2_acc_1_nl = conv_u2u_6_7({inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_3_5_mx0w1
      , inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_3_4_0_mx0w0}) + conv_u2u_6_7({FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_7_1_1
      , FpAdd_8U_23U_o_sign_2_lpi_1_dfm_7 , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_9});
  assign inp_lookup_2_FpMul_6U_10U_1_else_2_acc_1_nl = nl_inp_lookup_2_FpMul_6U_10U_1_else_2_acc_1_nl[6:0];
  assign nl_inp_lookup_2_FpMul_6U_10U_1_else_2_if_acc_nl = conv_u2u_6_7(readslicef_7_6_1((inp_lookup_2_FpMul_6U_10U_1_else_2_acc_1_nl)))
      + 7'b1010001;
  assign inp_lookup_2_FpMul_6U_10U_1_else_2_if_acc_nl = nl_inp_lookup_2_FpMul_6U_10U_1_else_2_if_acc_nl[6:0];
  assign inp_lookup_2_FpMul_6U_10U_1_else_2_if_acc_itm_6_1 = readslicef_7_1_6((inp_lookup_2_FpMul_6U_10U_1_else_2_if_acc_nl));
  assign nl_inp_lookup_2_FpMul_6U_10U_2_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_6U_10U_2_else_2_else_ac_int_cctor_2_sva_mx0w0[5:1])})
      + 6'b1;
  assign inp_lookup_2_FpMul_6U_10U_2_else_2_else_if_if_acc_1_nl = nl_inp_lookup_2_FpMul_6U_10U_2_else_2_else_if_if_acc_1_nl[5:0];
  assign inp_lookup_2_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1 = readslicef_6_1_5((inp_lookup_2_FpMul_6U_10U_2_else_2_else_if_if_acc_1_nl));
  assign FpMul_6U_10U_2_FpMul_6U_10U_2_and_22_nl = (FpMul_6U_10U_2_o_expo_2_lpi_1_dfm[5])
      & (~ FpMul_6U_10U_2_lor_10_lpi_1_dfm);
  assign FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_3_5_mx1w1 = MUX1HOT_s_1_3_2(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_2,
      FpMantRNE_22U_11U_1_else_carry_2_sva_1, (FpMul_6U_10U_2_FpMul_6U_10U_2_and_22_nl),
      {IsNaN_6U_10U_6_land_2_lpi_1_dfm_5 , FpMul_6U_10U_2_and_2_ssc , FpMul_6U_10U_2_FpMul_6U_10U_2_nor_1_ssc});
  assign nl_inp_lookup_3_FpAdd_8U_23U_if_3_if_acc_1_nl = ({1'b1 , (reg_FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_7_1_itm[7:1])})
      + 8'b1;
  assign inp_lookup_3_FpAdd_8U_23U_if_3_if_acc_1_nl = nl_inp_lookup_3_FpAdd_8U_23U_if_3_if_acc_1_nl[7:0];
  assign inp_lookup_3_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1 = readslicef_8_1_7((inp_lookup_3_FpAdd_8U_23U_if_3_if_acc_1_nl));
  assign inp_lookup_3_FpMantRNE_22U_11U_2_else_and_tmp = FpMantRNE_22U_11U_2_else_carry_3_sva_mx1w1
      & (FpMul_6U_10U_2_p_mant_20_1_3_lpi_1_dfm_3_mx0[19:10]==10'b1111111111);
  assign FpAdd_8U_23U_or_2_cse = FpMul_6U_10U_2_and_4_ssc | IsNaN_6U_10U_6_land_3_lpi_1_dfm_5;
  assign nl_inp_lookup_3_FpAdd_8U_23U_if_4_if_acc_nl = FpAdd_8U_23U_o_expo_3_lpi_1_dfm_10
      + 8'b1;
  assign inp_lookup_3_FpAdd_8U_23U_if_4_if_acc_nl = nl_inp_lookup_3_FpAdd_8U_23U_if_4_if_acc_nl[7:0];
  assign FpAdd_8U_23U_and_31_nl = (~(FpAdd_8U_23U_and_2_tmp | FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0))
      & FpMul_6U_10U_2_FpMul_6U_10U_2_nor_2_ssc;
  assign FpAdd_8U_23U_and_19_nl = FpAdd_8U_23U_and_2_tmp & (~ FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0)
      & FpMul_6U_10U_2_FpMul_6U_10U_2_nor_2_ssc;
  assign FpAdd_8U_23U_and_32_nl = FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0 & FpMul_6U_10U_2_FpMul_6U_10U_2_nor_2_ssc;
  assign FpAdd_8U_23U_o_expo_3_lpi_1_dfm_7_mx1w1 = MUX1HOT_v_8_4_2(FpAdd_8U_23U_o_expo_3_lpi_1_dfm_10,
      (inp_lookup_3_FpAdd_8U_23U_if_4_if_acc_nl), 8'b11111110, reg_chn_inp_in_crt_sva_3_574_544_reg,
      {(FpAdd_8U_23U_and_31_nl) , (FpAdd_8U_23U_and_19_nl) , (FpAdd_8U_23U_and_32_nl)
      , FpAdd_8U_23U_or_2_cse});
  assign inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_3_5_mx0w1 = inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_6_5_1
      & IsNaN_8U_23U_land_3_lpi_1_dfm_st_4;
  assign inp_lookup_else_if_a0_9_0_3_lpi_1_dfm_3_mx0w0 = FpFractionToFloat_35U_6U_10U_if_else_mux_10_itm_2
      & (signext_10_1(~ FpFractionToFloat_35U_6U_10U_is_zero_3_lpi_1_dfm_5)) & ({{9{IsNaN_8U_23U_land_3_lpi_1_dfm_st_4}},
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_4});
  assign nl_inp_lookup_3_FpMantRNE_22U_11U_2_else_acc_nl = FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_3_lpi_1_dfm_10
      + conv_u2u_1_10(FpMantRNE_22U_11U_1_else_carry_3_sva_1);
  assign inp_lookup_3_FpMantRNE_22U_11U_2_else_acc_nl = nl_inp_lookup_3_FpMantRNE_22U_11U_2_else_acc_nl[9:0];
  assign or_5848_nl = FpMantWidthDec_6U_21U_10U_0U_0U_2_if_1_unequal_tmp_2 | (~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_2);
  assign mux_2023_nl = MUX_v_10_2_2((signext_10_1(~ FpMantWidthDec_6U_21U_10U_0U_0U_2_if_1_unequal_tmp_2)),
      (inp_lookup_3_FpMantRNE_22U_11U_2_else_acc_nl), or_5848_nl);
  assign FpMul_6U_10U_2_nor_5_nl = ~(MUX_v_10_2_2((mux_2023_nl), 10'b1111111111,
      nor_1789_cse));
  assign FpMul_6U_10U_2_FpMul_6U_10U_2_FpMul_6U_10U_2_nor_6_nl = ~(MUX_v_10_2_2((FpMul_6U_10U_2_nor_5_nl),
      10'b1111111111, FpMul_6U_10U_2_lor_11_lpi_1_dfm));
  assign FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_3_mx1w1 = MUX_v_10_2_2((FpMul_6U_10U_2_FpMul_6U_10U_2_FpMul_6U_10U_2_nor_6_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_3_lpi_1_dfm_10, FpAdd_8U_23U_or_2_cse);
  assign nl_inp_lookup_3_FpMul_6U_10U_1_else_2_acc_1_nl = conv_u2u_6_7({inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_3_5_mx0w1
      , inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_3_4_0_mx0w0}) + conv_u2u_6_7({FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_7_1_1
      , FpAdd_8U_23U_o_sign_3_lpi_1_dfm_7 , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_9});
  assign inp_lookup_3_FpMul_6U_10U_1_else_2_acc_1_nl = nl_inp_lookup_3_FpMul_6U_10U_1_else_2_acc_1_nl[6:0];
  assign nl_inp_lookup_3_FpMul_6U_10U_1_else_2_if_acc_nl = conv_u2u_6_7(readslicef_7_6_1((inp_lookup_3_FpMul_6U_10U_1_else_2_acc_1_nl)))
      + 7'b1010001;
  assign inp_lookup_3_FpMul_6U_10U_1_else_2_if_acc_nl = nl_inp_lookup_3_FpMul_6U_10U_1_else_2_if_acc_nl[6:0];
  assign inp_lookup_3_FpMul_6U_10U_1_else_2_if_acc_itm_6_1 = readslicef_7_1_6((inp_lookup_3_FpMul_6U_10U_1_else_2_if_acc_nl));
  assign nl_inp_lookup_3_FpMul_6U_10U_2_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_6U_10U_2_else_2_else_ac_int_cctor_3_sva_mx0w0[5:1])})
      + 6'b1;
  assign inp_lookup_3_FpMul_6U_10U_2_else_2_else_if_if_acc_1_nl = nl_inp_lookup_3_FpMul_6U_10U_2_else_2_else_if_if_acc_1_nl[5:0];
  assign inp_lookup_3_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1 = readslicef_6_1_5((inp_lookup_3_FpMul_6U_10U_2_else_2_else_if_if_acc_1_nl));
  assign FpMul_6U_10U_2_FpMul_6U_10U_2_and_24_nl = (FpMul_6U_10U_2_o_expo_3_lpi_1_dfm[5])
      & (~ FpMul_6U_10U_2_lor_11_lpi_1_dfm);
  assign FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_3_5_mx1w1 = MUX1HOT_s_1_3_2(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_2,
      FpMantRNE_22U_11U_1_else_carry_3_sva_1, (FpMul_6U_10U_2_FpMul_6U_10U_2_and_24_nl),
      {IsNaN_6U_10U_6_land_3_lpi_1_dfm_5 , FpMul_6U_10U_2_and_4_ssc , FpMul_6U_10U_2_FpMul_6U_10U_2_nor_2_ssc});
  assign nl_inp_lookup_4_FpAdd_8U_23U_if_3_if_acc_1_nl = ({1'b1 , (reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_7_1_itm[7:1])})
      + 8'b1;
  assign inp_lookup_4_FpAdd_8U_23U_if_3_if_acc_1_nl = nl_inp_lookup_4_FpAdd_8U_23U_if_3_if_acc_1_nl[7:0];
  assign inp_lookup_4_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1 = readslicef_8_1_7((inp_lookup_4_FpAdd_8U_23U_if_3_if_acc_1_nl));
  assign inp_lookup_4_FpMantRNE_22U_11U_2_else_and_tmp = FpMantRNE_22U_11U_2_else_carry_sva_mx0w2
      & (FpMul_6U_10U_2_p_mant_20_1_lpi_1_dfm_3_mx0[19:10]==10'b1111111111);
  assign FpAdd_8U_23U_or_3_cse = FpMul_6U_10U_2_and_6_ssc | IsNaN_6U_10U_6_land_lpi_1_dfm_5;
  assign nl_inp_lookup_4_FpAdd_8U_23U_if_4_if_acc_nl = FpAdd_8U_23U_o_expo_lpi_1_dfm_10
      + 8'b1;
  assign inp_lookup_4_FpAdd_8U_23U_if_4_if_acc_nl = nl_inp_lookup_4_FpAdd_8U_23U_if_4_if_acc_nl[7:0];
  assign FpAdd_8U_23U_and_33_nl = (~(FpAdd_8U_23U_and_3_tmp | FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0))
      & FpMul_6U_10U_2_FpMul_6U_10U_2_nor_3_ssc;
  assign FpAdd_8U_23U_and_25_nl = FpAdd_8U_23U_and_3_tmp & (~ FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0)
      & FpMul_6U_10U_2_FpMul_6U_10U_2_nor_3_ssc;
  assign FpAdd_8U_23U_and_34_nl = FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0 & FpMul_6U_10U_2_FpMul_6U_10U_2_nor_3_ssc;
  assign FpAdd_8U_23U_o_expo_lpi_1_dfm_7_mx1w1 = MUX1HOT_v_8_4_2(FpAdd_8U_23U_o_expo_lpi_1_dfm_10,
      (inp_lookup_4_FpAdd_8U_23U_if_4_if_acc_nl), 8'b11111110, reg_chn_inp_in_crt_sva_3_606_576_reg,
      {(FpAdd_8U_23U_and_33_nl) , (FpAdd_8U_23U_and_25_nl) , (FpAdd_8U_23U_and_34_nl)
      , FpAdd_8U_23U_or_3_cse});
  assign inp_lookup_else_if_a0_15_10_lpi_1_dfm_3_5_mx0w1 = inp_lookup_else_if_a0_15_10_lpi_1_dfm_6_5_1
      & IsNaN_8U_23U_land_lpi_1_dfm_st_4;
  assign inp_lookup_else_if_a0_9_0_lpi_1_dfm_3_mx0w0 = FpFractionToFloat_35U_6U_10U_if_else_mux_14_itm_2
      & (signext_10_1(~ FpFractionToFloat_35U_6U_10U_is_zero_lpi_1_dfm_5)) & ({{9{IsNaN_8U_23U_land_lpi_1_dfm_st_4}},
      IsNaN_8U_23U_land_lpi_1_dfm_st_4});
  assign nl_inp_lookup_4_FpMul_6U_10U_1_else_2_acc_1_nl = conv_u2u_6_7({inp_lookup_else_if_a0_15_10_lpi_1_dfm_3_5_mx0w1
      , inp_lookup_else_if_a0_15_10_lpi_1_dfm_3_4_0_mx0w0}) + conv_u2u_6_7({FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_7_1_1
      , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_7_0_1 , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_9});
  assign inp_lookup_4_FpMul_6U_10U_1_else_2_acc_1_nl = nl_inp_lookup_4_FpMul_6U_10U_1_else_2_acc_1_nl[6:0];
  assign nl_inp_lookup_4_FpMul_6U_10U_1_else_2_if_acc_nl = conv_u2u_6_7(readslicef_7_6_1((inp_lookup_4_FpMul_6U_10U_1_else_2_acc_1_nl)))
      + 7'b1010001;
  assign inp_lookup_4_FpMul_6U_10U_1_else_2_if_acc_nl = nl_inp_lookup_4_FpMul_6U_10U_1_else_2_if_acc_nl[6:0];
  assign inp_lookup_4_FpMul_6U_10U_1_else_2_if_acc_itm_6_1 = readslicef_7_1_6((inp_lookup_4_FpMul_6U_10U_1_else_2_if_acc_nl));
  assign nl_inp_lookup_4_FpMul_6U_10U_2_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_6U_10U_2_else_2_else_ac_int_cctor_sva_mx0w0[5:1])})
      + 6'b1;
  assign inp_lookup_4_FpMul_6U_10U_2_else_2_else_if_if_acc_1_nl = nl_inp_lookup_4_FpMul_6U_10U_2_else_2_else_if_if_acc_1_nl[5:0];
  assign inp_lookup_4_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1 = readslicef_6_1_5((inp_lookup_4_FpMul_6U_10U_2_else_2_else_if_if_acc_1_nl));
  assign FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0 = ((~ FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_itm_23_1)
      & inp_lookup_1_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp) | FpAdd_8U_23U_1_is_a_greater_acc_itm_8_1;
  assign nl_FpMul_6U_10U_1_else_2_else_acc_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_8_1
      , FpAdd_8U_23U_o_sign_1_lpi_1_dfm_5 , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_10})
      + 6'b100001;
  assign FpMul_6U_10U_1_else_2_else_acc_nl = nl_FpMul_6U_10U_1_else_2_else_acc_nl[5:0];
  assign nl_FpMul_6U_10U_1_else_2_else_ac_int_cctor_1_sva_mx0w0 = (FpMul_6U_10U_1_else_2_else_acc_nl)
      + ({inp_lookup_1_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_itm_2
      , inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_7_4_0_1});
  assign FpMul_6U_10U_1_else_2_else_ac_int_cctor_1_sva_mx0w0 = nl_FpMul_6U_10U_1_else_2_else_ac_int_cctor_1_sva_mx0w0[5:0];
  assign nl_inp_lookup_1_FpMul_6U_10U_1_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_6U_10U_1_else_2_else_ac_int_cctor_1_sva_mx0w0[5:1])})
      + 6'b1;
  assign inp_lookup_1_FpMul_6U_10U_1_else_2_else_if_if_acc_1_nl = nl_inp_lookup_1_FpMul_6U_10U_1_else_2_else_if_if_acc_1_nl[5:0];
  assign inp_lookup_1_FpMul_6U_10U_1_else_2_else_if_if_acc_1_itm_5_1 = readslicef_6_1_5((inp_lookup_1_FpMul_6U_10U_1_else_2_else_if_if_acc_1_nl));
  assign FpMul_6U_10U_1_FpMul_6U_10U_1_and_20_nl = (FpMul_6U_10U_1_o_expo_1_lpi_1_dfm[5])
      & (~ FpMul_6U_10U_1_lor_9_lpi_1_dfm);
  assign FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_3_5_mx1w1 = MUX1HOT_s_1_3_2(inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_8_5_1,
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_9_1, (FpMul_6U_10U_1_FpMul_6U_10U_1_and_20_nl),
      {IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_16 , FpMul_6U_10U_1_and_ssc , FpMul_6U_10U_1_FpMul_6U_10U_1_nor_ssc});
  assign FpMul_6U_10U_2_FpMul_6U_10U_2_and_1_nl = (FpMul_6U_10U_2_o_expo_1_lpi_1_dfm[4])
      & (~ FpMul_6U_10U_2_lor_9_lpi_1_dfm);
  assign FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_3_4_mx0w0 = MUX1HOT_s_1_3_2((FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_7_4_0_1[4]),
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_2, (FpMul_6U_10U_2_FpMul_6U_10U_2_and_1_nl),
      {IsNaN_6U_10U_6_land_1_lpi_1_dfm_5 , FpMul_6U_10U_2_and_ssc , FpMul_6U_10U_2_FpMul_6U_10U_2_nor_ssc});
  assign FpMul_6U_10U_2_oelse_2_not_27_nl = ~ FpMul_6U_10U_2_lor_9_lpi_1_dfm;
  assign FpMul_6U_10U_2_FpMul_6U_10U_2_and_19_nl = MUX_v_4_2_2(4'b0000, (FpMul_6U_10U_2_o_expo_1_lpi_1_dfm[3:0]),
      (FpMul_6U_10U_2_oelse_2_not_27_nl));
  assign FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_3_3_0_mx0w0 = MUX1HOT_v_4_3_2((FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_7_4_0_1[3:0]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_11, (FpMul_6U_10U_2_FpMul_6U_10U_2_and_19_nl),
      {IsNaN_6U_10U_6_land_1_lpi_1_dfm_5 , FpMul_6U_10U_2_and_ssc , FpMul_6U_10U_2_FpMul_6U_10U_2_nor_ssc});
  assign FpMul_6U_10U_1_FpMul_6U_10U_1_and_1_nl = (FpMul_6U_10U_1_o_expo_1_lpi_1_dfm[4])
      & (~ FpMul_6U_10U_1_lor_9_lpi_1_dfm);
  assign FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_3_4_mx1w1 = MUX1HOT_s_1_3_2((inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_8_4_0_1[4]),
      FpAdd_8U_23U_o_sign_1_lpi_1_dfm_8, (FpMul_6U_10U_1_FpMul_6U_10U_1_and_1_nl),
      {IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_16 , FpMul_6U_10U_1_and_ssc , FpMul_6U_10U_1_FpMul_6U_10U_1_nor_ssc});
  assign inp_lookup_1_FpMantRNE_22U_11U_1_else_and_tmp = FpMantRNE_22U_11U_1_else_carry_1_sva
      & (FpMul_6U_10U_1_p_mant_20_1_1_lpi_1_dfm_3_mx0[19:10]==10'b1111111111);
  assign FpMul_6U_10U_1_oelse_2_not_27_nl = ~ FpMul_6U_10U_1_lor_9_lpi_1_dfm;
  assign FpMul_6U_10U_1_FpMul_6U_10U_1_and_19_nl = MUX_v_4_2_2(4'b0000, (FpMul_6U_10U_1_o_expo_1_lpi_1_dfm[3:0]),
      (FpMul_6U_10U_1_oelse_2_not_27_nl));
  assign FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_3_3_0_mx1w1 = MUX1HOT_v_4_3_2((inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_8_4_0_1[3:0]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_11, (FpMul_6U_10U_1_FpMul_6U_10U_1_and_19_nl),
      {IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_16 , FpMul_6U_10U_1_and_ssc , FpMul_6U_10U_1_FpMul_6U_10U_1_nor_ssc});
  assign IsNaN_8U_23U_3_IsNaN_8U_23U_3_nor_tmp = ~((~((FpAdd_8U_23U_o_mant_1_lpi_1_dfm_2_mx2!=23'b00000000000000000000000)))
      | (FpAdd_8U_23U_o_expo_1_lpi_1_dfm_7_mx1w1!=8'b11111111));
  assign FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0 = ((~ FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_1_itm_23_1)
      & inp_lookup_2_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp) | FpAdd_8U_23U_1_is_a_greater_acc_1_itm_8_1;
  assign nl_FpMul_6U_10U_1_else_2_else_acc_2_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_8_1
      , FpAdd_8U_23U_o_sign_2_lpi_1_dfm_5 , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_10})
      + 6'b100001;
  assign FpMul_6U_10U_1_else_2_else_acc_2_nl = nl_FpMul_6U_10U_1_else_2_else_acc_2_nl[5:0];
  assign nl_FpMul_6U_10U_1_else_2_else_ac_int_cctor_2_sva_mx0w0 = (FpMul_6U_10U_1_else_2_else_acc_2_nl)
      + ({inp_lookup_2_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_itm_2
      , inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_7_4_0_1});
  assign FpMul_6U_10U_1_else_2_else_ac_int_cctor_2_sva_mx0w0 = nl_FpMul_6U_10U_1_else_2_else_ac_int_cctor_2_sva_mx0w0[5:0];
  assign nl_inp_lookup_2_FpMul_6U_10U_1_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_6U_10U_1_else_2_else_ac_int_cctor_2_sva_mx0w0[5:1])})
      + 6'b1;
  assign inp_lookup_2_FpMul_6U_10U_1_else_2_else_if_if_acc_1_nl = nl_inp_lookup_2_FpMul_6U_10U_1_else_2_else_if_if_acc_1_nl[5:0];
  assign inp_lookup_2_FpMul_6U_10U_1_else_2_else_if_if_acc_1_itm_5_1 = readslicef_6_1_5((inp_lookup_2_FpMul_6U_10U_1_else_2_else_if_if_acc_1_nl));
  assign FpMul_6U_10U_1_FpMul_6U_10U_1_and_22_nl = (FpMul_6U_10U_1_o_expo_2_lpi_1_dfm[5])
      & (~ FpMul_6U_10U_1_lor_10_lpi_1_dfm);
  assign FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_3_5_mx1w1 = MUX1HOT_s_1_3_2(inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_8_5_1,
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_9_1, (FpMul_6U_10U_1_FpMul_6U_10U_1_and_22_nl),
      {IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_16 , FpMul_6U_10U_1_and_2_ssc , FpMul_6U_10U_1_FpMul_6U_10U_1_nor_1_ssc});
  assign FpMul_6U_10U_2_FpMul_6U_10U_2_and_5_nl = (FpMul_6U_10U_2_o_expo_2_lpi_1_dfm[4])
      & (~ FpMul_6U_10U_2_lor_10_lpi_1_dfm);
  assign FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_3_4_mx0w0 = MUX1HOT_s_1_3_2((FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_7_4_0_1[4]),
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_2, (FpMul_6U_10U_2_FpMul_6U_10U_2_and_5_nl),
      {IsNaN_6U_10U_6_land_2_lpi_1_dfm_5 , FpMul_6U_10U_2_and_2_ssc , FpMul_6U_10U_2_FpMul_6U_10U_2_nor_1_ssc});
  assign FpMul_6U_10U_2_oelse_2_not_26_nl = ~ FpMul_6U_10U_2_lor_10_lpi_1_dfm;
  assign FpMul_6U_10U_2_FpMul_6U_10U_2_and_21_nl = MUX_v_4_2_2(4'b0000, (FpMul_6U_10U_2_o_expo_2_lpi_1_dfm[3:0]),
      (FpMul_6U_10U_2_oelse_2_not_26_nl));
  assign FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_3_3_0_mx0w0 = MUX1HOT_v_4_3_2((FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_7_4_0_1[3:0]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_11, (FpMul_6U_10U_2_FpMul_6U_10U_2_and_21_nl),
      {IsNaN_6U_10U_6_land_2_lpi_1_dfm_5 , FpMul_6U_10U_2_and_2_ssc , FpMul_6U_10U_2_FpMul_6U_10U_2_nor_1_ssc});
  assign FpMul_6U_10U_1_FpMul_6U_10U_1_and_5_nl = (FpMul_6U_10U_1_o_expo_2_lpi_1_dfm[4])
      & (~ FpMul_6U_10U_1_lor_10_lpi_1_dfm);
  assign FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_3_4_mx1w1 = MUX1HOT_s_1_3_2((inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_8_4_0_1[4]),
      FpAdd_8U_23U_o_sign_2_lpi_1_dfm_8, (FpMul_6U_10U_1_FpMul_6U_10U_1_and_5_nl),
      {IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_16 , FpMul_6U_10U_1_and_2_ssc , FpMul_6U_10U_1_FpMul_6U_10U_1_nor_1_ssc});
  assign inp_lookup_2_FpMantRNE_22U_11U_1_else_and_tmp = FpMantRNE_22U_11U_1_else_carry_2_sva
      & (FpMul_6U_10U_1_p_mant_20_1_2_lpi_1_dfm_3_mx0[19:10]==10'b1111111111);
  assign FpMul_6U_10U_1_oelse_2_not_26_nl = ~ FpMul_6U_10U_1_lor_10_lpi_1_dfm;
  assign FpMul_6U_10U_1_FpMul_6U_10U_1_and_21_nl = MUX_v_4_2_2(4'b0000, (FpMul_6U_10U_1_o_expo_2_lpi_1_dfm[3:0]),
      (FpMul_6U_10U_1_oelse_2_not_26_nl));
  assign FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_3_3_0_mx1w1 = MUX1HOT_v_4_3_2((inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_8_4_0_1[3:0]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_11, (FpMul_6U_10U_1_FpMul_6U_10U_1_and_21_nl),
      {IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_16 , FpMul_6U_10U_1_and_2_ssc , FpMul_6U_10U_1_FpMul_6U_10U_1_nor_1_ssc});
  assign IsNaN_8U_23U_3_IsNaN_8U_23U_3_nor_1_tmp = ~((~((FpAdd_8U_23U_o_mant_2_lpi_1_dfm_2_mx2!=23'b00000000000000000000000)))
      | (FpAdd_8U_23U_o_expo_2_lpi_1_dfm_7_mx1w1!=8'b11111111));
  assign FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0 = ((~ FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_2_itm_23_1)
      & inp_lookup_3_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp) | FpAdd_8U_23U_1_is_a_greater_acc_2_itm_8_1;
  assign nl_FpMul_6U_10U_1_else_2_else_acc_3_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_8_1
      , FpAdd_8U_23U_o_sign_3_lpi_1_dfm_8 , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_10})
      + 6'b100001;
  assign FpMul_6U_10U_1_else_2_else_acc_3_nl = nl_FpMul_6U_10U_1_else_2_else_acc_3_nl[5:0];
  assign nl_FpMul_6U_10U_1_else_2_else_ac_int_cctor_3_sva_mx0w0 = (FpMul_6U_10U_1_else_2_else_acc_3_nl)
      + ({inp_lookup_3_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_itm_2
      , inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_7_4_0_1});
  assign FpMul_6U_10U_1_else_2_else_ac_int_cctor_3_sva_mx0w0 = nl_FpMul_6U_10U_1_else_2_else_ac_int_cctor_3_sva_mx0w0[5:0];
  assign nl_inp_lookup_3_FpMul_6U_10U_1_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_6U_10U_1_else_2_else_ac_int_cctor_3_sva_mx0w0[5:1])})
      + 6'b1;
  assign inp_lookup_3_FpMul_6U_10U_1_else_2_else_if_if_acc_1_nl = nl_inp_lookup_3_FpMul_6U_10U_1_else_2_else_if_if_acc_1_nl[5:0];
  assign inp_lookup_3_FpMul_6U_10U_1_else_2_else_if_if_acc_1_itm_5_1 = readslicef_6_1_5((inp_lookup_3_FpMul_6U_10U_1_else_2_else_if_if_acc_1_nl));
  assign FpMul_6U_10U_1_FpMul_6U_10U_1_and_24_nl = (FpMul_6U_10U_1_o_expo_3_lpi_1_dfm[5])
      & (~ FpMul_6U_10U_1_lor_11_lpi_1_dfm);
  assign FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_5_mx1w1 = MUX1HOT_s_1_3_2(inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_8_5_1,
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_9_1, (FpMul_6U_10U_1_FpMul_6U_10U_1_and_24_nl),
      {IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_16 , FpMul_6U_10U_1_and_4_ssc , FpMul_6U_10U_1_FpMul_6U_10U_1_nor_2_ssc});
  assign FpMul_6U_10U_2_FpMul_6U_10U_2_and_9_nl = (FpMul_6U_10U_2_o_expo_3_lpi_1_dfm[4])
      & (~ FpMul_6U_10U_2_lor_11_lpi_1_dfm);
  assign FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_3_4_mx0w0 = MUX1HOT_s_1_3_2((FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_7_4_0_1[4]),
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_2, (FpMul_6U_10U_2_FpMul_6U_10U_2_and_9_nl),
      {IsNaN_6U_10U_6_land_3_lpi_1_dfm_5 , FpMul_6U_10U_2_and_4_ssc , FpMul_6U_10U_2_FpMul_6U_10U_2_nor_2_ssc});
  assign FpMul_6U_10U_2_oelse_2_not_25_nl = ~ FpMul_6U_10U_2_lor_11_lpi_1_dfm;
  assign FpMul_6U_10U_2_FpMul_6U_10U_2_and_23_nl = MUX_v_4_2_2(4'b0000, (FpMul_6U_10U_2_o_expo_3_lpi_1_dfm[3:0]),
      (FpMul_6U_10U_2_oelse_2_not_25_nl));
  assign FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_3_3_0_mx0w0 = MUX1HOT_v_4_3_2((FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_7_4_0_1[3:0]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_3_lpi_1_dfm_11, (FpMul_6U_10U_2_FpMul_6U_10U_2_and_23_nl),
      {IsNaN_6U_10U_6_land_3_lpi_1_dfm_5 , FpMul_6U_10U_2_and_4_ssc , FpMul_6U_10U_2_FpMul_6U_10U_2_nor_2_ssc});
  assign nl_inp_lookup_3_FpMantRNE_22U_11U_1_else_acc_nl = FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_11
      + conv_u2u_1_10(FpAdd_8U_23U_o_sign_3_lpi_1_dfm_9);
  assign inp_lookup_3_FpMantRNE_22U_11U_1_else_acc_nl = nl_inp_lookup_3_FpMantRNE_22U_11U_1_else_acc_nl[9:0];
  assign or_5849_nl = FpMantWidthDec_6U_21U_10U_0U_0U_1_if_1_unequal_tmp_2 | (~ FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_9_1);
  assign mux_2024_nl = MUX_v_10_2_2((signext_10_1(~ FpMantWidthDec_6U_21U_10U_0U_0U_1_if_1_unequal_tmp_2)),
      (inp_lookup_3_FpMantRNE_22U_11U_1_else_acc_nl), or_5849_nl);
  assign FpMul_6U_10U_1_nor_5_nl = ~(MUX_v_10_2_2((mux_2024_nl), 10'b1111111111,
      nor_1191_cse));
  assign FpMul_6U_10U_1_FpMul_6U_10U_1_FpMul_6U_10U_1_nor_6_nl = ~(MUX_v_10_2_2((FpMul_6U_10U_1_nor_5_nl),
      10'b1111111111, FpMul_6U_10U_1_lor_11_lpi_1_dfm));
  assign FpMul_6U_10U_1_or_9_nl = FpMul_6U_10U_1_and_4_ssc | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_16;
  assign FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_3_mx0w1 = MUX_v_10_2_2((FpMul_6U_10U_1_FpMul_6U_10U_1_FpMul_6U_10U_1_nor_6_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_11, FpMul_6U_10U_1_or_9_nl);
  assign FpMul_6U_10U_1_FpMul_6U_10U_1_and_9_nl = (FpMul_6U_10U_1_o_expo_3_lpi_1_dfm[4])
      & (~ FpMul_6U_10U_1_lor_11_lpi_1_dfm);
  assign FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_4_mx1w1 = MUX1HOT_s_1_3_2((inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_8_4_0_1[4]),
      FpAdd_8U_23U_o_sign_3_lpi_1_dfm_9, (FpMul_6U_10U_1_FpMul_6U_10U_1_and_9_nl),
      {IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_16 , FpMul_6U_10U_1_and_4_ssc , FpMul_6U_10U_1_FpMul_6U_10U_1_nor_2_ssc});
  assign inp_lookup_3_FpMantRNE_22U_11U_1_else_and_tmp = FpMantRNE_22U_11U_1_else_carry_3_sva
      & (FpMul_6U_10U_1_p_mant_20_1_3_lpi_1_dfm_3_mx0[19:10]==10'b1111111111);
  assign FpMul_6U_10U_1_oelse_2_not_25_nl = ~ FpMul_6U_10U_1_lor_11_lpi_1_dfm;
  assign FpMul_6U_10U_1_FpMul_6U_10U_1_and_23_nl = MUX_v_4_2_2(4'b0000, (FpMul_6U_10U_1_o_expo_3_lpi_1_dfm[3:0]),
      (FpMul_6U_10U_1_oelse_2_not_25_nl));
  assign FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_3_0_mx1w1 = MUX1HOT_v_4_3_2((inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_8_4_0_1[3:0]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_11, (FpMul_6U_10U_1_FpMul_6U_10U_1_and_23_nl),
      {IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_16 , FpMul_6U_10U_1_and_4_ssc , FpMul_6U_10U_1_FpMul_6U_10U_1_nor_2_ssc});
  assign IsNaN_8U_23U_3_IsNaN_8U_23U_3_nor_2_tmp = ~((~((FpAdd_8U_23U_o_mant_3_lpi_1_dfm_2_mx2!=23'b00000000000000000000000)))
      | (FpAdd_8U_23U_o_expo_3_lpi_1_dfm_7_mx1w1!=8'b11111111));
  assign FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_1_mx0w0 = ((~ FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_3_itm_23_1)
      & inp_lookup_4_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp) | FpAdd_8U_23U_1_is_a_greater_acc_3_itm_8_1;
  assign nl_FpMul_6U_10U_1_else_2_else_acc_4_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_8_1
      , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_8_0 , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_10})
      + 6'b100001;
  assign FpMul_6U_10U_1_else_2_else_acc_4_nl = nl_FpMul_6U_10U_1_else_2_else_acc_4_nl[5:0];
  assign nl_FpMul_6U_10U_1_else_2_else_ac_int_cctor_sva_mx0w0 = (FpMul_6U_10U_1_else_2_else_acc_4_nl)
      + ({inp_lookup_4_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_itm_2
      , inp_lookup_else_if_a0_15_10_lpi_1_dfm_7_4_0_1});
  assign FpMul_6U_10U_1_else_2_else_ac_int_cctor_sva_mx0w0 = nl_FpMul_6U_10U_1_else_2_else_ac_int_cctor_sva_mx0w0[5:0];
  assign nl_inp_lookup_4_FpMul_6U_10U_1_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_6U_10U_1_else_2_else_ac_int_cctor_sva_mx0w0[5:1])})
      + 6'b1;
  assign inp_lookup_4_FpMul_6U_10U_1_else_2_else_if_if_acc_1_nl = nl_inp_lookup_4_FpMul_6U_10U_1_else_2_else_if_if_acc_1_nl[5:0];
  assign inp_lookup_4_FpMul_6U_10U_1_else_2_else_if_if_acc_1_itm_5_1 = readslicef_6_1_5((inp_lookup_4_FpMul_6U_10U_1_else_2_else_if_if_acc_1_nl));
  assign FpMul_6U_10U_1_FpMul_6U_10U_1_and_26_nl = (FpMul_6U_10U_1_o_expo_lpi_1_dfm[5])
      & (~ FpMul_6U_10U_1_lor_2_lpi_1_dfm);
  assign FpMul_6U_10U_1_o_expo_lpi_1_dfm_3_5_mx0w1 = MUX1HOT_s_1_3_2(inp_lookup_else_if_a0_15_10_lpi_1_dfm_8_5_1,
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_9_1, (FpMul_6U_10U_1_FpMul_6U_10U_1_and_26_nl),
      {IsNaN_6U_10U_4_land_lpi_1_dfm_5 , FpMul_6U_10U_1_and_6_ssc , IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0});
  assign FpMul_6U_10U_2_FpMul_6U_10U_2_and_26_nl = (FpMul_6U_10U_2_o_expo_lpi_1_dfm[5])
      & (~ FpMul_6U_10U_2_lor_2_lpi_1_dfm);
  assign FpMul_6U_10U_2_o_expo_lpi_1_dfm_3_5_mx0w0 = MUX1HOT_s_1_3_2(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_sva_2,
      FpMantRNE_22U_11U_1_else_carry_sva, (FpMul_6U_10U_2_FpMul_6U_10U_2_and_26_nl),
      {IsNaN_6U_10U_6_land_lpi_1_dfm_5 , FpMul_6U_10U_2_and_6_ssc , FpMul_6U_10U_2_FpMul_6U_10U_2_nor_3_ssc});
  assign FpMul_6U_10U_2_FpMul_6U_10U_2_and_13_nl = (FpMul_6U_10U_2_o_expo_lpi_1_dfm[4])
      & (~ FpMul_6U_10U_2_lor_2_lpi_1_dfm);
  assign FpMul_6U_10U_2_o_expo_lpi_1_dfm_3_4_mx0w0 = MUX1HOT_s_1_3_2((FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_7_4_0_1[4]),
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_sva_2, (FpMul_6U_10U_2_FpMul_6U_10U_2_and_13_nl),
      {IsNaN_6U_10U_6_land_lpi_1_dfm_5 , FpMul_6U_10U_2_and_6_ssc , FpMul_6U_10U_2_FpMul_6U_10U_2_nor_3_ssc});
  assign FpMul_6U_10U_2_oelse_2_not_24_nl = ~ FpMul_6U_10U_2_lor_2_lpi_1_dfm;
  assign FpMul_6U_10U_2_FpMul_6U_10U_2_and_25_nl = MUX_v_4_2_2(4'b0000, (FpMul_6U_10U_2_o_expo_lpi_1_dfm[3:0]),
      (FpMul_6U_10U_2_oelse_2_not_24_nl));
  assign FpMul_6U_10U_2_o_expo_lpi_1_dfm_3_3_0_mx0w0 = MUX1HOT_v_4_3_2((FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_7_4_0_1[3:0]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_11, (FpMul_6U_10U_2_FpMul_6U_10U_2_and_25_nl),
      {IsNaN_6U_10U_6_land_lpi_1_dfm_5 , FpMul_6U_10U_2_and_6_ssc , FpMul_6U_10U_2_FpMul_6U_10U_2_nor_3_ssc});
  assign IsNaN_8U_23U_3_IsNaN_8U_23U_3_nand_3_tmp = ~((FpAdd_8U_23U_o_expo_lpi_1_dfm_7_mx1w1==8'b11111111));
  assign FpMul_6U_10U_1_FpMul_6U_10U_1_and_13_nl = (FpMul_6U_10U_1_o_expo_lpi_1_dfm[4])
      & (~ FpMul_6U_10U_1_lor_2_lpi_1_dfm);
  assign FpMul_6U_10U_1_o_expo_lpi_1_dfm_3_4_mx0w1 = MUX1HOT_s_1_3_2((inp_lookup_else_if_a0_15_10_lpi_1_dfm_8_4_0_1[4]),
      FpAdd_8U_23U_o_sign_lpi_1_dfm_9, (FpMul_6U_10U_1_FpMul_6U_10U_1_and_13_nl),
      {IsNaN_6U_10U_4_land_lpi_1_dfm_5 , FpMul_6U_10U_1_and_6_ssc , IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0});
  assign inp_lookup_4_FpMantRNE_22U_11U_1_else_and_tmp = FpMantRNE_22U_11U_1_else_carry_sva_mx0w1
      & (FpMul_6U_10U_1_p_mant_20_1_lpi_1_dfm_3_mx0[19:10]==10'b1111111111);
  assign FpMul_6U_10U_1_oelse_2_not_24_nl = ~ FpMul_6U_10U_1_lor_2_lpi_1_dfm;
  assign FpMul_6U_10U_1_FpMul_6U_10U_1_and_25_nl = MUX_v_4_2_2(4'b0000, (FpMul_6U_10U_1_o_expo_lpi_1_dfm[3:0]),
      (FpMul_6U_10U_1_oelse_2_not_24_nl));
  assign FpMul_6U_10U_1_o_expo_lpi_1_dfm_3_3_0_mx0w1 = MUX1HOT_v_4_3_2((inp_lookup_else_if_a0_15_10_lpi_1_dfm_8_4_0_1[3:0]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_11, (FpMul_6U_10U_1_FpMul_6U_10U_1_and_25_nl),
      {IsNaN_6U_10U_4_land_lpi_1_dfm_5 , FpMul_6U_10U_1_and_6_ssc , IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0});
  assign IsNaN_8U_23U_3_nor_3_tmp = ~((FpAdd_8U_23U_o_mant_lpi_1_dfm_2_mx2!=23'b00000000000000000000000));
  assign inp_lookup_1_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp = ({FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_3_5_mx1w1
      , FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_3_4_mx1w1 , FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_3_3_0_mx1w1})
      == ({FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_5_1 , FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_4_1
      , FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_3_0_1});
  assign inp_lookup_2_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp = ({FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_3_5_mx1w1
      , FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_3_4_mx1w1 , FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_3_3_0_mx1w1})
      == ({FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_5_1 , FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_4_1
      , FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_3_0_1});
  assign inp_lookup_3_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp = ({FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_5_mx1w1
      , FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_4_mx1w1 , FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_3_0_mx1w1})
      == ({FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_5_1 , FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_4_1
      , FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_3_0_1});
  assign inp_lookup_4_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp = ({FpMul_6U_10U_1_o_expo_lpi_1_dfm_3_5_mx0w1
      , FpMul_6U_10U_1_o_expo_lpi_1_dfm_3_4_mx0w1 , FpMul_6U_10U_1_o_expo_lpi_1_dfm_3_3_0_mx0w1})
      == ({FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_5_1 , FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_4_1
      , FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_3_0_1});
  assign nl_inp_lookup_1_FpNormalize_8U_49U_1_else_acc_nl = reg_FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_7_1_itm
      + ({2'b11 , (~ libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_12)})
      + 8'b1;
  assign inp_lookup_1_FpNormalize_8U_49U_1_else_acc_nl = nl_inp_lookup_1_FpNormalize_8U_49U_1_else_acc_nl[7:0];
  assign FpNormalize_8U_49U_1_FpNormalize_8U_49U_1_and_nl = MUX_v_8_2_2(8'b00000000,
      (inp_lookup_1_FpNormalize_8U_49U_1_else_acc_nl), FpNormalize_8U_49U_1_oelse_not_9);
  assign nl_inp_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_nl = reg_FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_7_1_itm
      + 8'b1;
  assign inp_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_nl = nl_inp_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_nl[7:0];
  assign FpAdd_8U_23U_1_and_4_nl = (~ inp_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_1_itm_7_1)
      & (FpAdd_8U_23U_1_int_mant_p1_1_sva_3[49]);
  assign FpAdd_8U_23U_1_and_5_nl = inp_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_1_itm_7_1
      & (FpAdd_8U_23U_1_int_mant_p1_1_sva_3[49]);
  assign FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_2_mx0w0 = MUX1HOT_v_8_3_2((FpNormalize_8U_49U_1_FpNormalize_8U_49U_1_and_nl),
      reg_FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_7_1_itm, (inp_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_nl),
      {(~ (FpAdd_8U_23U_1_int_mant_p1_1_sva_3[49])) , (FpAdd_8U_23U_1_and_4_nl) ,
      (FpAdd_8U_23U_1_and_5_nl)});
  assign inp_lookup_1_FpMantRNE_49U_24U_1_else_and_tmp = FpMantRNE_49U_24U_1_else_carry_1_sva_mx0w2
      & (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign FpAdd_6U_10U_1_is_a_greater_oelse_FpAdd_6U_10U_1_is_a_greater_oelse_and_cse
      = (~ FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_itm_10) & IsNaN_8U_23U_2_land_1_lpi_1_dfm_9;
  assign FpAdd_6U_10U_1_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0 = FpAdd_6U_10U_1_is_a_greater_oelse_FpAdd_6U_10U_1_is_a_greater_oelse_and_cse
      | IsNaN_8U_23U_3_land_1_lpi_1_dfm_6;
  assign nl_inp_lookup_2_FpNormalize_8U_49U_1_else_acc_nl = reg_FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_7_1_itm
      + ({2'b11 , (~ libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_13)})
      + 8'b1;
  assign inp_lookup_2_FpNormalize_8U_49U_1_else_acc_nl = nl_inp_lookup_2_FpNormalize_8U_49U_1_else_acc_nl[7:0];
  assign FpNormalize_8U_49U_1_FpNormalize_8U_49U_1_and_2_nl = MUX_v_8_2_2(8'b00000000,
      (inp_lookup_2_FpNormalize_8U_49U_1_else_acc_nl), FpNormalize_8U_49U_1_oelse_not_11);
  assign nl_inp_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_nl = reg_FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_7_1_itm
      + 8'b1;
  assign inp_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_nl = nl_inp_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_nl[7:0];
  assign FpAdd_8U_23U_1_and_10_nl = (~ inp_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_1_itm_7_1)
      & (FpAdd_8U_23U_1_int_mant_p1_2_sva_3[49]);
  assign FpAdd_8U_23U_1_and_11_nl = inp_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_1_itm_7_1
      & (FpAdd_8U_23U_1_int_mant_p1_2_sva_3[49]);
  assign FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_2_mx0w0 = MUX1HOT_v_8_3_2((FpNormalize_8U_49U_1_FpNormalize_8U_49U_1_and_2_nl),
      reg_FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_7_1_itm, (inp_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_nl),
      {(~ (FpAdd_8U_23U_1_int_mant_p1_2_sva_3[49])) , (FpAdd_8U_23U_1_and_10_nl)
      , (FpAdd_8U_23U_1_and_11_nl)});
  assign inp_lookup_2_FpMantRNE_49U_24U_1_else_and_tmp = FpMantRNE_49U_24U_1_else_carry_2_sva_mx0w2
      & (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign FpAdd_6U_10U_1_is_a_greater_oelse_FpAdd_6U_10U_1_is_a_greater_oelse_and_1_cse
      = (~ FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_1_itm_10) & IsNaN_8U_23U_2_land_2_lpi_1_dfm_9;
  assign FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0 = FpAdd_6U_10U_1_is_a_greater_oelse_FpAdd_6U_10U_1_is_a_greater_oelse_and_1_cse
      | IsNaN_8U_23U_3_land_2_lpi_1_dfm_6;
  assign nl_inp_lookup_3_FpNormalize_8U_49U_1_else_acc_nl = reg_FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_7_1_itm
      + ({2'b11 , (~ libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_14)})
      + 8'b1;
  assign inp_lookup_3_FpNormalize_8U_49U_1_else_acc_nl = nl_inp_lookup_3_FpNormalize_8U_49U_1_else_acc_nl[7:0];
  assign FpNormalize_8U_49U_1_FpNormalize_8U_49U_1_and_4_nl = MUX_v_8_2_2(8'b00000000,
      (inp_lookup_3_FpNormalize_8U_49U_1_else_acc_nl), FpNormalize_8U_49U_1_oelse_not_13);
  assign nl_inp_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_nl = reg_FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_7_1_itm
      + 8'b1;
  assign inp_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_nl = nl_inp_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_nl[7:0];
  assign FpAdd_8U_23U_1_and_16_nl = (~ inp_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_1_itm_7)
      & (FpAdd_8U_23U_1_int_mant_p1_3_sva_3[49]);
  assign FpAdd_8U_23U_1_and_17_nl = inp_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_1_itm_7
      & (FpAdd_8U_23U_1_int_mant_p1_3_sva_3[49]);
  assign FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_2_mx0w0 = MUX1HOT_v_8_3_2((FpNormalize_8U_49U_1_FpNormalize_8U_49U_1_and_4_nl),
      reg_FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_7_1_itm, (inp_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_nl),
      {(~ (FpAdd_8U_23U_1_int_mant_p1_3_sva_3[49])) , (FpAdd_8U_23U_1_and_16_nl)
      , (FpAdd_8U_23U_1_and_17_nl)});
  assign inp_lookup_3_FpMantRNE_49U_24U_1_else_and_tmp = FpMantRNE_49U_24U_1_else_carry_3_sva_mx0w2
      & (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign FpAdd_6U_10U_1_is_a_greater_oelse_FpAdd_6U_10U_1_is_a_greater_oelse_and_2_cse
      = (~ FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_2_itm_10) & IsNaN_8U_23U_2_land_3_lpi_1_dfm_9;
  assign FpAdd_6U_10U_1_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0 = FpAdd_6U_10U_1_is_a_greater_oelse_FpAdd_6U_10U_1_is_a_greater_oelse_and_2_cse
      | IsNaN_8U_23U_3_land_3_lpi_1_dfm_6;
  assign nl_inp_lookup_4_FpNormalize_8U_49U_1_else_acc_nl = reg_FpMul_6U_10U_2_o_mant_lpi_1_dfm_7_1_reg
      + ({2'b11 , (~ libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_15)})
      + 8'b1;
  assign inp_lookup_4_FpNormalize_8U_49U_1_else_acc_nl = nl_inp_lookup_4_FpNormalize_8U_49U_1_else_acc_nl[7:0];
  assign FpNormalize_8U_49U_1_FpNormalize_8U_49U_1_and_6_nl = MUX_v_8_2_2(8'b00000000,
      (inp_lookup_4_FpNormalize_8U_49U_1_else_acc_nl), FpNormalize_8U_49U_1_oelse_not_15);
  assign nl_inp_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_nl = reg_FpMul_6U_10U_2_o_mant_lpi_1_dfm_7_1_reg
      + 8'b1;
  assign inp_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_nl = nl_inp_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_nl[7:0];
  assign FpAdd_8U_23U_1_and_22_nl = (~ inp_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_1_itm_7_1)
      & (FpAdd_8U_23U_1_int_mant_p1_sva_3[49]);
  assign FpAdd_8U_23U_1_and_23_nl = inp_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_1_itm_7_1
      & (FpAdd_8U_23U_1_int_mant_p1_sva_3[49]);
  assign FpAdd_8U_23U_1_o_expo_lpi_1_dfm_2_mx0w0 = MUX1HOT_v_8_3_2((FpNormalize_8U_49U_1_FpNormalize_8U_49U_1_and_6_nl),
      reg_FpMul_6U_10U_2_o_mant_lpi_1_dfm_7_1_reg, (inp_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_nl),
      {(~ (FpAdd_8U_23U_1_int_mant_p1_sva_3[49])) , (FpAdd_8U_23U_1_and_22_nl) ,
      (FpAdd_8U_23U_1_and_23_nl)});
  assign inp_lookup_4_FpMantRNE_49U_24U_1_else_and_tmp = FpMantRNE_49U_24U_1_else_carry_sva_mx0w2
      & (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign FpAdd_6U_10U_1_is_a_greater_lor_lpi_1_dfm_1_mx0w0 = ((~ FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_3_itm_10)
      & IsNaN_8U_23U_2_land_lpi_1_dfm_9) | IsNaN_8U_23U_3_land_lpi_1_dfm_5;
  assign nl_inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_nl = ({1'b1
      , (~ FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_7_mx0w0)}) + 9'b1100001;
  assign inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_nl = nl_inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_nl[8:0];
  assign inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8 = readslicef_9_1_8((inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_nl));
  assign inp_lookup_1_FpMantRNE_24U_11U_else_and_svs_mx0w0 = FpMantRNE_24U_11U_else_carry_1_sva
      & (FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_2_mx1[22:13]==10'b1111111111);
  assign nl_inp_lookup_1_FpMantRNE_49U_24U_1_else_acc_nl = reg_chn_inp_in_crt_sva_6_30_0_1_reg
      + conv_u2u_1_23(FpAdd_6U_10U_1_qr_2_lpi_1_dfm_3_5_1);
  assign inp_lookup_1_FpMantRNE_49U_24U_1_else_acc_nl = nl_inp_lookup_1_FpMantRNE_49U_24U_1_else_acc_nl[22:0];
  assign FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_4_itm = MUX_v_23_2_2((inp_lookup_1_FpMantRNE_49U_24U_1_else_acc_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_2_mx0);
  assign nl_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_2_sva_mx0w0
      = (~ (FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_7_mx0w0[3:1])) + 3'b1;
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_2_sva_mx0w0
      = nl_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_2_sva_mx0w0[2:0];
  assign nl_inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_nl = conv_u2u_7_8(FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_7_mx0w0[7:1])
      + 8'b11010101;
  assign inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_nl = nl_inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_nl[7:0];
  assign inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7 = readslicef_8_1_7((inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_nl));
  assign nl_inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_nl = conv_u2s_8_9(FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_7_mx0w0)
      + 9'b101100001;
  assign inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_nl = nl_inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_nl[8:0];
  assign inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8 = readslicef_9_1_8((inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_nl));
  assign inp_lookup_2_FpMantRNE_24U_11U_else_and_svs_mx0w0 = FpMantRNE_24U_11U_else_carry_2_sva_mx0w1
      & (FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_2_mx1[22:13]==10'b1111111111);
  assign nl_inp_lookup_2_FpMantRNE_49U_24U_1_else_acc_nl = reg_chn_inp_in_crt_sva_6_62_32_1_reg
      + conv_u2u_1_23(FpAdd_6U_10U_1_qr_3_lpi_1_dfm_3_5_1);
  assign inp_lookup_2_FpMantRNE_49U_24U_1_else_acc_nl = nl_inp_lookup_2_FpMantRNE_49U_24U_1_else_acc_nl[22:0];
  assign FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_5_itm = MUX_v_23_2_2((inp_lookup_2_FpMantRNE_49U_24U_1_else_acc_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_2_mx0);
  assign nl_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_3_sva_mx0w0
      = (~ (FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_7[3:1])) + 3'b1;
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_3_sva_mx0w0
      = nl_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_3_sva_mx0w0[2:0];
  assign nl_inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_nl = ({1'b1
      , (~ FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_7)}) + 9'b1100001;
  assign inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_nl = nl_inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_nl[8:0];
  assign inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8 = readslicef_9_1_8((inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_nl));
  assign nl_inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_nl = conv_u2u_7_8(FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_7[7:1])
      + 8'b11010101;
  assign inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_nl = nl_inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_nl[7:0];
  assign inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7 = readslicef_8_1_7((inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_nl));
  assign nl_inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_nl = conv_u2s_8_9(FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_7)
      + 9'b101100001;
  assign inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_nl = nl_inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_nl[8:0];
  assign inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8 = readslicef_9_1_8((inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_nl));
  assign IsNaN_8U_23U_4_IsNaN_8U_23U_4_nor_1_tmp = ~((~((FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_2_mx1!=23'b00000000000000000000000)))
      | (FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_7!=8'b11111111));
  assign inp_lookup_3_FpMantRNE_24U_11U_else_and_svs_mx0w0 = FpMantRNE_24U_11U_else_carry_3_sva_mx0w1
      & (FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx1[22:13]==10'b1111111111);
  assign nl_inp_lookup_3_FpMantRNE_49U_24U_1_else_acc_nl = reg_chn_inp_in_crt_sva_6_94_64_1_reg
      + conv_u2u_1_23(FpAdd_6U_10U_1_qr_4_lpi_1_dfm_3_5_1);
  assign inp_lookup_3_FpMantRNE_49U_24U_1_else_acc_nl = nl_inp_lookup_3_FpMantRNE_49U_24U_1_else_acc_nl[22:0];
  assign FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_6_nl = MUX_v_23_2_2((inp_lookup_3_FpMantRNE_49U_24U_1_else_acc_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_2_mx0);
  assign FpAdd_8U_23U_1_asn_40_mx0w1 = MUX_v_23_2_2((FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_6_nl),
      FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2, IsNaN_8U_23U_3_land_3_lpi_1_dfm_7);
  assign nl_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_4_sva_mx0w0
      = (~ (FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_7[3:1])) + 3'b1;
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_4_sva_mx0w0
      = nl_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_4_sva_mx0w0[2:0];
  assign nl_inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_nl = ({1'b1
      , (~ FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_7)}) + 9'b1100001;
  assign inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_nl = nl_inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_nl[8:0];
  assign inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8 = readslicef_9_1_8((inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_nl));
  assign nl_inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_nl = conv_u2u_7_8(FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_7[7:1])
      + 8'b11010101;
  assign inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_nl = nl_inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_nl[7:0];
  assign inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7 = readslicef_8_1_7((inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_nl));
  assign nl_inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_nl = conv_u2s_8_9(FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_7)
      + 9'b101100001;
  assign inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_nl = nl_inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_nl[8:0];
  assign inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8 = readslicef_9_1_8((inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_nl));
  assign IsNaN_8U_23U_4_IsNaN_8U_23U_4_nor_2_tmp = ~((~((FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx1!=23'b00000000000000000000000)))
      | (FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_7!=8'b11111111));
  assign inp_lookup_4_FpMantRNE_24U_11U_else_and_svs_mx0w0 = FpMantRNE_24U_11U_else_carry_sva_mx0w1
      & (FpAdd_8U_23U_1_o_mant_lpi_1_dfm_2_mx1[22:13]==10'b1111111111);
  assign nl_inp_lookup_4_FpMantRNE_49U_24U_1_else_acc_nl = reg_chn_inp_in_crt_sva_6_126_96_1_reg
      + conv_u2u_1_23(FpAdd_6U_10U_1_qr_lpi_1_dfm_3_5_1);
  assign inp_lookup_4_FpMantRNE_49U_24U_1_else_acc_nl = nl_inp_lookup_4_FpMantRNE_49U_24U_1_else_acc_nl[22:0];
  assign FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_7_itm = MUX_v_23_2_2((inp_lookup_4_FpMantRNE_49U_24U_1_else_acc_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_1_is_inf_lpi_1_dfm_2_mx0);
  assign nl_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_1_sva_mx0w0
      = (~ (FpAdd_8U_23U_1_o_expo_lpi_1_dfm_7[3:1])) + 3'b1;
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_1_sva_mx0w0
      = nl_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_1_sva_mx0w0[2:0];
  assign nl_inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_nl = ({1'b1
      , (~ FpAdd_8U_23U_1_o_expo_lpi_1_dfm_7)}) + 9'b1100001;
  assign inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_nl = nl_inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_nl[8:0];
  assign inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8 = readslicef_9_1_8((inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_nl));
  assign nl_inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_nl = conv_u2u_7_8(FpAdd_8U_23U_1_o_expo_lpi_1_dfm_7[7:1])
      + 8'b11010101;
  assign inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_nl = nl_inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_nl[7:0];
  assign inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7 = readslicef_8_1_7((inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_nl));
  assign nl_inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_nl = conv_u2s_8_9(FpAdd_8U_23U_1_o_expo_lpi_1_dfm_7)
      + 9'b101100001;
  assign inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_nl = nl_inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_nl[8:0];
  assign inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8 = readslicef_9_1_8((inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_nl));
  assign IsNaN_8U_23U_4_IsNaN_8U_23U_4_nor_3_tmp = ~((~((FpAdd_8U_23U_1_o_mant_lpi_1_dfm_2_mx1!=23'b00000000000000000000000)))
      | (FpAdd_8U_23U_1_o_expo_lpi_1_dfm_7!=8'b11111111));
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_else_mux_8_nl = MUX_s_1_2_2((~
      (FpAdd_6U_10U_1_qr_2_lpi_1_dfm_5[5])), (FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_sva_3[5]),
      inp_lookup_1_FpMantRNE_24U_11U_else_and_svs_2);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_7_5_mx0w0 = ((FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_else_mux_8_nl)
      & (~ FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_nor_ssc))
      | FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_1_lpi_1_dfm_3 | nor_1727_cse;
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_and_11_nl = (~ inp_lookup_1_FpMantRNE_24U_11U_else_and_svs_2)
      & FpWidthDec_8U_23U_6U_10U_0U_1U_and_1_m1c;
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_and_12_nl = inp_lookup_1_FpMantRNE_24U_11U_else_and_svs_2
      & FpWidthDec_8U_23U_6U_10U_0U_1U_and_1_m1c;
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_mux1h_nl =
      MUX1HOT_v_5_4_2(5'b1, (FpAdd_6U_10U_1_qr_2_lpi_1_dfm_5[4:0]), (FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_sva_3[4:0]),
      5'b11110, {FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_nor_ssc
      , (FpWidthDec_8U_23U_6U_10U_0U_1U_and_11_nl) , (FpWidthDec_8U_23U_6U_10U_0U_1U_and_12_nl)
      , FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_1_lpi_1_dfm_3});
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_not_8_nl = ~ FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_1_lpi_1_dfm_2;
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_and_nl
      = MUX_v_5_2_2(5'b00000, (FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_mux1h_nl),
      (FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_not_8_nl));
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_7_4_0_mx0w0 = MUX_v_5_2_2((FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_and_nl),
      5'b11111, nor_1727_cse);
  assign FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_tmp = FpNormalize_6U_23U_1_if_or_itm_2
      | (~((FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_1_lpi_1_dfm_5_mx1!=10'b0000000000)
      | FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_7_5_mx0w0 | (FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_7_4_0_mx0w0!=5'b00000)));
  assign FpAdd_6U_10U_1_or_12_cse = IsNaN_6U_10U_9_land_1_lpi_1_dfm_8 | IsNaN_6U_10U_8_land_1_lpi_1_dfm_7;
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_14_nl = MUX1HOT_s_1_3_2(FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_5,
      (FpAdd_6U_10U_1_o_expo_1_sva_4[5]), FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_8_5_1,
      {FpAdd_6U_10U_1_and_ssc , FpAdd_6U_10U_1_and_6_ssc , FpAdd_6U_10U_1_or_12_cse});
  assign FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_5_mx0w0 = (FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_14_nl)
      | FpAdd_6U_10U_1_and_28_ssc;
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_2_nl = MUX1HOT_s_1_3_2(FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_4,
      (FpAdd_6U_10U_1_o_expo_1_sva_4[4]), FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_8_4_1,
      {FpAdd_6U_10U_1_and_ssc , FpAdd_6U_10U_1_and_6_ssc , FpAdd_6U_10U_1_or_12_cse});
  assign FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_4_mx0w0 = (FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_2_nl)
      | FpAdd_6U_10U_1_and_28_ssc;
  assign FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_3_0_mx0w0 = MUX1HOT_v_4_4_2(FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_3_0,
      (FpAdd_6U_10U_1_o_expo_1_sva_4[3:0]), 4'b1110, ({reg_FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_8_3_0_itm
      , reg_FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_8_3_0_1_itm}), {FpAdd_6U_10U_1_and_ssc
      , FpAdd_6U_10U_1_and_6_ssc , FpAdd_6U_10U_1_and_28_ssc , FpAdd_6U_10U_1_or_12_cse});
  assign nl_inp_lookup_1_FpMantRNE_23U_11U_1_else_acc_nl = (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_1_else_carry_1_sva);
  assign inp_lookup_1_FpMantRNE_23U_11U_1_else_acc_nl = nl_inp_lookup_1_FpMantRNE_23U_11U_1_else_acc_nl[9:0];
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_itm_mx0w0 = MUX_v_10_2_2((inp_lookup_1_FpMantRNE_23U_11U_1_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_1_is_inf_1_lpi_1_dfm_2_mx0);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_else_mux_9_nl = MUX_s_1_2_2((~
      (FpAdd_6U_10U_1_qr_3_lpi_1_dfm_5[5])), (FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_sva_3[5]),
      inp_lookup_2_FpMantRNE_24U_11U_else_and_svs_2);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_7_5_mx0w0 = ((FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_else_mux_9_nl)
      & (~ FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_nor_1_ssc))
      | FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_2_lpi_1_dfm_3 | IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_5;
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_and_13_nl = (~ inp_lookup_2_FpMantRNE_24U_11U_else_and_svs_2)
      & FpWidthDec_8U_23U_6U_10U_0U_1U_and_3_m1c;
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_and_14_nl = inp_lookup_2_FpMantRNE_24U_11U_else_and_svs_2
      & FpWidthDec_8U_23U_6U_10U_0U_1U_and_3_m1c;
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_mux1h_1_nl
      = MUX1HOT_v_5_4_2(5'b1, (FpAdd_6U_10U_1_qr_3_lpi_1_dfm_5[4:0]), (FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_sva_3[4:0]),
      5'b11110, {FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_nor_1_ssc
      , (FpWidthDec_8U_23U_6U_10U_0U_1U_and_13_nl) , (FpWidthDec_8U_23U_6U_10U_0U_1U_and_14_nl)
      , FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_2_lpi_1_dfm_3});
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_not_9_nl = ~ FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_2_lpi_1_dfm_2;
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_and_2_nl
      = MUX_v_5_2_2(5'b00000, (FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_mux1h_1_nl),
      (FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_not_9_nl));
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_7_4_0_mx0w0 = MUX_v_5_2_2((FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_and_2_nl),
      5'b11111, IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_5);
  assign FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_2_tmp = FpNormalize_6U_23U_1_if_or_1_itm_2
      | (~((FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_2_lpi_1_dfm_5_mx0!=10'b0000000000)
      | FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_7_5_mx0w0 | (FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_7_4_0_mx0w0!=5'b00000)));
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_17_nl = MUX1HOT_s_1_3_2(FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_5,
      (FpAdd_6U_10U_1_o_expo_2_sva_4[5]), FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_8_5_1,
      {FpAdd_6U_10U_1_and_29_ssc , FpAdd_6U_10U_1_and_13_ssc , or_5680_cse});
  assign FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_5_mx0w0 = (FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_17_nl)
      | FpAdd_6U_10U_1_and_30_ssc;
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_5_nl = MUX1HOT_s_1_3_2(FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_4,
      (FpAdd_6U_10U_1_o_expo_2_sva_4[4]), FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_8_4_1,
      {FpAdd_6U_10U_1_and_29_ssc , FpAdd_6U_10U_1_and_13_ssc , or_5680_cse});
  assign FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_4_mx0w0 = (FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_5_nl)
      | FpAdd_6U_10U_1_and_30_ssc;
  assign FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_3_0_mx0w0 = MUX1HOT_v_4_4_2(FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_3_0,
      (FpAdd_6U_10U_1_o_expo_2_sva_4[3:0]), 4'b1110, ({reg_FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_8_3_0_itm
      , reg_FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_8_3_0_1_itm}), {FpAdd_6U_10U_1_and_29_ssc
      , FpAdd_6U_10U_1_and_13_ssc , FpAdd_6U_10U_1_and_30_ssc , or_5680_cse});
  assign nl_inp_lookup_2_FpMantRNE_23U_11U_1_else_acc_nl = (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_1_else_carry_2_sva);
  assign inp_lookup_2_FpMantRNE_23U_11U_1_else_acc_nl = nl_inp_lookup_2_FpMantRNE_23U_11U_1_else_acc_nl[9:0];
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_1_itm_mx0w0 = MUX_v_10_2_2((inp_lookup_2_FpMantRNE_23U_11U_1_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_1_is_inf_2_lpi_1_dfm_2_mx0);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_else_mux_10_nl = MUX_s_1_2_2((~
      (FpAdd_6U_10U_1_qr_4_lpi_1_dfm_5[5])), (FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_sva_3[5]),
      inp_lookup_3_FpMantRNE_24U_11U_else_and_svs_2);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_7_5_mx0w0 = ((FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_else_mux_10_nl)
      & (~ FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_nor_2_ssc))
      | FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_3_lpi_1_dfm_3 | IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_5;
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_and_15_nl = (~ inp_lookup_3_FpMantRNE_24U_11U_else_and_svs_2)
      & FpWidthDec_8U_23U_6U_10U_0U_1U_and_5_m1c;
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_and_16_nl = inp_lookup_3_FpMantRNE_24U_11U_else_and_svs_2
      & FpWidthDec_8U_23U_6U_10U_0U_1U_and_5_m1c;
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_mux1h_2_nl
      = MUX1HOT_v_5_4_2(5'b1, (FpAdd_6U_10U_1_qr_4_lpi_1_dfm_5[4:0]), (FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_sva_3[4:0]),
      5'b11110, {FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_nor_2_ssc
      , (FpWidthDec_8U_23U_6U_10U_0U_1U_and_15_nl) , (FpWidthDec_8U_23U_6U_10U_0U_1U_and_16_nl)
      , FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_3_lpi_1_dfm_3});
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_not_10_nl = ~ FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_3_lpi_1_dfm_2;
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_and_4_nl
      = MUX_v_5_2_2(5'b00000, (FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_mux1h_2_nl),
      (FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_not_10_nl));
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_7_4_0_mx0w0 = MUX_v_5_2_2((FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_and_4_nl),
      5'b11111, IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_5);
  assign FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_4_tmp = FpNormalize_6U_23U_1_if_or_2_itm_2
      | (~((FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_3_lpi_1_dfm_5_mx0!=10'b0000000000)
      | FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_7_5_mx0w0 | (FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_7_4_0_mx0w0!=5'b00000)));
  assign FpAdd_6U_10U_1_or_16_cse = IsNaN_6U_10U_9_land_3_lpi_1_dfm_8 | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_19;
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_20_nl = MUX1HOT_s_1_3_2(FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_5,
      (FpAdd_6U_10U_1_o_expo_3_sva_4[5]), FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_8_5_1,
      {FpAdd_6U_10U_1_and_31_ssc , FpAdd_6U_10U_1_and_19_ssc , FpAdd_6U_10U_1_or_16_cse});
  assign FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_5_mx0w0 = (FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_20_nl)
      | FpAdd_6U_10U_1_and_32_ssc;
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_8_nl = MUX1HOT_s_1_3_2(FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_4,
      (FpAdd_6U_10U_1_o_expo_3_sva_4[4]), FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_8_4_1,
      {FpAdd_6U_10U_1_and_31_ssc , FpAdd_6U_10U_1_and_19_ssc , FpAdd_6U_10U_1_or_16_cse});
  assign FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_4_mx0w0 = (FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_8_nl)
      | FpAdd_6U_10U_1_and_32_ssc;
  assign FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_3_0_mx0w0 = MUX1HOT_v_4_4_2(FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_3_0,
      (FpAdd_6U_10U_1_o_expo_3_sva_4[3:0]), 4'b1110, ({reg_FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_8_3_0_itm
      , reg_FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_8_3_0_1_itm}), {FpAdd_6U_10U_1_and_31_ssc
      , FpAdd_6U_10U_1_and_19_ssc , FpAdd_6U_10U_1_and_32_ssc , FpAdd_6U_10U_1_or_16_cse});
  assign nl_inp_lookup_3_FpMantRNE_23U_11U_1_else_acc_nl = (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_1_else_carry_3_sva);
  assign inp_lookup_3_FpMantRNE_23U_11U_1_else_acc_nl = nl_inp_lookup_3_FpMantRNE_23U_11U_1_else_acc_nl[9:0];
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_2_itm_mx0w0 = MUX_v_10_2_2((inp_lookup_3_FpMantRNE_23U_11U_1_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_1_is_inf_3_lpi_1_dfm_2_mx0);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_else_mux_11_nl = MUX_s_1_2_2((~
      (FpAdd_6U_10U_1_qr_lpi_1_dfm_5[5])), (FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_sva_3[5]),
      inp_lookup_4_FpMantRNE_24U_11U_else_and_svs_2);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_7_5_mx0w0 = ((FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_else_mux_11_nl)
      & (~ FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_nor_3_ssc))
      | FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_lpi_1_dfm_3 | IsNaN_6U_10U_8_land_lpi_1_dfm_st_5;
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_and_17_nl = (~ inp_lookup_4_FpMantRNE_24U_11U_else_and_svs_2)
      & FpWidthDec_8U_23U_6U_10U_0U_1U_and_7_m1c;
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_and_18_nl = inp_lookup_4_FpMantRNE_24U_11U_else_and_svs_2
      & FpWidthDec_8U_23U_6U_10U_0U_1U_and_7_m1c;
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_mux1h_3_nl
      = MUX1HOT_v_5_4_2(5'b1, (FpAdd_6U_10U_1_qr_lpi_1_dfm_5[4:0]), (FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_sva_3[4:0]),
      5'b11110, {FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_nor_3_ssc
      , (FpWidthDec_8U_23U_6U_10U_0U_1U_and_17_nl) , (FpWidthDec_8U_23U_6U_10U_0U_1U_and_18_nl)
      , FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_lpi_1_dfm_3});
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_not_11_nl = ~ FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_lpi_1_dfm_2;
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_and_6_nl
      = MUX_v_5_2_2(5'b00000, (FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_mux1h_3_nl),
      (FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_not_11_nl));
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_7_4_0_mx0w0 = MUX_v_5_2_2((FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_and_6_nl),
      5'b11111, IsNaN_6U_10U_8_land_lpi_1_dfm_st_5);
  assign FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_6_tmp = FpNormalize_6U_23U_1_if_or_3_itm_2
      | (~((FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_lpi_1_dfm_5_mx0!=10'b0000000000)
      | FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_7_5_mx0w0 | (FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_7_4_0_mx0w0!=5'b00000)));
  assign FpAdd_6U_10U_1_or_18_cse = IsNaN_6U_10U_9_land_lpi_1_dfm_8 | IsNaN_6U_10U_2_land_lpi_1_dfm_st_18;
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_23_nl = MUX1HOT_s_1_3_2(FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_5,
      (FpAdd_6U_10U_1_o_expo_sva_4[5]), FpMul_6U_10U_1_o_expo_lpi_1_dfm_8_5_1, {FpAdd_6U_10U_1_and_33_ssc
      , FpAdd_6U_10U_1_and_25_ssc , FpAdd_6U_10U_1_or_18_cse});
  assign FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_5_mx0w0 = (FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_23_nl)
      | FpAdd_6U_10U_1_and_34_ssc;
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_11_nl = MUX1HOT_s_1_3_2(FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_4,
      (FpAdd_6U_10U_1_o_expo_sva_4[4]), FpMul_6U_10U_1_o_expo_lpi_1_dfm_8_4_1, {FpAdd_6U_10U_1_and_33_ssc
      , FpAdd_6U_10U_1_and_25_ssc , FpAdd_6U_10U_1_or_18_cse});
  assign FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_4_mx0w0 = (FpAdd_6U_10U_1_FpAdd_6U_10U_1_mux1h_11_nl)
      | FpAdd_6U_10U_1_and_34_ssc;
  assign FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_3_0_mx0w0 = MUX1HOT_v_4_4_2(FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_3_0,
      (FpAdd_6U_10U_1_o_expo_sva_4[3:0]), 4'b1110, ({reg_FpMul_6U_10U_1_o_expo_lpi_1_dfm_8_3_0_itm
      , reg_FpMul_6U_10U_1_o_expo_lpi_1_dfm_8_3_0_1_itm}), {FpAdd_6U_10U_1_and_33_ssc
      , FpAdd_6U_10U_1_and_25_ssc , FpAdd_6U_10U_1_and_34_ssc , FpAdd_6U_10U_1_or_18_cse});
  assign nl_inp_lookup_4_FpMantRNE_23U_11U_1_else_acc_nl = (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_1_else_carry_sva);
  assign inp_lookup_4_FpMantRNE_23U_11U_1_else_acc_nl = nl_inp_lookup_4_FpMantRNE_23U_11U_1_else_acc_nl[9:0];
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_3_itm_mx0w0 = MUX_v_10_2_2((inp_lookup_4_FpMantRNE_23U_11U_1_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_1_is_inf_lpi_1_dfm_2_mx0);
  assign nl_inp_lookup_1_FpMul_6U_10U_else_2_acc_1_nl = conv_u2u_6_7({FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_10_5_1
      , FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_10_4_0_1}) + conv_u2u_6_7({FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_13_1_1
      , FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_5_1 , FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_3_0_1});
  assign inp_lookup_1_FpMul_6U_10U_else_2_acc_1_nl = nl_inp_lookup_1_FpMul_6U_10U_else_2_acc_1_nl[6:0];
  assign nl_inp_lookup_1_FpMul_6U_10U_else_2_if_acc_nl = conv_u2u_6_7(readslicef_7_6_1((inp_lookup_1_FpMul_6U_10U_else_2_acc_1_nl)))
      + 7'b1010001;
  assign inp_lookup_1_FpMul_6U_10U_else_2_if_acc_nl = nl_inp_lookup_1_FpMul_6U_10U_else_2_if_acc_nl[6:0];
  assign inp_lookup_1_FpMul_6U_10U_else_2_if_acc_itm_6_1 = readslicef_7_1_6((inp_lookup_1_FpMul_6U_10U_else_2_if_acc_nl));
  assign inp_lookup_1_FpMul_6U_10U_p_mant_p1_mul_tmp = conv_u2u_22_22(({1'b1 , FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_1_lpi_1_dfm_9})
      * ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_22}));
  assign nl_inp_lookup_2_FpMul_6U_10U_else_2_acc_1_nl = conv_u2u_6_7({FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_10_5_1
      , FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_10_4_0_1}) + conv_u2u_6_7({FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_13_1_1
      , FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_5_1 , FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_3_0_1});
  assign inp_lookup_2_FpMul_6U_10U_else_2_acc_1_nl = nl_inp_lookup_2_FpMul_6U_10U_else_2_acc_1_nl[6:0];
  assign nl_inp_lookup_2_FpMul_6U_10U_else_2_if_acc_nl = conv_u2u_6_7(readslicef_7_6_1((inp_lookup_2_FpMul_6U_10U_else_2_acc_1_nl)))
      + 7'b1010001;
  assign inp_lookup_2_FpMul_6U_10U_else_2_if_acc_nl = nl_inp_lookup_2_FpMul_6U_10U_else_2_if_acc_nl[6:0];
  assign inp_lookup_2_FpMul_6U_10U_else_2_if_acc_itm_6_1 = readslicef_7_1_6((inp_lookup_2_FpMul_6U_10U_else_2_if_acc_nl));
  assign inp_lookup_2_FpMul_6U_10U_p_mant_p1_mul_tmp = conv_u2u_22_22(({1'b1 , FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_2_lpi_1_dfm_9})
      * ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_22}));
  assign nl_inp_lookup_3_FpMul_6U_10U_else_2_acc_1_nl = conv_u2u_6_7({FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_10_5_1
      , FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_10_4_0_1}) + conv_u2u_6_7({FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_13_1_1
      , FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_5_1 , FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_3_0_1});
  assign inp_lookup_3_FpMul_6U_10U_else_2_acc_1_nl = nl_inp_lookup_3_FpMul_6U_10U_else_2_acc_1_nl[6:0];
  assign nl_inp_lookup_3_FpMul_6U_10U_else_2_if_acc_nl = conv_u2u_6_7(readslicef_7_6_1((inp_lookup_3_FpMul_6U_10U_else_2_acc_1_nl)))
      + 7'b1010001;
  assign inp_lookup_3_FpMul_6U_10U_else_2_if_acc_nl = nl_inp_lookup_3_FpMul_6U_10U_else_2_if_acc_nl[6:0];
  assign inp_lookup_3_FpMul_6U_10U_else_2_if_acc_itm_6_1 = readslicef_7_1_6((inp_lookup_3_FpMul_6U_10U_else_2_if_acc_nl));
  assign inp_lookup_3_FpMul_6U_10U_p_mant_p1_mul_tmp = conv_u2u_22_22(({1'b1 , FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_3_lpi_1_dfm_9})
      * ({1'b1 , FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_2_itm_2}));
  assign nl_inp_lookup_4_FpMul_6U_10U_else_2_acc_1_nl = conv_u2u_6_7({FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_10_5_1
      , FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_10_4_0_1}) + conv_u2u_6_7({FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_13_1_1
      , FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_5_1 , FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_3_0_1});
  assign inp_lookup_4_FpMul_6U_10U_else_2_acc_1_nl = nl_inp_lookup_4_FpMul_6U_10U_else_2_acc_1_nl[6:0];
  assign nl_inp_lookup_4_FpMul_6U_10U_else_2_if_acc_nl = conv_u2u_6_7(readslicef_7_6_1((inp_lookup_4_FpMul_6U_10U_else_2_acc_1_nl)))
      + 7'b1010001;
  assign inp_lookup_4_FpMul_6U_10U_else_2_if_acc_nl = nl_inp_lookup_4_FpMul_6U_10U_else_2_if_acc_nl[6:0];
  assign inp_lookup_4_FpMul_6U_10U_else_2_if_acc_itm_6_1 = readslicef_7_1_6((inp_lookup_4_FpMul_6U_10U_else_2_if_acc_nl));
  assign inp_lookup_4_FpMul_6U_10U_p_mant_p1_mul_tmp = conv_u2u_22_22(({1'b1 , FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_lpi_1_dfm_9})
      * ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_22}));
  assign inp_lookup_1_FpAdd_6U_10U_is_a_greater_oif_equal_tmp = ({reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_15_tmp
      , reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_15_tmp_1 , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_27})
      == ({reg_FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_5_4_tmp , reg_FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_5_4_tmp_1
      , FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_3_0_1});
  assign nl_inp_lookup_1_FpMantRNE_22U_11U_else_acc_nl = (FpMul_6U_10U_p_mant_20_1_1_lpi_1_dfm_3_mx0[19:10])
      + conv_u2u_1_10(FpMantRNE_22U_11U_else_carry_1_sva);
  assign inp_lookup_1_FpMantRNE_22U_11U_else_acc_nl = nl_inp_lookup_1_FpMantRNE_22U_11U_else_acc_nl[9:0];
  assign or_5850_nl = FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp | (~ inp_lookup_1_FpMantRNE_22U_11U_else_and_svs);
  assign mux_2025_nl = MUX_v_10_2_2((signext_10_1(~ FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp)),
      (inp_lookup_1_FpMantRNE_22U_11U_else_acc_nl), or_5850_nl);
  assign FpMul_6U_10U_nor_nl = ~(MUX_v_10_2_2((mux_2025_nl), 10'b1111111111, FpMul_6U_10U_is_inf_1_lpi_1_dfm_2));
  assign FpMul_6U_10U_FpMul_6U_10U_FpMul_6U_10U_nor_4_nl = ~(MUX_v_10_2_2((FpMul_6U_10U_nor_nl),
      10'b1111111111, FpMul_6U_10U_lor_9_lpi_1_dfm));
  assign FpMul_6U_10U_or_8_nl = FpMul_6U_10U_and_ssc | IsNaN_6U_10U_land_1_lpi_1_dfm_6;
  assign FpMul_6U_10U_o_mant_1_lpi_1_dfm_3_mx0w0 = MUX_v_10_2_2((FpMul_6U_10U_FpMul_6U_10U_FpMul_6U_10U_nor_4_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_23, FpMul_6U_10U_or_8_nl);
  assign FpMul_6U_10U_oelse_2_not_27_nl = ~ FpMul_6U_10U_lor_9_lpi_1_dfm;
  assign FpMul_6U_10U_FpMul_6U_10U_and_15_nl = MUX_v_4_2_2(4'b0000, (FpMul_6U_10U_o_expo_1_lpi_1_dfm[3:0]),
      (FpMul_6U_10U_oelse_2_not_27_nl));
  assign FpMul_6U_10U_o_expo_1_lpi_1_dfm_3_3_0_mx0w0 = MUX1HOT_v_4_3_2((FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_11_4_0_1[3:0]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_22, (FpMul_6U_10U_FpMul_6U_10U_and_15_nl),
      {IsNaN_6U_10U_land_1_lpi_1_dfm_6 , FpMul_6U_10U_and_ssc , FpMul_6U_10U_FpMul_6U_10U_nor_ssc});
  assign nl_FpAdd_6U_10U_is_a_greater_acc_nl = ({1'b1 , FpMul_6U_10U_o_expo_1_lpi_1_dfm_3_5_mx0w0
      , FpMul_6U_10U_o_expo_1_lpi_1_dfm_3_4_mx0w0 , FpMul_6U_10U_o_expo_1_lpi_1_dfm_3_3_0_mx0w0})
      + conv_u2u_6_7({(~ FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_14_1_1)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_14_0_1) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_26)})
      + 7'b1;
  assign FpAdd_6U_10U_is_a_greater_acc_nl = nl_FpAdd_6U_10U_is_a_greater_acc_nl[6:0];
  assign FpAdd_6U_10U_is_a_greater_acc_itm_6_1 = readslicef_7_1_6((FpAdd_6U_10U_is_a_greater_acc_nl));
  assign inp_lookup_2_FpAdd_6U_10U_is_a_greater_oif_equal_tmp = ({reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_15_tmp
      , reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_15_tmp_1 , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_27})
      == ({reg_FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_5_4_tmp , reg_FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_5_4_tmp_1
      , FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_3_0_1});
  assign nl_inp_lookup_2_FpMantRNE_22U_11U_else_acc_nl = (FpMul_6U_10U_p_mant_20_1_2_lpi_1_dfm_3_mx0[19:10])
      + conv_u2u_1_10(FpMantRNE_22U_11U_else_carry_2_sva);
  assign inp_lookup_2_FpMantRNE_22U_11U_else_acc_nl = nl_inp_lookup_2_FpMantRNE_22U_11U_else_acc_nl[9:0];
  assign or_5851_nl = FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp_1 | (~ inp_lookup_2_FpMantRNE_22U_11U_else_and_svs);
  assign mux_2026_nl = MUX_v_10_2_2((signext_10_1(~ FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp_1)),
      (inp_lookup_2_FpMantRNE_22U_11U_else_acc_nl), or_5851_nl);
  assign FpMul_6U_10U_nor_4_nl = ~(MUX_v_10_2_2((mux_2026_nl), 10'b1111111111, FpMul_6U_10U_is_inf_2_lpi_1_dfm_2));
  assign FpMul_6U_10U_FpMul_6U_10U_FpMul_6U_10U_nor_5_nl = ~(MUX_v_10_2_2((FpMul_6U_10U_nor_4_nl),
      10'b1111111111, FpMul_6U_10U_lor_10_lpi_1_dfm));
  assign FpMul_6U_10U_or_9_nl = FpMul_6U_10U_and_2_ssc | IsNaN_6U_10U_land_2_lpi_1_dfm_6;
  assign FpMul_6U_10U_o_mant_2_lpi_1_dfm_3_mx0w0 = MUX_v_10_2_2((FpMul_6U_10U_FpMul_6U_10U_FpMul_6U_10U_nor_5_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_23, FpMul_6U_10U_or_9_nl);
  assign FpMul_6U_10U_oelse_2_not_26_nl = ~ FpMul_6U_10U_lor_10_lpi_1_dfm;
  assign FpMul_6U_10U_FpMul_6U_10U_and_17_nl = MUX_v_4_2_2(4'b0000, (FpMul_6U_10U_o_expo_2_lpi_1_dfm[3:0]),
      (FpMul_6U_10U_oelse_2_not_26_nl));
  assign FpMul_6U_10U_o_expo_2_lpi_1_dfm_3_3_0_mx0w0 = MUX1HOT_v_4_3_2((FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_11_4_0_1[3:0]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_22, (FpMul_6U_10U_FpMul_6U_10U_and_17_nl),
      {IsNaN_6U_10U_land_2_lpi_1_dfm_6 , FpMul_6U_10U_and_2_ssc , FpMul_6U_10U_FpMul_6U_10U_nor_1_ssc});
  assign nl_FpAdd_6U_10U_is_a_greater_acc_1_nl = ({1'b1 , FpMul_6U_10U_o_expo_2_lpi_1_dfm_3_5_mx0w0
      , FpMul_6U_10U_o_expo_2_lpi_1_dfm_3_4_mx0w0 , FpMul_6U_10U_o_expo_2_lpi_1_dfm_3_3_0_mx0w0})
      + conv_u2u_6_7({(~ FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_14_1_1)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_14_0_1) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_26)})
      + 7'b1;
  assign FpAdd_6U_10U_is_a_greater_acc_1_nl = nl_FpAdd_6U_10U_is_a_greater_acc_1_nl[6:0];
  assign FpAdd_6U_10U_is_a_greater_acc_1_itm_6_1 = readslicef_7_1_6((FpAdd_6U_10U_is_a_greater_acc_1_nl));
  assign inp_lookup_3_FpAdd_6U_10U_is_a_greater_oif_equal_tmp = ({reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_15_tmp
      , reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_15_tmp_1 , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_27})
      == ({reg_FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_5_4_tmp , reg_FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_5_4_tmp_1
      , FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_3_0_1});
  assign nl_inp_lookup_3_FpMantRNE_22U_11U_else_acc_nl = (FpMul_6U_10U_p_mant_20_1_3_lpi_1_dfm_3_mx0[19:10])
      + conv_u2u_1_10(FpMantRNE_22U_11U_else_carry_3_sva);
  assign inp_lookup_3_FpMantRNE_22U_11U_else_acc_nl = nl_inp_lookup_3_FpMantRNE_22U_11U_else_acc_nl[9:0];
  assign or_5852_nl = FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp_2 | (~ inp_lookup_3_FpMantRNE_22U_11U_else_and_svs);
  assign mux_2027_nl = MUX_v_10_2_2((signext_10_1(~ FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp_2)),
      (inp_lookup_3_FpMantRNE_22U_11U_else_acc_nl), or_5852_nl);
  assign FpMul_6U_10U_nor_5_nl = ~(MUX_v_10_2_2((mux_2027_nl), 10'b1111111111, FpMul_6U_10U_is_inf_3_lpi_1_dfm_2));
  assign FpMul_6U_10U_FpMul_6U_10U_FpMul_6U_10U_nor_6_nl = ~(MUX_v_10_2_2((FpMul_6U_10U_nor_5_nl),
      10'b1111111111, FpMul_6U_10U_lor_11_lpi_1_dfm));
  assign FpMul_6U_10U_or_10_nl = FpMul_6U_10U_and_4_ssc | IsNaN_6U_10U_land_3_lpi_1_dfm_6;
  assign FpMul_6U_10U_o_mant_3_lpi_1_dfm_3_mx0w0 = MUX_v_10_2_2((FpMul_6U_10U_FpMul_6U_10U_FpMul_6U_10U_nor_6_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_22, FpMul_6U_10U_or_10_nl);
  assign FpMul_6U_10U_oelse_2_not_25_nl = ~ FpMul_6U_10U_lor_11_lpi_1_dfm;
  assign FpMul_6U_10U_FpMul_6U_10U_and_19_nl = MUX_v_4_2_2(4'b0000, (FpMul_6U_10U_o_expo_3_lpi_1_dfm[3:0]),
      (FpMul_6U_10U_oelse_2_not_25_nl));
  assign FpMul_6U_10U_o_expo_3_lpi_1_dfm_3_3_0_mx0w0 = MUX1HOT_v_4_3_2((FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_11_4_0_1[3:0]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_22, (FpMul_6U_10U_FpMul_6U_10U_and_19_nl),
      {IsNaN_6U_10U_land_3_lpi_1_dfm_6 , FpMul_6U_10U_and_4_ssc , FpMul_6U_10U_FpMul_6U_10U_nor_2_ssc});
  assign nl_FpAdd_6U_10U_is_a_greater_acc_2_nl = ({1'b1 , FpMul_6U_10U_o_expo_3_lpi_1_dfm_3_5_mx0w0
      , FpMul_6U_10U_o_expo_3_lpi_1_dfm_3_4_mx0w0 , FpMul_6U_10U_o_expo_3_lpi_1_dfm_3_3_0_mx0w0})
      + conv_u2u_6_7({(~ FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_14_1_1)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_14_0_1) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_26)})
      + 7'b1;
  assign FpAdd_6U_10U_is_a_greater_acc_2_nl = nl_FpAdd_6U_10U_is_a_greater_acc_2_nl[6:0];
  assign FpAdd_6U_10U_is_a_greater_acc_2_itm_6_1 = readslicef_7_1_6((FpAdd_6U_10U_is_a_greater_acc_2_nl));
  assign inp_lookup_4_FpAdd_6U_10U_is_a_greater_oif_equal_tmp = ({reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_15_tmp
      , reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_15_tmp_1 , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_27})
      == ({reg_FpMul_6U_10U_o_expo_lpi_1_dfm_6_5_4_tmp , reg_FpMul_6U_10U_o_expo_lpi_1_dfm_6_5_4_tmp_1
      , FpMul_6U_10U_o_expo_lpi_1_dfm_6_3_0_1});
  assign nl_inp_lookup_4_FpMantRNE_22U_11U_else_acc_nl = (FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0[19:10])
      + conv_u2u_1_10(FpMantRNE_22U_11U_else_carry_sva);
  assign inp_lookup_4_FpMantRNE_22U_11U_else_acc_nl = nl_inp_lookup_4_FpMantRNE_22U_11U_else_acc_nl[9:0];
  assign or_5853_nl = FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp_3 | (~ inp_lookup_4_FpMantRNE_22U_11U_else_and_svs);
  assign mux_2028_nl = MUX_v_10_2_2((signext_10_1(~ FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp_3)),
      (inp_lookup_4_FpMantRNE_22U_11U_else_acc_nl), or_5853_nl);
  assign FpMul_6U_10U_nor_6_nl = ~(MUX_v_10_2_2((mux_2028_nl), 10'b1111111111, FpMul_6U_10U_is_inf_lpi_1_dfm_2));
  assign FpMul_6U_10U_FpMul_6U_10U_FpMul_6U_10U_nor_7_nl = ~(MUX_v_10_2_2((FpMul_6U_10U_nor_6_nl),
      10'b1111111111, FpMul_6U_10U_lor_2_lpi_1_dfm));
  assign FpMul_6U_10U_or_11_nl = FpMul_6U_10U_and_6_ssc | IsNaN_6U_10U_land_lpi_1_dfm_6;
  assign FpMul_6U_10U_o_mant_lpi_1_dfm_3_mx0w0 = MUX_v_10_2_2((FpMul_6U_10U_FpMul_6U_10U_FpMul_6U_10U_nor_7_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_23, FpMul_6U_10U_or_11_nl);
  assign FpMul_6U_10U_oelse_2_not_24_nl = ~ FpMul_6U_10U_lor_2_lpi_1_dfm;
  assign FpMul_6U_10U_FpMul_6U_10U_and_21_nl = MUX_v_4_2_2(4'b0000, (FpMul_6U_10U_o_expo_lpi_1_dfm[3:0]),
      (FpMul_6U_10U_oelse_2_not_24_nl));
  assign FpMul_6U_10U_o_expo_lpi_1_dfm_3_3_0_mx0w0 = MUX1HOT_v_4_3_2((FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_11_4_0_1[3:0]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_22, (FpMul_6U_10U_FpMul_6U_10U_and_21_nl),
      {IsNaN_6U_10U_land_lpi_1_dfm_6 , FpMul_6U_10U_and_6_ssc , FpMul_6U_10U_FpMul_6U_10U_nor_3_ssc});
  assign nl_FpAdd_6U_10U_is_a_greater_acc_3_nl = ({1'b1 , FpMul_6U_10U_o_expo_lpi_1_dfm_3_5_mx0w0
      , FpMul_6U_10U_o_expo_lpi_1_dfm_3_4_mx0w0 , FpMul_6U_10U_o_expo_lpi_1_dfm_3_3_0_mx0w0})
      + conv_u2u_6_7({(~ FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_14_1_1)
      , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_14_0_1) , (~ FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_26)})
      + 7'b1;
  assign FpAdd_6U_10U_is_a_greater_acc_3_nl = nl_FpAdd_6U_10U_is_a_greater_acc_3_nl[6:0];
  assign FpAdd_6U_10U_is_a_greater_acc_3_itm_6_1 = readslicef_7_1_6((FpAdd_6U_10U_is_a_greater_acc_3_nl));
  assign FpAdd_6U_10U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0 = ((~ FpAdd_6U_10U_is_a_greater_oif_aelse_acc_itm_10_1)
      & inp_lookup_1_FpAdd_6U_10U_is_a_greater_oif_equal_tmp) | reg_inp_lookup_1_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse;
  assign FpAdd_6U_10U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0 = ((~ FpAdd_6U_10U_is_a_greater_oif_aelse_acc_1_itm_10_1)
      & inp_lookup_2_FpAdd_6U_10U_is_a_greater_oif_equal_tmp) | reg_inp_lookup_2_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse;
  assign FpAdd_6U_10U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0 = ((~ FpAdd_6U_10U_is_a_greater_oif_aelse_acc_2_itm_10_1)
      & inp_lookup_3_FpAdd_6U_10U_is_a_greater_oif_equal_tmp) | reg_inp_lookup_3_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse;
  assign FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_1_mx0w0 = ((~ FpAdd_6U_10U_is_a_greater_oif_aelse_acc_3_itm_10_1)
      & inp_lookup_4_FpAdd_6U_10U_is_a_greater_oif_equal_tmp) | reg_inp_lookup_4_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse;
  assign FpAdd_6U_10U_or_16_cse = IsNaN_6U_10U_3_land_1_lpi_1_dfm_8 | IsNaN_6U_10U_2_land_1_lpi_1_dfm_26;
  assign FpAdd_6U_10U_FpAdd_6U_10U_mux1h_13_nl = MUX1HOT_v_2_3_2(FpAdd_6U_10U_o_expo_1_lpi_1_dfm_2_5_4,
      (FpAdd_6U_10U_o_expo_1_sva_4[5:4]), ({reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_17_tmp
      , reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_17_tmp_1}), {FpAdd_6U_10U_and_ssc
      , FpAdd_6U_10U_and_6_ssc , FpAdd_6U_10U_or_16_cse});
  assign FpAdd_6U_10U_o_expo_1_lpi_1_dfm_7_5_4 = MUX_v_2_2_2((FpAdd_6U_10U_FpAdd_6U_10U_mux1h_13_nl),
      2'b11, FpAdd_6U_10U_and_28_ssc);
  assign IsInf_6U_23U_land_1_lpi_1_dfm_mx0w0 = ~((FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_22_13_1_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_9_0_1_lpi_1_dfm!=10'b0000000000)
      | IsNaN_6U_23U_IsNaN_6U_23U_nand_cse);
  assign IsInf_6U_23U_land_1_lpi_1_dfm_mx1 = MUX_s_1_2_2(IsInf_6U_23U_land_1_lpi_1_dfm_mx0w0,
      IsInf_6U_23U_land_1_lpi_1_dfm, or_dcpl_267);
  assign IsNaN_6U_23U_IsNaN_6U_23U_nor_tmp = ~((~((FpAdd_6U_10U_o_mant_1_lpi_1_dfm_2_mx0!=10'b0000000000)))
      | IsNaN_6U_23U_IsNaN_6U_23U_nand_cse);
  assign IsNaN_6U_23U_land_1_lpi_1_dfm_mx2 = MUX_s_1_2_2(IsNaN_6U_23U_IsNaN_6U_23U_nor_tmp,
      IsNaN_6U_23U_land_1_lpi_1_dfm, or_dcpl_267);
  assign nl_inp_lookup_1_FpAdd_6U_10U_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_3_5_4_tmp
      , reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_3_5_4_tmp_1 , (FpAdd_6U_10U_qr_2_lpi_1_dfm_3_3_0_1[3:1])})
      + 6'b1;
  assign inp_lookup_1_FpAdd_6U_10U_if_3_if_acc_1_nl = nl_inp_lookup_1_FpAdd_6U_10U_if_3_if_acc_1_nl[5:0];
  assign inp_lookup_1_FpAdd_6U_10U_if_3_if_acc_1_itm_5 = readslicef_6_1_5((inp_lookup_1_FpAdd_6U_10U_if_3_if_acc_1_nl));
  assign nl_FpAdd_6U_10U_asn_23_mx0w1 = ({1'b1 , (~ FpAdd_6U_10U_addend_smaller_qr_1_lpi_1_dfm_mx0)})
      + conv_u2u_23_24(FpAdd_6U_10U_addend_larger_qr_1_lpi_1_dfm_mx0) + 24'b1;
  assign FpAdd_6U_10U_asn_23_mx0w1 = nl_FpAdd_6U_10U_asn_23_mx0w1[23:0];
  assign nl_inp_lookup_1_FpNormalize_6U_23U_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_3_5_4_tmp)
      , (~ reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_3_5_4_tmp_1) , (~ FpAdd_6U_10U_qr_2_lpi_1_dfm_3_3_0_1)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_12)
      + 7'b1;
  assign inp_lookup_1_FpNormalize_6U_23U_acc_nl = nl_inp_lookup_1_FpNormalize_6U_23U_acc_nl[6:0];
  assign FpNormalize_6U_23U_if_FpNormalize_6U_23U_if_nand_tmp = ~(((FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_mx0[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((inp_lookup_1_FpNormalize_6U_23U_acc_nl))));
  assign FpAdd_6U_10U_or_17_cse = IsNaN_6U_10U_3_land_2_lpi_1_dfm_8 | IsNaN_6U_10U_2_land_2_lpi_1_dfm_26;
  assign FpAdd_6U_10U_FpAdd_6U_10U_mux1h_15_nl = MUX1HOT_v_2_3_2(FpAdd_6U_10U_o_expo_2_lpi_1_dfm_2_5_4,
      (FpAdd_6U_10U_o_expo_2_sva_4[5:4]), ({reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_17_tmp
      , reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_17_tmp_1}), {FpAdd_6U_10U_and_29_ssc
      , FpAdd_6U_10U_and_13_ssc , FpAdd_6U_10U_or_17_cse});
  assign FpAdd_6U_10U_o_expo_2_lpi_1_dfm_7_5_4 = MUX_v_2_2_2((FpAdd_6U_10U_FpAdd_6U_10U_mux1h_15_nl),
      2'b11, FpAdd_6U_10U_and_30_ssc);
  assign IsInf_6U_23U_land_2_lpi_1_dfm_mx0w0 = ~((FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_22_13_2_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_9_0_2_lpi_1_dfm!=10'b0000000000)
      | IsNaN_6U_23U_IsNaN_6U_23U_nand_1_cse);
  assign IsInf_6U_23U_land_2_lpi_1_dfm_mx1 = MUX_s_1_2_2(IsInf_6U_23U_land_2_lpi_1_dfm_mx0w0,
      IsInf_6U_23U_land_2_lpi_1_dfm, or_dcpl_269);
  assign IsNaN_6U_23U_IsNaN_6U_23U_nor_1_tmp = ~((~((FpAdd_6U_10U_o_mant_2_lpi_1_dfm_2_mx0!=10'b0000000000)))
      | IsNaN_6U_23U_IsNaN_6U_23U_nand_1_cse);
  assign IsNaN_6U_23U_land_2_lpi_1_dfm_mx2 = MUX_s_1_2_2(IsNaN_6U_23U_IsNaN_6U_23U_nor_1_tmp,
      IsNaN_6U_23U_land_2_lpi_1_dfm, or_dcpl_269);
  assign nl_inp_lookup_2_FpAdd_6U_10U_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_3_5_4_tmp
      , reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_3_5_4_tmp_1 , (FpAdd_6U_10U_qr_3_lpi_1_dfm_3_3_0_1[3:1])})
      + 6'b1;
  assign inp_lookup_2_FpAdd_6U_10U_if_3_if_acc_1_nl = nl_inp_lookup_2_FpAdd_6U_10U_if_3_if_acc_1_nl[5:0];
  assign inp_lookup_2_FpAdd_6U_10U_if_3_if_acc_1_itm_5 = readslicef_6_1_5((inp_lookup_2_FpAdd_6U_10U_if_3_if_acc_1_nl));
  assign nl_FpAdd_6U_10U_asn_20_mx0w1 = ({1'b1 , (~ FpAdd_6U_10U_addend_smaller_qr_2_lpi_1_dfm_mx0)})
      + conv_u2u_23_24(FpAdd_6U_10U_addend_larger_qr_2_lpi_1_dfm_mx0) + 24'b1;
  assign FpAdd_6U_10U_asn_20_mx0w1 = nl_FpAdd_6U_10U_asn_20_mx0w1[23:0];
  assign nl_inp_lookup_2_FpNormalize_6U_23U_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_3_5_4_tmp)
      , (~ reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_3_5_4_tmp_1) , (~ FpAdd_6U_10U_qr_3_lpi_1_dfm_3_3_0_1)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_13)
      + 7'b1;
  assign inp_lookup_2_FpNormalize_6U_23U_acc_nl = nl_inp_lookup_2_FpNormalize_6U_23U_acc_nl[6:0];
  assign FpNormalize_6U_23U_if_FpNormalize_6U_23U_if_nand_1_tmp = ~(((FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_mx0[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((inp_lookup_2_FpNormalize_6U_23U_acc_nl))));
  assign FpAdd_6U_10U_or_18_cse = IsNaN_6U_10U_3_land_3_lpi_1_dfm_8 | IsNaN_6U_10U_2_land_3_lpi_1_dfm_26;
  assign FpAdd_6U_10U_FpAdd_6U_10U_mux1h_17_nl = MUX1HOT_v_2_3_2(FpAdd_6U_10U_o_expo_3_lpi_1_dfm_2_5_4,
      (FpAdd_6U_10U_o_expo_3_sva_4[5:4]), ({reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_17_tmp
      , reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_17_tmp_1}), {FpAdd_6U_10U_and_31_ssc
      , FpAdd_6U_10U_and_19_ssc , FpAdd_6U_10U_or_18_cse});
  assign FpAdd_6U_10U_o_expo_3_lpi_1_dfm_7_5_4 = MUX_v_2_2_2((FpAdd_6U_10U_FpAdd_6U_10U_mux1h_17_nl),
      2'b11, FpAdd_6U_10U_and_32_ssc);
  assign IsInf_6U_23U_land_3_lpi_1_dfm_mx0w0 = ~((FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_22_13_3_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_9_0_3_lpi_1_dfm!=10'b0000000000)
      | IsNaN_6U_23U_IsNaN_6U_23U_nand_2_cse);
  assign IsInf_6U_23U_land_3_lpi_1_dfm_mx1 = MUX_s_1_2_2(IsInf_6U_23U_land_3_lpi_1_dfm_mx0w0,
      IsInf_6U_23U_land_3_lpi_1_dfm, or_dcpl_276);
  assign IsNaN_6U_23U_IsNaN_6U_23U_nor_2_tmp = ~((~((FpAdd_6U_10U_o_mant_3_lpi_1_dfm_2_mx0!=10'b0000000000)))
      | IsNaN_6U_23U_IsNaN_6U_23U_nand_2_cse);
  assign IsNaN_6U_23U_land_3_lpi_1_dfm_mx1 = MUX_s_1_2_2(IsNaN_6U_23U_IsNaN_6U_23U_nor_2_tmp,
      IsNaN_6U_23U_land_3_lpi_1_dfm, or_dcpl_276);
  assign nl_inp_lookup_3_FpAdd_6U_10U_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_3_5_4_tmp
      , reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_3_5_4_tmp_1 , (FpAdd_6U_10U_qr_4_lpi_1_dfm_3_3_0_1[3:1])})
      + 6'b1;
  assign inp_lookup_3_FpAdd_6U_10U_if_3_if_acc_1_nl = nl_inp_lookup_3_FpAdd_6U_10U_if_3_if_acc_1_nl[5:0];
  assign inp_lookup_3_FpAdd_6U_10U_if_3_if_acc_1_itm_5 = readslicef_6_1_5((inp_lookup_3_FpAdd_6U_10U_if_3_if_acc_1_nl));
  assign nl_FpAdd_6U_10U_asn_17_mx0w1 = ({1'b1 , (~ FpAdd_6U_10U_addend_smaller_qr_3_lpi_1_dfm_mx0)})
      + conv_u2u_23_24(FpAdd_6U_10U_addend_larger_qr_3_lpi_1_dfm_mx0) + 24'b1;
  assign FpAdd_6U_10U_asn_17_mx0w1 = nl_FpAdd_6U_10U_asn_17_mx0w1[23:0];
  assign nl_inp_lookup_3_FpNormalize_6U_23U_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_3_5_4_tmp)
      , (~ reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_3_5_4_tmp_1) , (~ FpAdd_6U_10U_qr_4_lpi_1_dfm_3_3_0_1)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_14)
      + 7'b1;
  assign inp_lookup_3_FpNormalize_6U_23U_acc_nl = nl_inp_lookup_3_FpNormalize_6U_23U_acc_nl[6:0];
  assign FpNormalize_6U_23U_if_FpNormalize_6U_23U_if_nand_2_tmp = ~(((FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_mx0[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((inp_lookup_3_FpNormalize_6U_23U_acc_nl))));
  assign FpAdd_6U_10U_or_19_cse = IsNaN_6U_10U_3_land_lpi_1_dfm_8 | IsNaN_6U_10U_2_land_lpi_1_dfm_26;
  assign FpAdd_6U_10U_FpAdd_6U_10U_mux1h_19_nl = MUX1HOT_v_2_3_2(FpAdd_6U_10U_o_expo_lpi_1_dfm_2_5_4,
      (FpAdd_6U_10U_o_expo_sva_4[5:4]), ({reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_17_tmp
      , reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_17_tmp_1}), {FpAdd_6U_10U_and_33_ssc
      , FpAdd_6U_10U_and_25_ssc , FpAdd_6U_10U_or_19_cse});
  assign FpAdd_6U_10U_o_expo_lpi_1_dfm_7_5_4 = MUX_v_2_2_2((FpAdd_6U_10U_FpAdd_6U_10U_mux1h_19_nl),
      2'b11, FpAdd_6U_10U_and_34_ssc);
  assign IsInf_6U_23U_land_lpi_1_dfm_mx0w0 = ~((FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_22_13_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_9_0_lpi_1_dfm!=10'b0000000000) |
      IsNaN_6U_23U_IsNaN_6U_23U_nand_3_cse);
  assign IsInf_6U_23U_land_lpi_1_dfm_mx1 = MUX_s_1_2_2(IsInf_6U_23U_land_lpi_1_dfm_mx0w0,
      IsInf_6U_23U_land_lpi_1_dfm, or_dcpl_278);
  assign IsNaN_6U_23U_IsNaN_6U_23U_nor_3_tmp = ~((~((FpAdd_6U_10U_o_mant_lpi_1_dfm_2_mx0!=10'b0000000000)))
      | IsNaN_6U_23U_IsNaN_6U_23U_nand_3_cse);
  assign IsNaN_6U_23U_land_lpi_1_dfm_mx1 = MUX_s_1_2_2(IsNaN_6U_23U_IsNaN_6U_23U_nor_3_tmp,
      IsNaN_6U_23U_land_lpi_1_dfm, or_dcpl_278);
  assign nl_inp_lookup_4_FpAdd_6U_10U_if_3_if_acc_1_nl = ({1'b1 , reg_FpAdd_6U_10U_qr_lpi_1_dfm_3_5_4_tmp
      , reg_FpAdd_6U_10U_qr_lpi_1_dfm_3_5_4_tmp_1 , (FpAdd_6U_10U_qr_lpi_1_dfm_3_3_0_1[3:1])})
      + 6'b1;
  assign inp_lookup_4_FpAdd_6U_10U_if_3_if_acc_1_nl = nl_inp_lookup_4_FpAdd_6U_10U_if_3_if_acc_1_nl[5:0];
  assign inp_lookup_4_FpAdd_6U_10U_if_3_if_acc_1_itm_5 = readslicef_6_1_5((inp_lookup_4_FpAdd_6U_10U_if_3_if_acc_1_nl));
  assign nl_FpAdd_6U_10U_asn_mx0w1 = ({1'b1 , (~ FpAdd_6U_10U_addend_smaller_qr_lpi_1_dfm_mx0)})
      + conv_u2u_23_24(FpAdd_6U_10U_addend_larger_qr_lpi_1_dfm_mx0) + 24'b1;
  assign FpAdd_6U_10U_asn_mx0w1 = nl_FpAdd_6U_10U_asn_mx0w1[23:0];
  assign nl_inp_lookup_4_FpNormalize_6U_23U_acc_nl = ({1'b1 , (~ reg_FpAdd_6U_10U_qr_lpi_1_dfm_3_5_4_tmp)
      , (~ reg_FpAdd_6U_10U_qr_lpi_1_dfm_3_5_4_tmp_1) , (~ FpAdd_6U_10U_qr_lpi_1_dfm_3_3_0_1)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_15)
      + 7'b1;
  assign inp_lookup_4_FpNormalize_6U_23U_acc_nl = nl_inp_lookup_4_FpNormalize_6U_23U_acc_nl[6:0];
  assign FpNormalize_6U_23U_if_FpNormalize_6U_23U_if_nand_3_tmp = ~(((FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_mx0[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((inp_lookup_4_FpNormalize_6U_23U_acc_nl))));
  assign IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_tmp = ~((FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_7_mx0w0==8'b11111111));
  assign IsNaN_8U_23U_4_nor_tmp = ~((FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_2_mx1!=23'b00000000000000000000000));
  assign FpMantRNE_24U_11U_else_carry_1_sva = (FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_2_mx1[12])
      & ((FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_2_mx1[0]) | (FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_2_mx1[1])
      | (FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_2_mx1[2]) | (FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_2_mx1[3])
      | (FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_2_mx1[4]) | (FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_2_mx1[5])
      | (FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_2_mx1[6]) | (FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_2_mx1[7])
      | (FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_2_mx1[8]) | (FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_2_mx1[9])
      | (FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_2_mx1[10]) | (FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_2_mx1[11])
      | (FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_2_mx1[13]));
  assign nl_inp_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_nl = FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_12
      + 8'b1;
  assign inp_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_nl = nl_inp_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_nl[7:0];
  assign FpAdd_8U_23U_1_or_nl = ((~(FpAdd_8U_23U_1_and_tmp | FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_2_mx0))
      & FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_5_m1c) | (IsNaN_8U_23U_3_land_1_lpi_1_dfm_7
      & (~ IsNaN_6U_10U_8_land_1_lpi_1_dfm_st_3));
  assign FpAdd_8U_23U_1_and_6_nl = FpAdd_8U_23U_1_and_tmp & (~ FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_2_mx0)
      & FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_5_m1c;
  assign FpAdd_8U_23U_1_and_28_nl = FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_2_mx0 & FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_5_m1c;
  assign FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_7_mx0w0 = MUX1HOT_v_8_4_2(FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_12,
      (inp_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_nl), 8'b11111110, reg_chn_inp_in_crt_sva_6_30_0_reg,
      {(FpAdd_8U_23U_1_or_nl) , (FpAdd_8U_23U_1_and_6_nl) , (FpAdd_8U_23U_1_and_28_nl)
      , IsNaN_6U_10U_8_land_1_lpi_1_dfm_st_3});
  assign or_6234_nl = IsNaN_8U_23U_3_land_1_lpi_1_dfm_7 | IsNaN_6U_10U_8_land_1_lpi_1_dfm_st_3;
  assign FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_2_mx1 = MUX_v_23_2_2(FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_4_itm,
      reg_chn_inp_in_crt_sva_6_30_0_1_reg, or_6234_nl);
  assign or_6233_nl = IsNaN_8U_23U_3_land_2_lpi_1_dfm_7 | IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_4;
  assign FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_2_mx1 = MUX_v_23_2_2(FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_5_itm,
      reg_chn_inp_in_crt_sva_6_62_32_1_reg, or_6233_nl);
  assign FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx1 = MUX_v_23_2_2(FpAdd_8U_23U_1_asn_40_mx0w1,
      reg_chn_inp_in_crt_sva_6_94_64_1_reg, IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_4);
  assign or_6232_nl = IsNaN_8U_23U_3_land_lpi_1_dfm_6 | IsNaN_6U_10U_8_land_lpi_1_dfm_st_4;
  assign FpAdd_8U_23U_1_o_mant_lpi_1_dfm_2_mx1 = MUX_v_23_2_2(FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_7_itm,
      reg_chn_inp_in_crt_sva_6_126_96_1_reg, or_6232_nl);
  assign nl_inp_lookup_1_FpMantRNE_22U_11U_2_else_acc_nl = inp_lookup_1_FpMantWidthDec_6U_21U_10U_0U_0U_1_overflow_slc_FpMantRNE_22U_11U_i_data_1_20_1_19_10_itm
      + conv_u2u_1_10(FpMantRNE_22U_11U_1_else_carry_1_sva_1);
  assign inp_lookup_1_FpMantRNE_22U_11U_2_else_acc_nl = nl_inp_lookup_1_FpMantRNE_22U_11U_2_else_acc_nl[9:0];
  assign or_5854_nl = FpMantWidthDec_6U_21U_10U_0U_0U_2_if_1_unequal_tmp | (~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_2);
  assign mux_2029_nl = MUX_v_10_2_2((signext_10_1(~ FpMantWidthDec_6U_21U_10U_0U_0U_2_if_1_unequal_tmp)),
      (inp_lookup_1_FpMantRNE_22U_11U_2_else_acc_nl), or_5854_nl);
  assign FpMul_6U_10U_2_nor_nl = ~(MUX_v_10_2_2((mux_2029_nl), 10'b1111111111, nor_1274_cse));
  assign FpMul_6U_10U_2_FpMul_6U_10U_2_FpMul_6U_10U_2_nor_4_nl = ~(MUX_v_10_2_2((FpMul_6U_10U_2_nor_nl),
      10'b1111111111, FpMul_6U_10U_2_lor_9_lpi_1_dfm));
  assign FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_3_mx0w0 = MUX_v_10_2_2((FpMul_6U_10U_2_FpMul_6U_10U_2_FpMul_6U_10U_2_nor_4_nl),
      ({reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_8_reg , reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_8_1_reg}),
      FpAdd_8U_23U_or_cse);
  assign nl_inp_lookup_2_FpMantRNE_22U_11U_2_else_acc_nl = FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_10
      + conv_u2u_1_10(FpMantRNE_22U_11U_1_else_carry_2_sva_1);
  assign inp_lookup_2_FpMantRNE_22U_11U_2_else_acc_nl = nl_inp_lookup_2_FpMantRNE_22U_11U_2_else_acc_nl[9:0];
  assign or_5855_nl = FpMantWidthDec_6U_21U_10U_0U_0U_2_if_1_unequal_tmp_1 | (~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_2);
  assign mux_2030_nl = MUX_v_10_2_2((signext_10_1(~ FpMantWidthDec_6U_21U_10U_0U_0U_2_if_1_unequal_tmp_1)),
      (inp_lookup_2_FpMantRNE_22U_11U_2_else_acc_nl), or_5855_nl);
  assign FpMul_6U_10U_2_nor_4_nl = ~(MUX_v_10_2_2((mux_2030_nl), 10'b1111111111,
      nor_1790_cse));
  assign FpMul_6U_10U_2_FpMul_6U_10U_2_FpMul_6U_10U_2_nor_5_itm = ~(MUX_v_10_2_2((FpMul_6U_10U_2_nor_4_nl),
      10'b1111111111, FpMul_6U_10U_2_lor_10_lpi_1_dfm));
  assign FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_3_mx0w0 = MUX_v_10_2_2(FpMul_6U_10U_2_FpMul_6U_10U_2_FpMul_6U_10U_2_nor_5_itm,
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_10, FpAdd_8U_23U_or_1_cse);
  assign nl_inp_lookup_4_FpMantRNE_22U_11U_2_else_acc_nl = inp_lookup_4_FpMantWidthDec_6U_21U_10U_0U_0U_1_overflow_slc_FpMantRNE_22U_11U_i_data_1_20_1_19_10_itm
      + conv_u2u_1_10(FpMantRNE_22U_11U_1_else_carry_sva);
  assign inp_lookup_4_FpMantRNE_22U_11U_2_else_acc_nl = nl_inp_lookup_4_FpMantRNE_22U_11U_2_else_acc_nl[9:0];
  assign or_5856_nl = FpMantWidthDec_6U_21U_10U_0U_0U_2_if_1_unequal_tmp_3 | (~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_sva_2);
  assign mux_2031_nl = MUX_v_10_2_2((signext_10_1(~ FpMantWidthDec_6U_21U_10U_0U_0U_2_if_1_unequal_tmp_3)),
      (inp_lookup_4_FpMantRNE_22U_11U_2_else_acc_nl), or_5856_nl);
  assign FpMul_6U_10U_2_nor_6_nl = ~(MUX_v_10_2_2((mux_2031_nl), 10'b1111111111,
      nor_1238_cse));
  assign FpMul_6U_10U_2_FpMul_6U_10U_2_FpMul_6U_10U_2_nor_7_nl = ~(MUX_v_10_2_2((FpMul_6U_10U_2_nor_6_nl),
      10'b1111111111, FpMul_6U_10U_2_lor_2_lpi_1_dfm));
  assign FpMul_6U_10U_2_o_mant_lpi_1_dfm_3_mx0w0 = MUX_v_10_2_2((FpMul_6U_10U_2_FpMul_6U_10U_2_FpMul_6U_10U_2_nor_7_nl),
      ({reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_8_reg , reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_8_1_reg}),
      FpAdd_8U_23U_or_3_cse);
  assign FpMantRNE_22U_11U_1_else_carry_1_sva = (FpMul_6U_10U_1_p_mant_20_1_1_lpi_1_dfm_3_mx0[9])
      & (((FpMul_6U_10U_1_p_mant_p1_1_sva_mx1_20_0[0]) & FpMul_6U_10U_1_p_mant_p1_1_sva_mx2_21)
      | (FpMul_6U_10U_1_p_mant_20_1_1_lpi_1_dfm_3_mx0[0]) | (FpMul_6U_10U_1_p_mant_20_1_1_lpi_1_dfm_3_mx0[1])
      | (FpMul_6U_10U_1_p_mant_20_1_1_lpi_1_dfm_3_mx0[2]) | (FpMul_6U_10U_1_p_mant_20_1_1_lpi_1_dfm_3_mx0[3])
      | (FpMul_6U_10U_1_p_mant_20_1_1_lpi_1_dfm_3_mx0[4]) | (FpMul_6U_10U_1_p_mant_20_1_1_lpi_1_dfm_3_mx0[5])
      | (FpMul_6U_10U_1_p_mant_20_1_1_lpi_1_dfm_3_mx0[6]) | (FpMul_6U_10U_1_p_mant_20_1_1_lpi_1_dfm_3_mx0[7])
      | (FpMul_6U_10U_1_p_mant_20_1_1_lpi_1_dfm_3_mx0[8]) | (FpMul_6U_10U_1_p_mant_20_1_1_lpi_1_dfm_3_mx0[10]));
  assign FpMantRNE_22U_11U_2_else_carry_1_sva_mx1w1 = (FpMul_6U_10U_2_p_mant_20_1_1_lpi_1_dfm_3_mx0[9])
      & (((FpMul_6U_10U_2_p_mant_p1_1_sva_mx1_20_0[0]) & FpMul_6U_10U_2_p_mant_p1_1_sva_mx2_21)
      | (FpMul_6U_10U_2_p_mant_20_1_1_lpi_1_dfm_3_mx0[0]) | (FpMul_6U_10U_2_p_mant_20_1_1_lpi_1_dfm_3_mx0[1])
      | (FpMul_6U_10U_2_p_mant_20_1_1_lpi_1_dfm_3_mx0[2]) | (FpMul_6U_10U_2_p_mant_20_1_1_lpi_1_dfm_3_mx0[3])
      | (FpMul_6U_10U_2_p_mant_20_1_1_lpi_1_dfm_3_mx0[4]) | (FpMul_6U_10U_2_p_mant_20_1_1_lpi_1_dfm_3_mx0[5])
      | (FpMul_6U_10U_2_p_mant_20_1_1_lpi_1_dfm_3_mx0[6]) | (FpMul_6U_10U_2_p_mant_20_1_1_lpi_1_dfm_3_mx0[7])
      | (FpMul_6U_10U_2_p_mant_20_1_1_lpi_1_dfm_3_mx0[8]) | (FpMul_6U_10U_2_p_mant_20_1_1_lpi_1_dfm_3_mx0[10]));
  assign inp_lookup_else_if_not_nl = ~ IsNaN_8U_23U_land_1_lpi_1_dfm_st_4;
  assign inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_3_4_0_mx0w0 = MUX_v_5_2_2(inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_4_0_1,
      5'b11111, (inp_lookup_else_if_not_nl));
  assign inp_lookup_else_if_not_1_nl = ~ IsNaN_8U_23U_land_2_lpi_1_dfm_st_4;
  assign inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_3_4_0_mx0w0 = MUX_v_5_2_2(inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_6_4_0_1,
      5'b11111, (inp_lookup_else_if_not_1_nl));
  assign FpMantRNE_22U_11U_1_else_carry_3_sva = (FpMul_6U_10U_1_p_mant_20_1_3_lpi_1_dfm_3_mx0[9])
      & (((FpMul_6U_10U_1_p_mant_p1_3_sva_mx1_20_0[0]) & FpMul_6U_10U_1_p_mant_p1_3_sva_mx2_21)
      | (FpMul_6U_10U_1_p_mant_20_1_3_lpi_1_dfm_3_mx0[0]) | (FpMul_6U_10U_1_p_mant_20_1_3_lpi_1_dfm_3_mx0[1])
      | (FpMul_6U_10U_1_p_mant_20_1_3_lpi_1_dfm_3_mx0[2]) | (FpMul_6U_10U_1_p_mant_20_1_3_lpi_1_dfm_3_mx0[3])
      | (FpMul_6U_10U_1_p_mant_20_1_3_lpi_1_dfm_3_mx0[4]) | (FpMul_6U_10U_1_p_mant_20_1_3_lpi_1_dfm_3_mx0[5])
      | (FpMul_6U_10U_1_p_mant_20_1_3_lpi_1_dfm_3_mx0[6]) | (FpMul_6U_10U_1_p_mant_20_1_3_lpi_1_dfm_3_mx0[7])
      | (FpMul_6U_10U_1_p_mant_20_1_3_lpi_1_dfm_3_mx0[8]) | (FpMul_6U_10U_1_p_mant_20_1_3_lpi_1_dfm_3_mx0[10]));
  assign FpMantRNE_22U_11U_2_else_carry_3_sva_mx1w1 = (FpMul_6U_10U_2_p_mant_20_1_3_lpi_1_dfm_3_mx0[9])
      & (((FpMul_6U_10U_2_p_mant_p1_3_sva_mx1_20_0[0]) & FpMul_6U_10U_2_p_mant_p1_3_sva_mx2_21)
      | (FpMul_6U_10U_2_p_mant_20_1_3_lpi_1_dfm_3_mx0[0]) | (FpMul_6U_10U_2_p_mant_20_1_3_lpi_1_dfm_3_mx0[1])
      | (FpMul_6U_10U_2_p_mant_20_1_3_lpi_1_dfm_3_mx0[2]) | (FpMul_6U_10U_2_p_mant_20_1_3_lpi_1_dfm_3_mx0[3])
      | (FpMul_6U_10U_2_p_mant_20_1_3_lpi_1_dfm_3_mx0[4]) | (FpMul_6U_10U_2_p_mant_20_1_3_lpi_1_dfm_3_mx0[5])
      | (FpMul_6U_10U_2_p_mant_20_1_3_lpi_1_dfm_3_mx0[6]) | (FpMul_6U_10U_2_p_mant_20_1_3_lpi_1_dfm_3_mx0[7])
      | (FpMul_6U_10U_2_p_mant_20_1_3_lpi_1_dfm_3_mx0[8]) | (FpMul_6U_10U_2_p_mant_20_1_3_lpi_1_dfm_3_mx0[10]));
  assign inp_lookup_else_if_not_2_nl = ~ IsNaN_8U_23U_land_3_lpi_1_dfm_st_4;
  assign inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_3_4_0_mx0w0 = MUX_v_5_2_2(inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_6_4_0_1,
      5'b11111, (inp_lookup_else_if_not_2_nl));
  assign inp_lookup_else_if_not_3_nl = ~ IsNaN_8U_23U_land_lpi_1_dfm_st_4;
  assign inp_lookup_else_if_a0_15_10_lpi_1_dfm_3_4_0_mx0w0 = MUX_v_5_2_2(inp_lookup_else_if_a0_15_10_lpi_1_dfm_6_4_0_1,
      5'b11111, (inp_lookup_else_if_not_3_nl));
  assign IsZero_5U_10U_3_aelse_not_23_nl = ~ IsZero_5U_10U_3_land_1_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_and_nl
      = MUX_v_10_2_2(10'b0000000000, (chn_inp_in_rsci_d_mxwt[341:332]), (IsZero_5U_10U_3_aelse_not_23_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_mux_4_nl = MUX_v_10_2_2(z_out_16, (FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_and_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_or_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_3_mux_4_nl), 10'b1111111111,
      IsInf_5U_10U_3_land_1_lpi_1_dfm);
  assign IsZero_5U_10U_3_aelse_not_22_nl = ~ IsZero_5U_10U_3_land_2_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_and_3_nl
      = MUX_v_10_2_2(10'b0000000000, (chn_inp_in_rsci_d_mxwt[357:348]), (IsZero_5U_10U_3_aelse_not_22_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_mux_36_nl = MUX_v_10_2_2(inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_itm,
      (FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_and_3_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_1_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_or_4_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_3_mux_36_nl), 10'b1111111111,
      IsInf_5U_10U_3_land_2_lpi_1_dfm);
  assign IsZero_5U_10U_3_aelse_not_21_nl = ~ IsZero_5U_10U_3_land_3_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_and_6_nl
      = MUX_v_10_2_2(10'b0000000000, (chn_inp_in_rsci_d_mxwt[373:364]), (IsZero_5U_10U_3_aelse_not_21_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_mux_37_nl = MUX_v_10_2_2(z_out_17, (FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_and_6_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_2_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_or_8_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_3_mux_37_nl), 10'b1111111111,
      IsInf_5U_10U_3_land_3_lpi_1_dfm);
  assign IsZero_5U_10U_3_aelse_not_20_nl = ~ IsZero_5U_10U_3_land_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_and_9_nl
      = MUX_v_10_2_2(10'b0000000000, (chn_inp_in_rsci_d_mxwt[389:380]), (IsZero_5U_10U_3_aelse_not_20_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_mux_38_nl = MUX_v_10_2_2(inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_lshift_itm,
      (FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_and_9_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_3_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_or_12_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_3_mux_38_nl), 10'b1111111111,
      IsInf_5U_10U_3_land_lpi_1_dfm);
  assign nl_FpMantRNE_36U_11U_1_else_ac_int_cctor_2_sva_mx0w0 = (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[35:25])
      + conv_u2u_1_11(FpMantRNE_36U_11U_1_else_carry_1_sva);
  assign FpMantRNE_36U_11U_1_else_ac_int_cctor_2_sva_mx0w0 = nl_FpMantRNE_36U_11U_1_else_ac_int_cctor_2_sva_mx0w0[10:0];
  assign nl_FpMantRNE_36U_11U_1_else_ac_int_cctor_3_sva_mx0w0 = (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[35:25])
      + conv_u2u_1_11(FpMantRNE_36U_11U_1_else_carry_2_sva);
  assign FpMantRNE_36U_11U_1_else_ac_int_cctor_3_sva_mx0w0 = nl_FpMantRNE_36U_11U_1_else_ac_int_cctor_3_sva_mx0w0[10:0];
  assign nl_FpMantRNE_36U_11U_1_else_ac_int_cctor_4_sva_mx0w0 = (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[35:25])
      + conv_u2u_1_11(FpMantRNE_36U_11U_1_else_carry_3_sva);
  assign FpMantRNE_36U_11U_1_else_ac_int_cctor_4_sva_mx0w0 = nl_FpMantRNE_36U_11U_1_else_ac_int_cctor_4_sva_mx0w0[10:0];
  assign nl_FpMantRNE_36U_11U_1_else_ac_int_cctor_sva_mx0w0 = (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[35:25])
      + conv_u2u_1_11(FpMantRNE_36U_11U_1_else_carry_sva);
  assign FpMantRNE_36U_11U_1_else_ac_int_cctor_sva_mx0w0 = nl_FpMantRNE_36U_11U_1_else_ac_int_cctor_sva_mx0w0[10:0];
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_4_nl
      = ~((chn_inp_in_rsci_d_mxwt[282]) | IsZero_5U_10U_2_land_1_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_18_nl = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_4_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_1_sva[4]), IsDenorm_5U_10U_2_land_1_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_3_0_mx0w0 = (FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_18_nl)
      | IsInf_5U_10U_1_land_1_lpi_1_dfm | IsNaN_5U_10U_1_land_1_lpi_1_dfm;
  assign IsZero_5U_10U_1_aelse_not_27_nl = ~ IsZero_5U_10U_2_land_1_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_16_nl
      = MUX_v_4_2_2(4'b0000, (chn_inp_in_rsci_d_mxwt[281:278]), (IsZero_5U_10U_1_aelse_not_27_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux1h_4_nl
      = MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_16_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_1_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_cse
      , IsDenorm_5U_10U_2_land_1_lpi_1_dfm , IsInf_5U_10U_1_land_1_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux1h_4_nl),
      4'b1111, IsNaN_5U_10U_1_land_1_lpi_1_dfm);
  assign inp_lookup_2_IsZero_6U_10U_5_IsZero_6U_10U_5_nor_mx0w1 = ~((chn_inp_in_rsci_d_mxwt[298])
      | FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_3_0_mx0w0 | (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_3_mx0w0!=4'b0000));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_6_nl
      = ~((chn_inp_in_rsci_d_mxwt[298]) | IsZero_5U_10U_2_land_2_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_20_nl = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_6_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_2_sva[4]), IsDenorm_5U_10U_2_land_2_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_3_0_mx0w0 = (FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_20_nl)
      | IsInf_5U_10U_1_land_2_lpi_1_dfm | IsNaN_5U_10U_1_land_2_lpi_1_dfm;
  assign IsZero_5U_10U_1_aelse_not_26_nl = ~ IsZero_5U_10U_2_land_2_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_18_nl
      = MUX_v_4_2_2(4'b0000, (chn_inp_in_rsci_d_mxwt[297:294]), (IsZero_5U_10U_1_aelse_not_26_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux1h_6_nl
      = MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_18_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_2_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_1_cse
      , IsDenorm_5U_10U_2_land_2_lpi_1_dfm , IsInf_5U_10U_1_land_2_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux1h_6_nl),
      4'b1111, IsNaN_5U_10U_1_land_2_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_8_nl
      = ~((chn_inp_in_rsci_d_mxwt[314]) | IsZero_5U_10U_2_land_3_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_22_nl = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_8_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_3_sva[4]), IsDenorm_5U_10U_2_land_3_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_3_0_mx0w0 = (FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_22_nl)
      | IsInf_5U_10U_1_land_3_lpi_1_dfm | IsNaN_5U_10U_1_land_3_lpi_1_dfm;
  assign IsZero_5U_10U_1_aelse_not_25_nl = ~ IsZero_5U_10U_2_land_3_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_20_nl
      = MUX_v_4_2_2(4'b0000, (chn_inp_in_rsci_d_mxwt[313:310]), (IsZero_5U_10U_1_aelse_not_25_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux1h_8_nl
      = MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_20_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_3_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_2_cse
      , IsDenorm_5U_10U_2_land_3_lpi_1_dfm , IsInf_5U_10U_1_land_3_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux1h_8_nl),
      4'b1111, IsNaN_5U_10U_1_land_3_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_10_nl
      = ~((chn_inp_in_rsci_d_mxwt[330]) | IsZero_5U_10U_2_land_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_24_nl = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_nor_10_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_sva[4]), IsDenorm_5U_10U_2_land_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_3_0_mx0w0 = (FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_mux_24_nl)
      | IsInf_5U_10U_1_land_lpi_1_dfm | IsNaN_5U_10U_1_land_lpi_1_dfm;
  assign inp_lookup_4_IsZero_6U_10U_5_IsZero_6U_10U_5_nor_mx0w1 = ~((chn_inp_in_rsci_d_mxwt[330])
      | FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_3_0_mx0w0 | (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_3_mx0w0!=4'b0000));
  assign IsZero_5U_10U_1_aelse_not_24_nl = ~ IsZero_5U_10U_2_land_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_22_nl
      = MUX_v_4_2_2(4'b0000, (chn_inp_in_rsci_d_mxwt[329:326]), (IsZero_5U_10U_1_aelse_not_24_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux1h_10_nl
      = MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_and_22_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_3_cse
      , IsDenorm_5U_10U_2_land_lpi_1_dfm , IsInf_5U_10U_1_land_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux1h_10_nl),
      4'b1111, IsNaN_5U_10U_1_land_lpi_1_dfm);
  assign FpMul_6U_10U_2_p_mant_p1_1_sva_mx1_20_0 = MUX_v_21_2_2((FpMul_6U_10U_2_p_mant_p1_1_sva_mx3[20:0]),
      (FpMul_6U_10U_2_p_mant_p1_1_sva[20:0]), FpMul_6U_10U_2_lor_6_lpi_1_dfm_st_3);
  assign FpMul_6U_10U_2_p_mant_p1_1_sva_mx2_21 = MUX_s_1_2_2((FpMul_6U_10U_2_p_mant_p1_1_sva_mx3[21]),
      (FpMul_6U_10U_2_p_mant_p1_1_sva[21]), FpMul_6U_10U_2_lor_6_lpi_1_dfm_st_3);
  assign inp_lookup_1_FpMul_6U_10U_2_p_mant_p1_mul_tmp = conv_u2u_22_22(({1'b1 ,
      FpFractionToFloat_35U_6U_10U_1_o_mant_1_lpi_1_dfm_8}) * ({1'b1 , reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_7_itm
      , reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_7_1_itm}));
  assign FpMul_6U_10U_2_p_mant_p1_1_sva_mx3 = MUX_v_22_2_2(FpMul_6U_10U_2_p_mant_p1_1_sva,
      inp_lookup_1_FpMul_6U_10U_2_p_mant_p1_mul_tmp, inp_lookup_1_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs);
  assign FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_3_5_mx0w0 = (IntLeadZero_35U_1_leading_sign_35_0_rtn_1_sva_2[5])
      & (~(FpFractionToFloat_35U_6U_10U_1_if_else_else_if_slc_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_5_mdf_1_sva_2
      & (~ inp_lookup_1_FpMantRNE_36U_11U_1_else_and_svs_2) & FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_st_2))
      & (~ FpFractionToFloat_35U_6U_10U_1_is_zero_1_lpi_1_dfm_1);
  assign nl_inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_else_else_else_acc_nl
      = (~ (IntLeadZero_35U_1_leading_sign_35_0_rtn_1_sva_2[4:0])) + 5'b11111;
  assign inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_else_else_else_acc_nl = nl_inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_else_else_else_acc_nl[4:0];
  assign FpFractionToFloat_35U_6U_10U_1_and_nl = inp_lookup_1_FpMantRNE_36U_11U_1_else_and_svs_2
      & FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_st_2;
  assign FpFractionToFloat_35U_6U_10U_1_mux_tmp = MUX_v_5_2_2((inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_else_else_else_acc_nl),
      (~ (IntLeadZero_35U_1_leading_sign_35_0_rtn_1_sva_2[4:0])), FpFractionToFloat_35U_6U_10U_1_and_nl);
  assign FpFractionToFloat_35U_6U_10U_1_nor_4_nl = ~(MUX_v_5_2_2(FpFractionToFloat_35U_6U_10U_1_mux_tmp,
      5'b11111, FpFractionToFloat_35U_6U_10U_1_is_zero_1_lpi_1_dfm_1));
  assign FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_3_4_0_mx0w0 = ~(MUX_v_5_2_2((FpFractionToFloat_35U_6U_10U_1_nor_4_nl),
      5'b11111, FpFractionToFloat_35U_6U_10U_1_is_zero_1_lpi_1_dfm_1));
  assign FpMul_6U_10U_2_p_mant_p1_2_sva_mx1_20_0 = MUX_v_21_2_2((FpMul_6U_10U_2_p_mant_p1_2_sva_mx3[20:0]),
      (FpMul_6U_10U_2_p_mant_p1_2_sva[20:0]), FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_3);
  assign FpMul_6U_10U_2_p_mant_p1_2_sva_mx2_21 = MUX_s_1_2_2((FpMul_6U_10U_2_p_mant_p1_2_sva_mx3[21]),
      (FpMul_6U_10U_2_p_mant_p1_2_sva[21]), FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_3);
  assign inp_lookup_2_FpMul_6U_10U_2_p_mant_p1_mul_tmp = conv_u2u_22_22(({1'b1 ,
      FpFractionToFloat_35U_6U_10U_1_o_mant_2_lpi_1_dfm_8}) * ({1'b1 , reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_7_itm
      , reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_7_1_itm}));
  assign FpMul_6U_10U_2_p_mant_p1_2_sva_mx3 = MUX_v_22_2_2(FpMul_6U_10U_2_p_mant_p1_2_sva,
      inp_lookup_2_FpMul_6U_10U_2_p_mant_p1_mul_tmp, inp_lookup_2_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs);
  assign FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_3_5_mx0w0 = (IntLeadZero_35U_1_leading_sign_35_0_rtn_2_sva_2[5])
      & (~(FpFractionToFloat_35U_6U_10U_1_if_else_else_if_slc_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_5_mdf_2_sva_2
      & (~ inp_lookup_2_FpMantRNE_36U_11U_1_else_and_svs_2) & FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_st_2))
      & (~ FpFractionToFloat_35U_6U_10U_1_is_zero_2_lpi_1_dfm_1);
  assign FpFractionToFloat_35U_6U_10U_1_and_1_cse = inp_lookup_2_FpMantRNE_36U_11U_1_else_and_svs_2
      & FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_st_2;
  assign nl_inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_else_else_else_acc_nl
      = (~ (IntLeadZero_35U_1_leading_sign_35_0_rtn_2_sva_2[4:0])) + 5'b11111;
  assign inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_else_else_else_acc_nl = nl_inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_else_else_else_acc_nl[4:0];
  assign FpFractionToFloat_35U_6U_10U_1_mux_40_tmp = MUX_v_5_2_2((inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_else_else_else_acc_nl),
      (~ (IntLeadZero_35U_1_leading_sign_35_0_rtn_2_sva_2[4:0])), FpFractionToFloat_35U_6U_10U_1_and_1_cse);
  assign FpFractionToFloat_35U_6U_10U_1_nor_nl = ~(MUX_v_5_2_2(FpFractionToFloat_35U_6U_10U_1_mux_40_tmp,
      5'b11111, FpFractionToFloat_35U_6U_10U_1_is_zero_2_lpi_1_dfm_1));
  assign FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_3_4_0_mx0w0 = ~(MUX_v_5_2_2((FpFractionToFloat_35U_6U_10U_1_nor_nl),
      5'b11111, FpFractionToFloat_35U_6U_10U_1_is_zero_2_lpi_1_dfm_1));
  assign FpMul_6U_10U_2_p_mant_p1_3_sva_mx1_20_0 = MUX_v_21_2_2((FpMul_6U_10U_2_p_mant_p1_3_sva_mx3[20:0]),
      (FpMul_6U_10U_2_p_mant_p1_3_sva[20:0]), FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_3);
  assign FpMul_6U_10U_2_p_mant_p1_3_sva_mx2_21 = MUX_s_1_2_2((FpMul_6U_10U_2_p_mant_p1_3_sva_mx3[21]),
      (FpMul_6U_10U_2_p_mant_p1_3_sva[21]), FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_3);
  assign inp_lookup_3_FpMul_6U_10U_2_p_mant_p1_mul_tmp = conv_u2u_22_22(({1'b1 ,
      FpFractionToFloat_35U_6U_10U_1_o_mant_3_lpi_1_dfm_8}) * ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_3_lpi_1_dfm_9}));
  assign FpMul_6U_10U_2_p_mant_p1_3_sva_mx3 = MUX_v_22_2_2(FpMul_6U_10U_2_p_mant_p1_3_sva,
      inp_lookup_3_FpMul_6U_10U_2_p_mant_p1_mul_tmp, inp_lookup_3_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs);
  assign FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_3_5_mx0w0 = (IntLeadZero_35U_1_leading_sign_35_0_rtn_3_sva_2[5])
      & (~(FpFractionToFloat_35U_6U_10U_1_if_else_else_if_slc_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_5_mdf_3_sva_2
      & (~ inp_lookup_3_FpMantRNE_36U_11U_1_else_and_svs_2) & FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_st_2))
      & (~ FpFractionToFloat_35U_6U_10U_1_is_zero_3_lpi_1_dfm_1);
  assign FpFractionToFloat_35U_6U_10U_1_and_2_cse = inp_lookup_3_FpMantRNE_36U_11U_1_else_and_svs_2
      & FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_st_2;
  assign nl_inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_else_else_else_acc_nl
      = (~ (IntLeadZero_35U_1_leading_sign_35_0_rtn_3_sva_2[4:0])) + 5'b11111;
  assign inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_else_else_else_acc_nl = nl_inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_else_else_else_acc_nl[4:0];
  assign FpFractionToFloat_35U_6U_10U_1_mux_41_tmp = MUX_v_5_2_2((inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_else_else_else_acc_nl),
      (~ (IntLeadZero_35U_1_leading_sign_35_0_rtn_3_sva_2[4:0])), FpFractionToFloat_35U_6U_10U_1_and_2_cse);
  assign FpFractionToFloat_35U_6U_10U_1_nor_5_nl = ~(MUX_v_5_2_2(FpFractionToFloat_35U_6U_10U_1_mux_41_tmp,
      5'b11111, FpFractionToFloat_35U_6U_10U_1_is_zero_3_lpi_1_dfm_1));
  assign FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_3_4_0_mx0w0 = ~(MUX_v_5_2_2((FpFractionToFloat_35U_6U_10U_1_nor_5_nl),
      5'b11111, FpFractionToFloat_35U_6U_10U_1_is_zero_3_lpi_1_dfm_1));
  assign FpMul_6U_10U_2_p_mant_p1_sva_mx1_20_0 = MUX_v_21_2_2((FpMul_6U_10U_2_p_mant_p1_sva_mx3[20:0]),
      (FpMul_6U_10U_2_p_mant_p1_sva[20:0]), FpMul_6U_10U_2_lor_1_lpi_1_dfm_st_3);
  assign FpMul_6U_10U_2_p_mant_p1_sva_mx2_21 = MUX_s_1_2_2((FpMul_6U_10U_2_p_mant_p1_sva_mx3[21]),
      (FpMul_6U_10U_2_p_mant_p1_sva[21]), FpMul_6U_10U_2_lor_1_lpi_1_dfm_st_3);
  assign inp_lookup_4_FpMul_6U_10U_2_p_mant_p1_mul_tmp = conv_u2u_22_22(({1'b1 ,
      FpFractionToFloat_35U_6U_10U_1_o_mant_lpi_1_dfm_8}) * ({1'b1 , reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_7_itm
      , reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_7_1_itm}));
  assign FpMul_6U_10U_2_p_mant_p1_sva_mx3 = MUX_v_22_2_2(FpMul_6U_10U_2_p_mant_p1_sva,
      inp_lookup_4_FpMul_6U_10U_2_p_mant_p1_mul_tmp, inp_lookup_4_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs);
  assign FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_3_5_mx0w0 = (IntLeadZero_35U_1_leading_sign_35_0_rtn_sva_2[5])
      & (~(FpFractionToFloat_35U_6U_10U_1_if_else_else_if_slc_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_5_mdf_sva_2
      & (~ inp_lookup_4_FpMantRNE_36U_11U_1_else_and_svs_2) & FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2))
      & (~ FpFractionToFloat_35U_6U_10U_1_is_zero_lpi_1_dfm_1);
  assign nl_inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_else_else_else_acc_nl
      = (~ (IntLeadZero_35U_1_leading_sign_35_0_rtn_sva_2[4:0])) + 5'b11111;
  assign inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_else_else_else_acc_nl = nl_inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_else_else_else_acc_nl[4:0];
  assign FpFractionToFloat_35U_6U_10U_1_and_3_nl = inp_lookup_4_FpMantRNE_36U_11U_1_else_and_svs_2
      & FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2;
  assign FpFractionToFloat_35U_6U_10U_1_mux_42_tmp = MUX_v_5_2_2((inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_else_else_else_acc_nl),
      (~ (IntLeadZero_35U_1_leading_sign_35_0_rtn_sva_2[4:0])), FpFractionToFloat_35U_6U_10U_1_and_3_nl);
  assign FpFractionToFloat_35U_6U_10U_1_nor_6_nl = ~(MUX_v_5_2_2(FpFractionToFloat_35U_6U_10U_1_mux_42_tmp,
      5'b11111, FpFractionToFloat_35U_6U_10U_1_is_zero_lpi_1_dfm_1));
  assign FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_3_4_0_mx0w0 = ~(MUX_v_5_2_2((FpFractionToFloat_35U_6U_10U_1_nor_6_nl),
      5'b11111, FpFractionToFloat_35U_6U_10U_1_is_zero_lpi_1_dfm_1));
  assign nl_inp_lookup_1_FpNormalize_8U_49U_acc_nl = ({1'b1 , (~ reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_7_1_itm)})
      + conv_u2s_6_9(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_8)
      + 9'b1;
  assign inp_lookup_1_FpNormalize_8U_49U_acc_nl = nl_inp_lookup_1_FpNormalize_8U_49U_acc_nl[8:0];
  assign FpNormalize_8U_49U_if_FpNormalize_8U_49U_if_nand_tmp = ~(((z_out[48:0]!=49'b0000000000000000000000000000000000000000000000000))
      & (readslicef_9_1_8((inp_lookup_1_FpNormalize_8U_49U_acc_nl))));
  assign inp_lookup_1_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_tmp
      = (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_19!=10'b0000000000);
  assign nl_inp_lookup_2_FpNormalize_8U_49U_acc_nl = ({1'b1 , (~ reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_7_1_itm)})
      + conv_u2s_6_9(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_9)
      + 9'b1;
  assign inp_lookup_2_FpNormalize_8U_49U_acc_nl = nl_inp_lookup_2_FpNormalize_8U_49U_acc_nl[8:0];
  assign FpNormalize_8U_49U_if_FpNormalize_8U_49U_if_nand_1_tmp = ~(((z_out_1[48:0]!=49'b0000000000000000000000000000000000000000000000000))
      & (readslicef_9_1_8((inp_lookup_2_FpNormalize_8U_49U_acc_nl))));
  assign inp_lookup_2_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_tmp
      = (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_19!=10'b0000000000);
  assign nl_inp_lookup_3_FpNormalize_8U_49U_acc_nl = ({1'b1 , (~ reg_FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_7_1_itm)})
      + conv_u2s_6_9(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_10)
      + 9'b1;
  assign inp_lookup_3_FpNormalize_8U_49U_acc_nl = nl_inp_lookup_3_FpNormalize_8U_49U_acc_nl[8:0];
  assign FpNormalize_8U_49U_if_FpNormalize_8U_49U_if_nand_2_tmp = ~(((z_out_2[48:0]!=49'b0000000000000000000000000000000000000000000000000))
      & (readslicef_9_1_8((inp_lookup_3_FpNormalize_8U_49U_acc_nl))));
  assign inp_lookup_3_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_tmp
      = (reg_FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_7_itm!=2'b00) |
      (reg_FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_7_1_itm!=8'b00000000);
  assign nl_inp_lookup_4_FpNormalize_8U_49U_acc_nl = ({1'b1 , (~ reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_7_1_itm)})
      + conv_u2s_6_9(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_11)
      + 9'b1;
  assign inp_lookup_4_FpNormalize_8U_49U_acc_nl = nl_inp_lookup_4_FpNormalize_8U_49U_acc_nl[8:0];
  assign FpNormalize_8U_49U_if_FpNormalize_8U_49U_if_nand_3_tmp = ~(((z_out_3[48:0]!=49'b0000000000000000000000000000000000000000000000000))
      & (readslicef_9_1_8((inp_lookup_4_FpNormalize_8U_49U_acc_nl))));
  assign inp_lookup_4_IsNaN_6U_10U_5_aif_IsNaN_6U_10U_5_aelse_IsNaN_6U_10U_5_aelse_or_tmp
      = (FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_19!=10'b0000000000);
  assign inp_lookup_1_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp = (chn_inp_in_crt_sva_3_127_0_1[30:23])
      == FpAdd_8U_23U_o_expo_1_lpi_1_dfm_7_mx1w1;
  assign FpMul_6U_10U_1_p_mant_p1_1_sva_mx1_20_0 = MUX_v_21_2_2((FpMul_6U_10U_1_p_mant_p1_1_sva_mx3[20:0]),
      (FpMul_6U_10U_1_p_mant_p1_1_sva[20:0]), FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_3);
  assign FpMul_6U_10U_1_p_mant_p1_1_sva_mx2_21 = MUX_s_1_2_2((FpMul_6U_10U_1_p_mant_p1_1_sva_mx3[21]),
      (FpMul_6U_10U_1_p_mant_p1_1_sva[21]), FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_3);
  assign inp_lookup_1_FpMul_6U_10U_1_p_mant_p1_mul_tmp = conv_u2u_22_22(({1'b1 ,
      inp_lookup_else_if_a0_9_0_1_lpi_1_dfm_10}) * ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_20}));
  assign FpMul_6U_10U_1_p_mant_p1_1_sva_mx3 = MUX_v_22_2_2(FpMul_6U_10U_1_p_mant_p1_1_sva,
      inp_lookup_1_FpMul_6U_10U_1_p_mant_p1_mul_tmp, inp_lookup_1_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs);
  assign nl_FpMul_6U_10U_2_else_2_else_acc_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_7_1_1
      , FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_7_0_1 , FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_10})
      + 6'b100001;
  assign FpMul_6U_10U_2_else_2_else_acc_nl = nl_FpMul_6U_10U_2_else_2_else_acc_nl[5:0];
  assign nl_FpMul_6U_10U_2_else_2_else_ac_int_cctor_1_sva_mx0w0 = (FpMul_6U_10U_2_else_2_else_acc_nl)
      + ({FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_6_5_1 , FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_6_4_0_1});
  assign FpMul_6U_10U_2_else_2_else_ac_int_cctor_1_sva_mx0w0 = nl_FpMul_6U_10U_2_else_2_else_ac_int_cctor_1_sva_mx0w0[5:0];
  assign inp_lookup_2_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp = (chn_inp_in_crt_sva_3_127_0_1[62:55])
      == FpAdd_8U_23U_o_expo_2_lpi_1_dfm_7_mx1w1;
  assign FpMul_6U_10U_1_p_mant_p1_2_sva_mx1_20_0 = MUX_v_21_2_2((FpMul_6U_10U_1_p_mant_p1_2_sva_mx3[20:0]),
      (FpMul_6U_10U_1_p_mant_p1_2_sva[20:0]), FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_3);
  assign FpMul_6U_10U_1_p_mant_p1_2_sva_mx2_21 = MUX_s_1_2_2((FpMul_6U_10U_1_p_mant_p1_2_sva_mx3[21]),
      (FpMul_6U_10U_1_p_mant_p1_2_sva[21]), FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_3);
  assign inp_lookup_2_FpMul_6U_10U_1_p_mant_p1_mul_tmp = conv_u2u_22_22(({1'b1 ,
      inp_lookup_else_if_a0_9_0_2_lpi_1_dfm_10}) * ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_20}));
  assign FpMul_6U_10U_1_p_mant_p1_2_sva_mx3 = MUX_v_22_2_2(FpMul_6U_10U_1_p_mant_p1_2_sva,
      inp_lookup_2_FpMul_6U_10U_1_p_mant_p1_mul_tmp, inp_lookup_2_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs);
  assign nl_FpMul_6U_10U_2_else_2_else_acc_2_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_7_1_1
      , FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_7_0_1 , FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_10})
      + 6'b100001;
  assign FpMul_6U_10U_2_else_2_else_acc_2_nl = nl_FpMul_6U_10U_2_else_2_else_acc_2_nl[5:0];
  assign nl_FpMul_6U_10U_2_else_2_else_ac_int_cctor_2_sva_mx0w0 = (FpMul_6U_10U_2_else_2_else_acc_2_nl)
      + ({FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_6_5_1 , FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_6_4_0_1});
  assign FpMul_6U_10U_2_else_2_else_ac_int_cctor_2_sva_mx0w0 = nl_FpMul_6U_10U_2_else_2_else_ac_int_cctor_2_sva_mx0w0[5:0];
  assign inp_lookup_3_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp = (chn_inp_in_crt_sva_3_127_0_1[94:87])
      == FpAdd_8U_23U_o_expo_3_lpi_1_dfm_7_mx1w1;
  assign FpMul_6U_10U_1_p_mant_p1_3_sva_mx1_20_0 = MUX_v_21_2_2((FpMul_6U_10U_1_p_mant_p1_3_sva_mx3[20:0]),
      (FpMul_6U_10U_1_p_mant_p1_3_sva[20:0]), FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_3);
  assign FpMul_6U_10U_1_p_mant_p1_3_sva_mx2_21 = MUX_s_1_2_2((FpMul_6U_10U_1_p_mant_p1_3_sva_mx3[21]),
      (FpMul_6U_10U_1_p_mant_p1_3_sva[21]), FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_3);
  assign inp_lookup_3_FpMul_6U_10U_1_p_mant_p1_mul_tmp = conv_u2u_22_22(({1'b1 ,
      inp_lookup_else_if_a0_9_0_3_lpi_1_dfm_10}) * ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_10}));
  assign FpMul_6U_10U_1_p_mant_p1_3_sva_mx3 = MUX_v_22_2_2(FpMul_6U_10U_1_p_mant_p1_3_sva,
      inp_lookup_3_FpMul_6U_10U_1_p_mant_p1_mul_tmp, inp_lookup_3_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs);
  assign nl_FpMul_6U_10U_2_else_2_else_acc_3_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_7_1_1
      , FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_7_0_1 , FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_3_lpi_1_dfm_10})
      + 6'b100001;
  assign FpMul_6U_10U_2_else_2_else_acc_3_nl = nl_FpMul_6U_10U_2_else_2_else_acc_3_nl[5:0];
  assign nl_FpMul_6U_10U_2_else_2_else_ac_int_cctor_3_sva_mx0w0 = (FpMul_6U_10U_2_else_2_else_acc_3_nl)
      + ({FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_6_5_1 , FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_6_4_0_1});
  assign FpMul_6U_10U_2_else_2_else_ac_int_cctor_3_sva_mx0w0 = nl_FpMul_6U_10U_2_else_2_else_ac_int_cctor_3_sva_mx0w0[5:0];
  assign inp_lookup_4_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp = (chn_inp_in_crt_sva_3_127_0_1[126:119])
      == FpAdd_8U_23U_o_expo_lpi_1_dfm_7_mx1w1;
  assign FpMul_6U_10U_1_p_mant_p1_sva_mx1_20_0 = MUX_v_21_2_2((FpMul_6U_10U_1_p_mant_p1_sva_mx3[20:0]),
      (FpMul_6U_10U_1_p_mant_p1_sva[20:0]), FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_3);
  assign FpMul_6U_10U_1_p_mant_p1_sva_mx2_21 = MUX_s_1_2_2((FpMul_6U_10U_1_p_mant_p1_sva_mx3[21]),
      (FpMul_6U_10U_1_p_mant_p1_sva[21]), FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_3);
  assign inp_lookup_4_FpMul_6U_10U_1_p_mant_p1_mul_tmp = conv_u2u_22_22(({1'b1 ,
      inp_lookup_else_if_a0_9_0_lpi_1_dfm_10}) * ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_20}));
  assign FpMul_6U_10U_1_p_mant_p1_sva_mx3 = MUX_v_22_2_2(FpMul_6U_10U_1_p_mant_p1_sva,
      inp_lookup_4_FpMul_6U_10U_1_p_mant_p1_mul_tmp, inp_lookup_4_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs);
  assign nl_FpMul_6U_10U_2_else_2_else_acc_4_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_7_1_1
      , FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_7_0_1 , FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_10})
      + 6'b100001;
  assign FpMul_6U_10U_2_else_2_else_acc_4_nl = nl_FpMul_6U_10U_2_else_2_else_acc_4_nl[5:0];
  assign nl_FpMul_6U_10U_2_else_2_else_ac_int_cctor_sva_mx0w0 = (FpMul_6U_10U_2_else_2_else_acc_4_nl)
      + ({FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_6_5_1 , FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_6_4_0_1});
  assign FpMul_6U_10U_2_else_2_else_ac_int_cctor_sva_mx0w0 = nl_FpMul_6U_10U_2_else_2_else_ac_int_cctor_sva_mx0w0[5:0];
  assign nl_inp_lookup_1_FpMantRNE_49U_24U_else_acc_nl = (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[47:25])
      + conv_u2u_1_23(FpMantRNE_49U_24U_else_carry_1_sva);
  assign inp_lookup_1_FpMantRNE_49U_24U_else_acc_nl = nl_inp_lookup_1_FpMantRNE_49U_24U_else_acc_nl[22:0];
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_4_itm = MUX_v_23_2_2((inp_lookup_1_FpMantRNE_49U_24U_else_acc_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0);
  assign nl_inp_lookup_2_FpMantRNE_49U_24U_else_acc_nl = (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[47:25])
      + conv_u2u_1_23(FpMantRNE_49U_24U_else_carry_2_sva);
  assign inp_lookup_2_FpMantRNE_49U_24U_else_acc_nl = nl_inp_lookup_2_FpMantRNE_49U_24U_else_acc_nl[22:0];
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_5_itm = MUX_v_23_2_2((inp_lookup_2_FpMantRNE_49U_24U_else_acc_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0);
  assign nl_inp_lookup_3_FpMantRNE_49U_24U_else_acc_nl = (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[47:25])
      + conv_u2u_1_23(FpMantRNE_49U_24U_else_carry_3_sva);
  assign inp_lookup_3_FpMantRNE_49U_24U_else_acc_nl = nl_inp_lookup_3_FpMantRNE_49U_24U_else_acc_nl[22:0];
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_6_itm = MUX_v_23_2_2((inp_lookup_3_FpMantRNE_49U_24U_else_acc_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0);
  assign nl_inp_lookup_4_FpMantRNE_49U_24U_else_acc_nl = (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[47:25])
      + conv_u2u_1_23(FpMantRNE_49U_24U_else_carry_sva);
  assign inp_lookup_4_FpMantRNE_49U_24U_else_acc_nl = nl_inp_lookup_4_FpMantRNE_49U_24U_else_acc_nl[22:0];
  assign FpAdd_8U_23U_FpAdd_8U_23U_or_7_itm = MUX_v_23_2_2((inp_lookup_4_FpMantRNE_49U_24U_else_acc_nl),
      23'b11111111111111111111111, FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0);
  assign IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0 = ~(IsNaN_6U_10U_5_land_lpi_1_dfm_6
      | IsNaN_6U_10U_4_land_lpi_1_dfm_5);
  assign nl_FpAdd_6U_10U_1_is_a_greater_acc_3_nl = ({1'b1 , FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_5_1
      , FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_4_1 , FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_3_0_1})
      + conv_u2u_6_7({(~ FpMul_6U_10U_1_o_expo_lpi_1_dfm_3_5_mx0w1) , (~ FpMul_6U_10U_1_o_expo_lpi_1_dfm_3_4_mx0w1)
      , (~ FpMul_6U_10U_1_o_expo_lpi_1_dfm_3_3_0_mx0w1)}) + 7'b1;
  assign FpAdd_6U_10U_1_is_a_greater_acc_3_nl = nl_FpAdd_6U_10U_1_is_a_greater_acc_3_nl[6:0];
  assign FpAdd_6U_10U_1_is_a_greater_acc_3_itm_6_1 = readslicef_7_1_6((FpAdd_6U_10U_1_is_a_greater_acc_3_nl));
  assign nl_FpAdd_6U_10U_1_is_a_greater_acc_2_nl = ({1'b1 , FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_5_1
      , FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_4_1 , FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_3_0_1})
      + conv_u2u_6_7({(~ FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_5_mx1w1) , (~ FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_4_mx1w1)
      , (~ FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_3_0_mx1w1)}) + 7'b1;
  assign FpAdd_6U_10U_1_is_a_greater_acc_2_nl = nl_FpAdd_6U_10U_1_is_a_greater_acc_2_nl[6:0];
  assign FpAdd_6U_10U_1_is_a_greater_acc_2_itm_6 = readslicef_7_1_6((FpAdd_6U_10U_1_is_a_greater_acc_2_nl));
  assign nl_FpAdd_6U_10U_1_is_a_greater_acc_1_nl = ({1'b1 , FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_5_1
      , FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_4_1 , FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_3_0_1})
      + conv_u2u_6_7({(~ FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_3_5_mx1w1) , (~ FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_3_4_mx1w1)
      , (~ FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_3_3_0_mx1w1)}) + 7'b1;
  assign FpAdd_6U_10U_1_is_a_greater_acc_1_nl = nl_FpAdd_6U_10U_1_is_a_greater_acc_1_nl[6:0];
  assign FpAdd_6U_10U_1_is_a_greater_acc_1_itm_6 = readslicef_7_1_6((FpAdd_6U_10U_1_is_a_greater_acc_1_nl));
  assign nl_FpAdd_6U_10U_1_is_a_greater_acc_nl = ({1'b1 , FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_5_1
      , FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_4_1 , FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_3_0_1})
      + conv_u2u_6_7({(~ FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_3_5_mx1w1) , (~ FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_3_4_mx1w1)
      , (~ FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_3_3_0_mx1w1)}) + 7'b1;
  assign FpAdd_6U_10U_1_is_a_greater_acc_nl = nl_FpAdd_6U_10U_1_is_a_greater_acc_nl[6:0];
  assign FpAdd_6U_10U_1_is_a_greater_acc_itm_6 = readslicef_7_1_6((FpAdd_6U_10U_1_is_a_greater_acc_nl));
  assign FpMantRNE_49U_24U_1_else_carry_1_sva_mx0w2 = (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[25]));
  assign FpMantRNE_49U_24U_1_else_carry_2_sva_mx0w2 = (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[25]));
  assign FpMantRNE_49U_24U_1_else_carry_3_sva_mx0w2 = (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[25]));
  assign FpMantRNE_49U_24U_1_else_carry_sva_mx0w2 = (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[25]));
  assign FpMantRNE_24U_11U_else_carry_2_sva_mx0w1 = (FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_2_mx1[12])
      & ((FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_2_mx1[0]) | (FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_2_mx1[1])
      | (FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_2_mx1[2]) | (FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_2_mx1[3])
      | (FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_2_mx1[4]) | (FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_2_mx1[5])
      | (FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_2_mx1[6]) | (FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_2_mx1[7])
      | (FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_2_mx1[8]) | (FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_2_mx1[9])
      | (FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_2_mx1[10]) | (FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_2_mx1[11])
      | (FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_2_mx1[13]));
  assign FpMantRNE_24U_11U_else_carry_3_sva_mx0w1 = (FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx1[12])
      & ((FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx1[0]) | (FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx1[1])
      | (FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx1[2]) | (FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx1[3])
      | (FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx1[4]) | (FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx1[5])
      | (FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx1[6]) | (FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx1[7])
      | (FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx1[8]) | (FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx1[9])
      | (FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx1[10]) | (FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx1[11])
      | (FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx1[13]));
  assign FpMantRNE_24U_11U_else_carry_sva_mx0w1 = (FpAdd_8U_23U_1_o_mant_lpi_1_dfm_2_mx1[12])
      & ((FpAdd_8U_23U_1_o_mant_lpi_1_dfm_2_mx1[0]) | (FpAdd_8U_23U_1_o_mant_lpi_1_dfm_2_mx1[1])
      | (FpAdd_8U_23U_1_o_mant_lpi_1_dfm_2_mx1[2]) | (FpAdd_8U_23U_1_o_mant_lpi_1_dfm_2_mx1[3])
      | (FpAdd_8U_23U_1_o_mant_lpi_1_dfm_2_mx1[4]) | (FpAdd_8U_23U_1_o_mant_lpi_1_dfm_2_mx1[5])
      | (FpAdd_8U_23U_1_o_mant_lpi_1_dfm_2_mx1[6]) | (FpAdd_8U_23U_1_o_mant_lpi_1_dfm_2_mx1[7])
      | (FpAdd_8U_23U_1_o_mant_lpi_1_dfm_2_mx1[8]) | (FpAdd_8U_23U_1_o_mant_lpi_1_dfm_2_mx1[9])
      | (FpAdd_8U_23U_1_o_mant_lpi_1_dfm_2_mx1[10]) | (FpAdd_8U_23U_1_o_mant_lpi_1_dfm_2_mx1[11])
      | (FpAdd_8U_23U_1_o_mant_lpi_1_dfm_2_mx1[13]));
  assign nl_inp_lookup_1_FpMantRNE_24U_11U_else_acc_nl = (FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_6[22:13])
      + conv_u2u_1_10(FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_8_5_1);
  assign inp_lookup_1_FpMantRNE_24U_11U_else_acc_nl = nl_inp_lookup_1_FpMantRNE_24U_11U_else_acc_nl[9:0];
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_mux_1_nl = MUX_v_10_2_2((FpMantDecShiftRight_23U_8U_10U_o_mant_sum_1_sva[9:0]),
      (inp_lookup_1_FpMantRNE_24U_11U_else_acc_nl), inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_2);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_nl = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_mux_1_nl),
      10'b1111111111, FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_1_lpi_1_dfm_3));
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_mx0w1
      = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_nl), 10'b1111111111,
      FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_1_lpi_1_dfm_2));
  assign nl_inp_lookup_2_FpMantRNE_24U_11U_else_acc_nl = (FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_6[22:13])
      + conv_u2u_1_10(FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_8_5_1);
  assign inp_lookup_2_FpMantRNE_24U_11U_else_acc_nl = nl_inp_lookup_2_FpMantRNE_24U_11U_else_acc_nl[9:0];
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_mux_14_nl = MUX_v_10_2_2((FpMantDecShiftRight_23U_8U_10U_o_mant_sum_2_sva[9:0]),
      (inp_lookup_2_FpMantRNE_24U_11U_else_acc_nl), IsNaN_6U_10U_9_land_2_lpi_1_dfm_8);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_1_nl = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_mux_14_nl),
      10'b1111111111, FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_2_lpi_1_dfm_3));
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_1_mx0w1
      = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_1_nl), 10'b1111111111,
      FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_2_lpi_1_dfm_2));
  assign nl_inp_lookup_3_FpMantRNE_24U_11U_else_acc_nl = (FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_6[22:13])
      + conv_u2u_1_10(FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_8_5_1);
  assign inp_lookup_3_FpMantRNE_24U_11U_else_acc_nl = nl_inp_lookup_3_FpMantRNE_24U_11U_else_acc_nl[9:0];
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_mux_27_nl = MUX_v_10_2_2((FpMantDecShiftRight_23U_8U_10U_o_mant_sum_3_sva[9:0]),
      (inp_lookup_3_FpMantRNE_24U_11U_else_acc_nl), IsNaN_6U_10U_9_land_3_lpi_1_dfm_8);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_2_nl = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_mux_27_nl),
      10'b1111111111, FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_3_lpi_1_dfm_3));
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_2_mx0w1
      = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_2_nl), 10'b1111111111,
      FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_3_lpi_1_dfm_2));
  assign nl_inp_lookup_4_FpMantRNE_24U_11U_else_acc_nl = (FpAdd_8U_23U_1_o_mant_lpi_1_dfm_6[22:13])
      + conv_u2u_1_10(FpMul_6U_10U_1_o_expo_lpi_1_dfm_8_5_1);
  assign inp_lookup_4_FpMantRNE_24U_11U_else_acc_nl = nl_inp_lookup_4_FpMantRNE_24U_11U_else_acc_nl[9:0];
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_mux_40_nl = MUX_v_10_2_2((FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva[9:0]),
      (inp_lookup_4_FpMantRNE_24U_11U_else_acc_nl), IsNaN_6U_10U_9_land_lpi_1_dfm_8);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_3_nl = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_mux_40_nl),
      10'b1111111111, FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_lpi_1_dfm_3));
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_3_mx0w1
      = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_3_nl), 10'b1111111111,
      FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_lpi_1_dfm_2));
  assign inp_lookup_if_unequal_tmp_1_mx0w0 = ~((cfg_precision_1_sva_20==2'b10));
  assign IsNaN_6U_10U_3_IsNaN_6U_10U_3_nor_tmp = ~((~((FpMul_6U_10U_o_mant_1_lpi_1_dfm_3_mx0w0!=10'b0000000000)))
      | (~(FpMul_6U_10U_o_expo_1_lpi_1_dfm_3_5_mx0w0 & FpMul_6U_10U_o_expo_1_lpi_1_dfm_3_4_mx0w0
      & (FpMul_6U_10U_o_expo_1_lpi_1_dfm_3_3_0_mx0w0==4'b1111))));
  assign IsNaN_6U_10U_3_IsNaN_6U_10U_3_nor_1_tmp = ~((~((FpMul_6U_10U_o_mant_2_lpi_1_dfm_3_mx0w0!=10'b0000000000)))
      | (~(FpMul_6U_10U_o_expo_2_lpi_1_dfm_3_5_mx0w0 & FpMul_6U_10U_o_expo_2_lpi_1_dfm_3_4_mx0w0
      & (FpMul_6U_10U_o_expo_2_lpi_1_dfm_3_3_0_mx0w0==4'b1111))));
  assign IsNaN_6U_10U_3_IsNaN_6U_10U_3_nor_2_tmp = ~((~((FpMul_6U_10U_o_mant_3_lpi_1_dfm_3_mx0w0!=10'b0000000000)))
      | (~(FpMul_6U_10U_o_expo_3_lpi_1_dfm_3_5_mx0w0 & FpMul_6U_10U_o_expo_3_lpi_1_dfm_3_4_mx0w0
      & (FpMul_6U_10U_o_expo_3_lpi_1_dfm_3_3_0_mx0w0==4'b1111))));
  assign IsNaN_6U_10U_3_IsNaN_6U_10U_3_nor_3_tmp = ~((~((FpMul_6U_10U_o_mant_lpi_1_dfm_3_mx0w0!=10'b0000000000)))
      | (~(FpMul_6U_10U_o_expo_lpi_1_dfm_3_5_mx0w0 & FpMul_6U_10U_o_expo_lpi_1_dfm_3_4_mx0w0
      & (FpMul_6U_10U_o_expo_lpi_1_dfm_3_3_0_mx0w0==4'b1111))));
  assign FpMantRNE_22U_11U_1_else_carry_2_sva = (FpMul_6U_10U_1_p_mant_20_1_2_lpi_1_dfm_3_mx0[9])
      & (((FpMul_6U_10U_1_p_mant_p1_2_sva_mx1_20_0[0]) & FpMul_6U_10U_1_p_mant_p1_2_sva_mx2_21)
      | (FpMul_6U_10U_1_p_mant_20_1_2_lpi_1_dfm_3_mx0[0]) | (FpMul_6U_10U_1_p_mant_20_1_2_lpi_1_dfm_3_mx0[1])
      | (FpMul_6U_10U_1_p_mant_20_1_2_lpi_1_dfm_3_mx0[2]) | (FpMul_6U_10U_1_p_mant_20_1_2_lpi_1_dfm_3_mx0[3])
      | (FpMul_6U_10U_1_p_mant_20_1_2_lpi_1_dfm_3_mx0[4]) | (FpMul_6U_10U_1_p_mant_20_1_2_lpi_1_dfm_3_mx0[5])
      | (FpMul_6U_10U_1_p_mant_20_1_2_lpi_1_dfm_3_mx0[6]) | (FpMul_6U_10U_1_p_mant_20_1_2_lpi_1_dfm_3_mx0[7])
      | (FpMul_6U_10U_1_p_mant_20_1_2_lpi_1_dfm_3_mx0[8]) | (FpMul_6U_10U_1_p_mant_20_1_2_lpi_1_dfm_3_mx0[10]));
  assign FpMantRNE_22U_11U_2_else_carry_2_sva_mx1w1 = (FpMul_6U_10U_2_p_mant_20_1_2_lpi_1_dfm_3_mx0[9])
      & (((FpMul_6U_10U_2_p_mant_p1_2_sva_mx1_20_0[0]) & FpMul_6U_10U_2_p_mant_p1_2_sva_mx2_21)
      | (FpMul_6U_10U_2_p_mant_20_1_2_lpi_1_dfm_3_mx0[0]) | (FpMul_6U_10U_2_p_mant_20_1_2_lpi_1_dfm_3_mx0[1])
      | (FpMul_6U_10U_2_p_mant_20_1_2_lpi_1_dfm_3_mx0[2]) | (FpMul_6U_10U_2_p_mant_20_1_2_lpi_1_dfm_3_mx0[3])
      | (FpMul_6U_10U_2_p_mant_20_1_2_lpi_1_dfm_3_mx0[4]) | (FpMul_6U_10U_2_p_mant_20_1_2_lpi_1_dfm_3_mx0[5])
      | (FpMul_6U_10U_2_p_mant_20_1_2_lpi_1_dfm_3_mx0[6]) | (FpMul_6U_10U_2_p_mant_20_1_2_lpi_1_dfm_3_mx0[7])
      | (FpMul_6U_10U_2_p_mant_20_1_2_lpi_1_dfm_3_mx0[8]) | (FpMul_6U_10U_2_p_mant_20_1_2_lpi_1_dfm_3_mx0[10]));
  assign FpMantRNE_22U_11U_1_else_carry_sva_mx0w1 = (FpMul_6U_10U_1_p_mant_20_1_lpi_1_dfm_3_mx0[9])
      & (((FpMul_6U_10U_1_p_mant_p1_sva_mx1_20_0[0]) & FpMul_6U_10U_1_p_mant_p1_sva_mx2_21)
      | (FpMul_6U_10U_1_p_mant_20_1_lpi_1_dfm_3_mx0[0]) | (FpMul_6U_10U_1_p_mant_20_1_lpi_1_dfm_3_mx0[1])
      | (FpMul_6U_10U_1_p_mant_20_1_lpi_1_dfm_3_mx0[2]) | (FpMul_6U_10U_1_p_mant_20_1_lpi_1_dfm_3_mx0[3])
      | (FpMul_6U_10U_1_p_mant_20_1_lpi_1_dfm_3_mx0[4]) | (FpMul_6U_10U_1_p_mant_20_1_lpi_1_dfm_3_mx0[5])
      | (FpMul_6U_10U_1_p_mant_20_1_lpi_1_dfm_3_mx0[6]) | (FpMul_6U_10U_1_p_mant_20_1_lpi_1_dfm_3_mx0[7])
      | (FpMul_6U_10U_1_p_mant_20_1_lpi_1_dfm_3_mx0[8]) | (FpMul_6U_10U_1_p_mant_20_1_lpi_1_dfm_3_mx0[10]));
  assign FpMantRNE_22U_11U_2_else_carry_sva_mx0w2 = (FpMul_6U_10U_2_p_mant_20_1_lpi_1_dfm_3_mx0[9])
      & (((FpMul_6U_10U_2_p_mant_p1_sva_mx1_20_0[0]) & FpMul_6U_10U_2_p_mant_p1_sva_mx2_21)
      | (FpMul_6U_10U_2_p_mant_20_1_lpi_1_dfm_3_mx0[0]) | (FpMul_6U_10U_2_p_mant_20_1_lpi_1_dfm_3_mx0[1])
      | (FpMul_6U_10U_2_p_mant_20_1_lpi_1_dfm_3_mx0[2]) | (FpMul_6U_10U_2_p_mant_20_1_lpi_1_dfm_3_mx0[3])
      | (FpMul_6U_10U_2_p_mant_20_1_lpi_1_dfm_3_mx0[4]) | (FpMul_6U_10U_2_p_mant_20_1_lpi_1_dfm_3_mx0[5])
      | (FpMul_6U_10U_2_p_mant_20_1_lpi_1_dfm_3_mx0[6]) | (FpMul_6U_10U_2_p_mant_20_1_lpi_1_dfm_3_mx0[7])
      | (FpMul_6U_10U_2_p_mant_20_1_lpi_1_dfm_3_mx0[8]) | (FpMul_6U_10U_2_p_mant_20_1_lpi_1_dfm_3_mx0[10]));
  assign IsZero_5U_10U_1_aelse_not_21_nl = ~ IsZero_5U_10U_2_land_3_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_26_nl
      = MUX_v_10_2_2(10'b0000000000, (chn_inp_in_rsci_d_mxwt[309:300]), (IsZero_5U_10U_1_aelse_not_21_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux_47_nl = MUX_v_10_2_2(inp_lookup_3_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_itm,
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_26_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_2_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_or_8_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux_47_nl), 10'b1111111111,
      IsInf_5U_10U_1_land_3_lpi_1_dfm);
  assign inp_lookup_3_IsNaN_6U_10U_7_aif_IsNaN_6U_10U_7_aelse_IsNaN_6U_10U_7_aelse_or_tmp
      = (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_3_lpi_1_dfm_8!=10'b0000000000);
  assign nl_inp_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_8U_23U_1_o_expo_lpi_1_dfm_2_mx0w0[7:1])})
      + 8'b1;
  assign inp_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_1_nl = nl_inp_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_1_nl[7:0];
  assign inp_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_1_itm_7_1 = readslicef_8_1_7((inp_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_1_nl));
  assign nl_inp_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_2_mx0w0[7:1])})
      + 8'b1;
  assign inp_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_1_nl = nl_inp_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_1_nl[7:0];
  assign inp_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_1_itm_7 = readslicef_8_1_7((inp_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_1_nl));
  assign nl_inp_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_2_mx0w0[7:1])})
      + 8'b1;
  assign inp_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_1_nl = nl_inp_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_1_nl[7:0];
  assign inp_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_1_itm_7_1 = readslicef_8_1_7((inp_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_1_nl));
  assign nl_inp_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_2_mx0w0[7:1])})
      + 8'b1;
  assign inp_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_1_nl = nl_inp_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_1_nl[7:0];
  assign inp_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_1_itm_7_1 = readslicef_8_1_7((inp_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_1_nl));
  assign IsNaN_6U_10U_IsNaN_6U_10U_nor_tmp = ~((~((FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_1_lpi_1_dfm_5_mx1!=10'b0000000000)))
      | (~(FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_7_5_mx0w0 & (FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_7_4_0_mx0w0==5'b11111))));
  assign inp_lookup_1_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp
      = (FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_21!=10'b0000000000);
  assign IsNaN_6U_10U_1_land_1_lpi_1_dfm_mx0w0 = inp_lookup_1_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp
      & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_12_1_1 & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_12_0_1
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_21==4'b1111);
  assign IsNaN_6U_10U_IsNaN_6U_10U_nor_1_tmp = ~((~((FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_2_lpi_1_dfm_5_mx0!=10'b0000000000)))
      | (~(FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_7_5_mx0w0 & (FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_7_4_0_mx0w0==5'b11111))));
  assign inp_lookup_2_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp
      = (FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_21!=10'b0000000000);
  assign IsNaN_6U_10U_1_land_2_lpi_1_dfm_mx0w0 = inp_lookup_2_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp
      & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_12_1_1 & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_12_0_1
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_21==4'b1111);
  assign IsNaN_6U_10U_IsNaN_6U_10U_nor_2_tmp = ~((~((FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_3_lpi_1_dfm_5_mx0!=10'b0000000000)))
      | (~(FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_7_5_mx0w0 & (FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_7_4_0_mx0w0==5'b11111))));
  assign inp_lookup_3_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp
      = (FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_21!=10'b0000000000);
  assign IsNaN_6U_10U_1_land_3_lpi_1_dfm_mx0w0 = inp_lookup_3_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp
      & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_12_1_1 & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_12_0_1
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_21==4'b1111);
  assign IsNaN_6U_10U_IsNaN_6U_10U_nor_3_tmp = ~((~((FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_lpi_1_dfm_5_mx0!=10'b0000000000)))
      | (~(FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_7_5_mx0w0 & (FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_7_4_0_mx0w0==5'b11111))));
  assign inp_lookup_4_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp
      = (FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_21!=10'b0000000000);
  assign IsNaN_6U_10U_1_land_lpi_1_dfm_mx0w0 = inp_lookup_4_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp
      & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_12_1_1 & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_12_0_1
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_21==4'b1111);
  assign FpMul_6U_10U_FpMul_6U_10U_and_16_nl = (FpMul_6U_10U_o_expo_1_lpi_1_dfm[5])
      & (~ FpMul_6U_10U_lor_9_lpi_1_dfm);
  assign FpMul_6U_10U_o_expo_1_lpi_1_dfm_3_5_mx0w0 = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_14_0_1,
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_14_1_1, (FpMul_6U_10U_FpMul_6U_10U_and_16_nl),
      {IsNaN_6U_10U_land_1_lpi_1_dfm_6 , FpMul_6U_10U_and_ssc , FpMul_6U_10U_FpMul_6U_10U_nor_ssc});
  assign FpMul_6U_10U_FpMul_6U_10U_and_1_nl = (FpMul_6U_10U_o_expo_1_lpi_1_dfm[4])
      & (~ FpMul_6U_10U_lor_9_lpi_1_dfm);
  assign FpMul_6U_10U_o_expo_1_lpi_1_dfm_3_4_mx0w0 = MUX1HOT_s_1_3_2((FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_11_4_0_1[4]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_14_0_1, (FpMul_6U_10U_FpMul_6U_10U_and_1_nl),
      {IsNaN_6U_10U_land_1_lpi_1_dfm_6 , FpMul_6U_10U_and_ssc , FpMul_6U_10U_FpMul_6U_10U_nor_ssc});
  assign FpMul_6U_10U_FpMul_6U_10U_and_18_nl = (FpMul_6U_10U_o_expo_2_lpi_1_dfm[5])
      & (~ FpMul_6U_10U_lor_10_lpi_1_dfm);
  assign FpMul_6U_10U_o_expo_2_lpi_1_dfm_3_5_mx0w0 = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_14_0_1,
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_14_1_1, (FpMul_6U_10U_FpMul_6U_10U_and_18_nl),
      {IsNaN_6U_10U_land_2_lpi_1_dfm_6 , FpMul_6U_10U_and_2_ssc , FpMul_6U_10U_FpMul_6U_10U_nor_1_ssc});
  assign FpMul_6U_10U_FpMul_6U_10U_and_4_nl = (FpMul_6U_10U_o_expo_2_lpi_1_dfm[4])
      & (~ FpMul_6U_10U_lor_10_lpi_1_dfm);
  assign FpMul_6U_10U_o_expo_2_lpi_1_dfm_3_4_mx0w0 = MUX1HOT_s_1_3_2((FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_11_4_0_1[4]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_14_0_1, (FpMul_6U_10U_FpMul_6U_10U_and_4_nl),
      {IsNaN_6U_10U_land_2_lpi_1_dfm_6 , FpMul_6U_10U_and_2_ssc , FpMul_6U_10U_FpMul_6U_10U_nor_1_ssc});
  assign FpMul_6U_10U_FpMul_6U_10U_and_20_nl = (FpMul_6U_10U_o_expo_3_lpi_1_dfm[5])
      & (~ FpMul_6U_10U_lor_11_lpi_1_dfm);
  assign FpMul_6U_10U_o_expo_3_lpi_1_dfm_3_5_mx0w0 = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_14_0_1,
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_14_1_1, (FpMul_6U_10U_FpMul_6U_10U_and_20_nl),
      {IsNaN_6U_10U_land_3_lpi_1_dfm_6 , FpMul_6U_10U_and_4_ssc , FpMul_6U_10U_FpMul_6U_10U_nor_2_ssc});
  assign FpMul_6U_10U_FpMul_6U_10U_and_7_nl = (FpMul_6U_10U_o_expo_3_lpi_1_dfm[4])
      & (~ FpMul_6U_10U_lor_11_lpi_1_dfm);
  assign FpMul_6U_10U_o_expo_3_lpi_1_dfm_3_4_mx0w0 = MUX1HOT_s_1_3_2((FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_11_4_0_1[4]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_14_0_1, (FpMul_6U_10U_FpMul_6U_10U_and_7_nl),
      {IsNaN_6U_10U_land_3_lpi_1_dfm_6 , FpMul_6U_10U_and_4_ssc , FpMul_6U_10U_FpMul_6U_10U_nor_2_ssc});
  assign FpMul_6U_10U_FpMul_6U_10U_and_22_nl = (FpMul_6U_10U_o_expo_lpi_1_dfm[5])
      & (~ FpMul_6U_10U_lor_2_lpi_1_dfm);
  assign FpMul_6U_10U_o_expo_lpi_1_dfm_3_5_mx0w0 = MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_14_0_1,
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_14_1_1, (FpMul_6U_10U_FpMul_6U_10U_and_22_nl),
      {IsNaN_6U_10U_land_lpi_1_dfm_6 , FpMul_6U_10U_and_6_ssc , FpMul_6U_10U_FpMul_6U_10U_nor_3_ssc});
  assign FpMul_6U_10U_FpMul_6U_10U_and_10_nl = (FpMul_6U_10U_o_expo_lpi_1_dfm[4])
      & (~ FpMul_6U_10U_lor_2_lpi_1_dfm);
  assign FpMul_6U_10U_o_expo_lpi_1_dfm_3_4_mx0w0 = MUX1HOT_s_1_3_2((FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_11_4_0_1[4]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_14_0_1, (FpMul_6U_10U_FpMul_6U_10U_and_10_nl),
      {IsNaN_6U_10U_land_lpi_1_dfm_6 , FpMul_6U_10U_and_6_ssc , FpMul_6U_10U_FpMul_6U_10U_nor_3_ssc});
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_1_lpi_1_dfm_5_mx1 = MUX_v_10_2_2((FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_6[9:0]),
      FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_mx0w1,
      FpAdd_6U_10U_1_or_12_cse);
  assign inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0
      = ~(FpMul_6U_10U_1_o_sign_1_lpi_1_dfm_mx0w0 ^ FpMul_6U_10U_2_o_sign_1_lpi_1_dfm_mx0w0);
  assign inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0
      = ~(FpMul_6U_10U_1_o_sign_2_lpi_1_dfm_mx0w0 ^ FpMul_6U_10U_2_o_sign_2_lpi_1_dfm_mx0w0);
  assign inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0
      = ~(FpMul_6U_10U_1_o_sign_3_lpi_1_dfm_mx0w0 ^ FpMul_6U_10U_2_o_sign_3_lpi_1_dfm_mx0w0);
  assign inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0
      = ~(FpMul_6U_10U_1_o_sign_lpi_1_dfm_mx0w0 ^ FpMul_6U_10U_2_o_sign_lpi_1_dfm_mx0w0);
  assign IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_3_tmp = ~((~((FpMul_6U_10U_1_o_mant_lpi_1_dfm_3_mx0w0!=10'b0000000000)))
      | (~(FpMul_6U_10U_1_o_expo_lpi_1_dfm_3_5_mx0w1 & FpMul_6U_10U_1_o_expo_lpi_1_dfm_3_4_mx0w1
      & (FpMul_6U_10U_1_o_expo_lpi_1_dfm_3_3_0_mx0w1==4'b1111))));
  assign IsNaN_6U_10U_9_nor_3_tmp = ~((FpMul_6U_10U_2_o_mant_lpi_1_dfm_7!=10'b0000000000));
  assign IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_2_tmp = ~((~((FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_3_mx0w1!=10'b0000000000)))
      | (~(FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_5_mx1w1 & FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_4_mx1w1
      & (FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_3_0_mx1w1==4'b1111))));
  assign IsNaN_6U_10U_9_nor_2_tmp = ~((FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_8!=10'b0000000000));
  assign IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_1_tmp = ~((~((FpMul_6U_10U_1_o_mant_2_lpi_1_dfm_3!=10'b0000000000)))
      | (~(FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_3_5_mx1w1 & FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_3_4_mx1w1
      & (FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_3_3_0_mx1w1==4'b1111))));
  assign IsNaN_6U_10U_9_nor_1_tmp = ~((FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_8!=10'b0000000000));
  assign IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_tmp = ~((~((FpMul_6U_10U_1_o_mant_1_lpi_1_dfm_3!=10'b0000000000)))
      | (~(FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_3_5_mx1w1 & FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_3_4_mx1w1
      & (FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_3_3_0_mx1w1==4'b1111))));
  assign IsNaN_6U_10U_9_nor_tmp = ~((FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_8!=10'b0000000000));
  assign IsNaN_6U_23U_2_aelse_not_11_nl = ~ IsNaN_6U_23U_2_land_lpi_1_dfm;
  assign FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_22_13_lpi_1_dfm_mx0w1 = MUX_v_10_2_2(10'b0000000000,
      FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_3_itm_2, (IsNaN_6U_23U_2_aelse_not_11_nl));
  assign IsNaN_6U_23U_2_aelse_not_10_nl = ~ IsNaN_6U_23U_2_land_3_lpi_1_dfm;
  assign FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_22_13_3_lpi_1_dfm_mx0w1 = MUX_v_10_2_2(10'b0000000000,
      FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_2_itm_2, (IsNaN_6U_23U_2_aelse_not_10_nl));
  assign IsNaN_6U_23U_2_aelse_not_9_nl = ~ IsNaN_6U_23U_2_land_2_lpi_1_dfm;
  assign FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_22_13_2_lpi_1_dfm_mx0w1 = MUX_v_10_2_2(10'b0000000000,
      FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_1_itm_2, (IsNaN_6U_23U_2_aelse_not_9_nl));
  assign IsNaN_6U_23U_2_aelse_not_8_nl = ~ IsNaN_6U_23U_2_land_1_lpi_1_dfm;
  assign FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_22_13_1_lpi_1_dfm_mx0w1 = MUX_v_10_2_2(10'b0000000000,
      FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_itm_2, (IsNaN_6U_23U_2_aelse_not_8_nl));
  assign nl_inp_lookup_1_FpMantRNE_22U_11U_1_else_acc_nl = FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_21
      + conv_u2u_1_10(FpAdd_8U_23U_o_sign_1_lpi_1_dfm_8);
  assign inp_lookup_1_FpMantRNE_22U_11U_1_else_acc_nl = nl_inp_lookup_1_FpMantRNE_22U_11U_1_else_acc_nl[9:0];
  assign or_5857_nl = FpMantWidthDec_6U_21U_10U_0U_0U_1_if_1_unequal_tmp | (~ FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_9_1);
  assign mux_2032_nl = MUX_v_10_2_2((signext_10_1(~ FpMantWidthDec_6U_21U_10U_0U_0U_1_if_1_unequal_tmp)),
      (inp_lookup_1_FpMantRNE_22U_11U_1_else_acc_nl), or_5857_nl);
  assign FpMul_6U_10U_1_nor_nl = ~(MUX_v_10_2_2((mux_2032_nl), 10'b1111111111, nor_1225_cse));
  assign FpMul_6U_10U_1_FpMul_6U_10U_1_FpMul_6U_10U_1_nor_4_itm = ~(MUX_v_10_2_2((FpMul_6U_10U_1_nor_nl),
      10'b1111111111, FpMul_6U_10U_1_lor_9_lpi_1_dfm));
  assign FpMul_6U_10U_1_or_11_itm = FpMul_6U_10U_1_and_ssc | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_16;
  assign FpMul_6U_10U_1_o_mant_1_lpi_1_dfm_3 = MUX_v_10_2_2(FpMul_6U_10U_1_FpMul_6U_10U_1_FpMul_6U_10U_1_nor_4_itm,
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_21, FpMul_6U_10U_1_or_11_itm);
  assign nl_inp_lookup_2_FpMantRNE_22U_11U_1_else_acc_nl = FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_21
      + conv_u2u_1_10(FpAdd_8U_23U_o_sign_2_lpi_1_dfm_8);
  assign inp_lookup_2_FpMantRNE_22U_11U_1_else_acc_nl = nl_inp_lookup_2_FpMantRNE_22U_11U_1_else_acc_nl[9:0];
  assign or_5858_nl = FpMantWidthDec_6U_21U_10U_0U_0U_1_if_1_unequal_tmp_1 | (~ FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_9_1);
  assign mux_2033_nl = MUX_v_10_2_2((signext_10_1(~ FpMantWidthDec_6U_21U_10U_0U_0U_1_if_1_unequal_tmp_1)),
      (inp_lookup_2_FpMantRNE_22U_11U_1_else_acc_nl), or_5858_nl);
  assign FpMul_6U_10U_1_nor_4_nl = ~(MUX_v_10_2_2((mux_2033_nl), 10'b1111111111,
      nor_1208_cse));
  assign FpMul_6U_10U_1_FpMul_6U_10U_1_FpMul_6U_10U_1_nor_5_itm = ~(MUX_v_10_2_2((FpMul_6U_10U_1_nor_4_nl),
      10'b1111111111, FpMul_6U_10U_1_lor_10_lpi_1_dfm));
  assign FpMul_6U_10U_1_or_10_itm = FpMul_6U_10U_1_and_2_ssc | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_16;
  assign FpMul_6U_10U_1_o_mant_2_lpi_1_dfm_3 = MUX_v_10_2_2(FpMul_6U_10U_1_FpMul_6U_10U_1_FpMul_6U_10U_1_nor_5_itm,
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_21, FpMul_6U_10U_1_or_10_itm);
  assign nl_inp_lookup_4_FpMantRNE_22U_11U_1_else_acc_nl = FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_21
      + conv_u2u_1_10(FpAdd_8U_23U_o_sign_lpi_1_dfm_9);
  assign inp_lookup_4_FpMantRNE_22U_11U_1_else_acc_nl = nl_inp_lookup_4_FpMantRNE_22U_11U_1_else_acc_nl[9:0];
  assign or_5859_nl = FpMantWidthDec_6U_21U_10U_0U_0U_1_if_1_unequal_tmp_3 | (~ FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_9_1);
  assign mux_2034_nl = MUX_v_10_2_2((signext_10_1(~ FpMantWidthDec_6U_21U_10U_0U_0U_1_if_1_unequal_tmp_3)),
      (inp_lookup_4_FpMantRNE_22U_11U_1_else_acc_nl), or_5859_nl);
  assign FpMul_6U_10U_1_nor_6_nl = ~(MUX_v_10_2_2((mux_2034_nl), 10'b1111111111,
      nor_1180_cse));
  assign FpMul_6U_10U_1_FpMul_6U_10U_1_FpMul_6U_10U_1_nor_7_itm = ~(MUX_v_10_2_2((FpMul_6U_10U_1_nor_6_nl),
      10'b1111111111, FpMul_6U_10U_1_lor_2_lpi_1_dfm));
  assign FpMul_6U_10U_1_or_8_itm = FpMul_6U_10U_1_and_6_ssc | IsNaN_6U_10U_4_land_lpi_1_dfm_5;
  assign FpMul_6U_10U_1_o_mant_lpi_1_dfm_3_mx0w0 = MUX_v_10_2_2(FpMul_6U_10U_1_FpMul_6U_10U_1_FpMul_6U_10U_1_nor_7_itm,
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_21, FpMul_6U_10U_1_or_8_itm);
  assign or_6231_cse = IsNaN_6U_10U_7_land_1_lpi_1_dfm_6 | IsNaN_6U_10U_6_land_1_lpi_1_dfm_5;
  assign FpAdd_8U_23U_o_mant_1_lpi_1_dfm_2_mx2 = MUX_v_23_2_2(FpAdd_8U_23U_FpAdd_8U_23U_or_4_itm,
      reg_chn_inp_in_crt_sva_3_510_480_1_reg, or_6231_cse);
  assign or_6230_cse = IsNaN_6U_10U_7_land_2_lpi_1_dfm_6 | IsNaN_6U_10U_6_land_2_lpi_1_dfm_5;
  assign FpAdd_8U_23U_o_mant_2_lpi_1_dfm_2_mx2 = MUX_v_23_2_2(FpAdd_8U_23U_FpAdd_8U_23U_or_5_itm,
      reg_chn_inp_in_crt_sva_3_542_512_1_reg, or_6230_cse);
  assign or_6229_cse = IsNaN_6U_10U_7_land_3_lpi_1_dfm_6 | IsNaN_6U_10U_6_land_3_lpi_1_dfm_5;
  assign FpAdd_8U_23U_o_mant_3_lpi_1_dfm_2_mx2 = MUX_v_23_2_2(FpAdd_8U_23U_FpAdd_8U_23U_or_6_itm,
      reg_chn_inp_in_crt_sva_3_574_544_1_reg, or_6229_cse);
  assign or_6166_nl = IsNaN_6U_10U_7_land_lpi_1_dfm_6 | IsNaN_6U_10U_6_land_lpi_1_dfm_5;
  assign FpAdd_8U_23U_o_mant_lpi_1_dfm_2_mx2 = MUX_v_23_2_2(FpAdd_8U_23U_FpAdd_8U_23U_or_7_itm,
      reg_chn_inp_in_crt_sva_3_606_576_1_reg, or_6166_nl);
  assign IsInf_6U_23U_1_land_1_lpi_1_dfm_mx0w0 = ~((FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_22_13_1_lpi_1_dfm_mx0w1!=10'b0000000000)
      | (FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_9_0_1_lpi_1_dfm!=10'b0000000000)
      | (~ FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_13_1_1));
  assign IsInf_6U_23U_1_land_2_lpi_1_dfm_mx0w0 = ~((FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_22_13_2_lpi_1_dfm_mx0w1!=10'b0000000000)
      | (FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_9_0_2_lpi_1_dfm!=10'b0000000000)
      | (~ FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_13_1_1));
  assign IsInf_6U_23U_1_land_3_lpi_1_dfm_mx0w0 = ~((FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_22_13_3_lpi_1_dfm_mx0w1!=10'b0000000000)
      | (FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_9_0_3_lpi_1_dfm!=10'b0000000000)
      | (~ FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_13_1_1));
  assign IsInf_6U_23U_1_land_lpi_1_dfm_mx0w0 = ~((FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_22_13_lpi_1_dfm_mx0w1!=10'b0000000000)
      | (FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_9_0_lpi_1_dfm!=10'b0000000000)
      | (~ FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_13_1_1));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_3_mx1 = MUX_v_10_2_2((chn_inp_in_rsci_d_mxwt[341:332]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_or_mx0w1,
      or_dcpl_499);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_3_mx1 = MUX_v_10_2_2((chn_inp_in_rsci_d_mxwt[357:348]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_or_4_mx0w1,
      or_dcpl_542);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_3_lpi_1_dfm_3_mx1 = MUX_v_10_2_2((chn_inp_in_rsci_d_mxwt[373:364]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_or_8_mx0w1,
      or_dcpl_585);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_3_mx1 = MUX_v_10_2_2((chn_inp_in_rsci_d_mxwt[389:380]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_or_12_mx0w1,
      or_dcpl_628);
  assign IsNaN_6U_10U_4_nor_tmp = ~((inp_lookup_else_if_a0_9_0_1_lpi_1_dfm_3_mx0w0!=10'b0000000000));
  assign IsNaN_6U_10U_4_land_1_lpi_1_dfm_mx0w1 = ~(IsNaN_6U_10U_4_nor_tmp | (~(inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_3_5_mx0w1
      & (inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_3_4_0_mx0w0==5'b11111))));
  assign IsNaN_6U_10U_4_nor_1_tmp = ~((inp_lookup_else_if_a0_9_0_2_lpi_1_dfm_3_mx0w0!=10'b0000000000));
  assign IsNaN_6U_10U_4_land_2_lpi_1_dfm_mx0w1 = ~(IsNaN_6U_10U_4_nor_1_tmp | (~(inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_3_5_mx0w1
      & (inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_3_4_0_mx0w0==5'b11111))));
  assign IsNaN_6U_10U_4_nor_2_tmp = ~((inp_lookup_else_if_a0_9_0_3_lpi_1_dfm_3_mx0w0!=10'b0000000000));
  assign IsNaN_6U_10U_4_land_3_lpi_1_dfm_mx0w1 = ~(IsNaN_6U_10U_4_nor_2_tmp | (~(inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_3_5_mx0w1
      & (inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_3_4_0_mx0w0==5'b11111))));
  assign IsNaN_6U_10U_4_nor_3_tmp = ~((inp_lookup_else_if_a0_9_0_lpi_1_dfm_3_mx0w0!=10'b0000000000));
  assign IsNaN_6U_10U_4_land_lpi_1_dfm_mx0w1 = ~(IsNaN_6U_10U_4_nor_3_tmp | (~(inp_lookup_else_if_a0_15_10_lpi_1_dfm_3_5_mx0w1
      & (inp_lookup_else_if_a0_15_10_lpi_1_dfm_3_4_0_mx0w0==5'b11111))));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_nl
      = ~((chn_inp_in_rsci_d_mxwt[410]) | IsZero_5U_10U_land_1_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_mux_2_nl = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_1_sva[4]), IsDenorm_5U_10U_land_1_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3_0_mx0w0 = (FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_mux_2_nl)
      | IsInf_5U_10U_land_1_lpi_1_dfm | IsNaN_5U_10U_land_1_lpi_1_dfm;
  assign IsZero_5U_10U_aelse_not_27_nl = ~ IsZero_5U_10U_land_1_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_2_nl =
      MUX_v_4_2_2(4'b0000, (chn_inp_in_rsci_d_mxwt[409:406]), (IsZero_5U_10U_aelse_not_27_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_mux1h_nl =
      MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_2_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_1_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_cse
      , IsDenorm_5U_10U_land_1_lpi_1_dfm , IsInf_5U_10U_land_1_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_mux1h_nl),
      4'b1111, IsNaN_5U_10U_land_1_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_1_nl
      = ~((chn_inp_in_rsci_d_mxwt[426]) | IsZero_5U_10U_land_2_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_mux_7_nl = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_1_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_2_sva[4]), IsDenorm_5U_10U_land_2_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3_0_mx0w0 = (FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_mux_7_nl)
      | IsInf_5U_10U_land_2_lpi_1_dfm | IsNaN_5U_10U_land_2_lpi_1_dfm;
  assign IsZero_5U_10U_aelse_not_26_nl = ~ IsZero_5U_10U_land_2_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_5_nl =
      MUX_v_4_2_2(4'b0000, (chn_inp_in_rsci_d_mxwt[425:422]), (IsZero_5U_10U_aelse_not_26_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_mux1h_1_nl
      = MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_5_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_2_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_1_cse
      , IsDenorm_5U_10U_land_2_lpi_1_dfm , IsInf_5U_10U_land_2_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_mux1h_1_nl),
      4'b1111, IsNaN_5U_10U_land_2_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_2_nl
      = ~((chn_inp_in_rsci_d_mxwt[442]) | IsZero_5U_10U_land_3_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_mux_12_nl = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_2_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_3_sva[4]), IsDenorm_5U_10U_land_3_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3_0_mx0w0 = (FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_mux_12_nl)
      | IsInf_5U_10U_land_3_lpi_1_dfm | IsNaN_5U_10U_land_3_lpi_1_dfm;
  assign IsZero_5U_10U_aelse_not_25_nl = ~ IsZero_5U_10U_land_3_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_8_nl =
      MUX_v_4_2_2(4'b0000, (chn_inp_in_rsci_d_mxwt[441:438]), (IsZero_5U_10U_aelse_not_25_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_mux1h_2_nl
      = MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_8_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_3_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_2_cse
      , IsDenorm_5U_10U_land_3_lpi_1_dfm , IsInf_5U_10U_land_3_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_mux1h_2_nl),
      4'b1111, IsNaN_5U_10U_land_3_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_3_nl
      = ~((chn_inp_in_rsci_d_mxwt[458]) | IsZero_5U_10U_land_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_mux_17_nl = MUX_s_1_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_3_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_sva[4]), IsDenorm_5U_10U_land_lpi_1_dfm);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3_0_mx0w0 = (FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_mux_17_nl)
      | IsInf_5U_10U_land_lpi_1_dfm | IsNaN_5U_10U_land_lpi_1_dfm;
  assign IsZero_5U_10U_aelse_not_24_nl = ~ IsZero_5U_10U_land_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_11_nl
      = MUX_v_4_2_2(4'b0000, (chn_inp_in_rsci_d_mxwt[457:454]), (IsZero_5U_10U_aelse_not_24_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_mux1h_3_nl
      = MUX1HOT_v_4_3_2((FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_11_nl),
      (FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_sva[3:0]), 4'b1110, {FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_3_cse
      , IsDenorm_5U_10U_land_lpi_1_dfm , IsInf_5U_10U_land_lpi_1_dfm});
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w0 = MUX_v_4_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_mux1h_3_nl),
      4'b1111, IsNaN_5U_10U_land_lpi_1_dfm);
  assign IsNaN_6U_10U_6_nor_tmp = ~((FpFractionToFloat_35U_6U_10U_1_o_mant_1_lpi_1_dfm_3_mx0w0!=10'b0000000000));
  assign IsNaN_6U_10U_6_nor_1_tmp = ~((FpFractionToFloat_35U_6U_10U_1_o_mant_2_lpi_1_dfm_3_mx0w0!=10'b0000000000));
  assign IsNaN_6U_10U_6_nor_2_tmp = ~((FpFractionToFloat_35U_6U_10U_1_o_mant_3_lpi_1_dfm_3_mx0w0!=10'b0000000000));
  assign IsNaN_6U_10U_6_nor_3_tmp = ~((FpFractionToFloat_35U_6U_10U_1_o_mant_lpi_1_dfm_3_mx0w0!=10'b0000000000));
  assign IsZero_5U_10U_aelse_not_23_nl = ~ IsZero_5U_10U_land_1_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_nl = MUX_v_10_2_2(10'b0000000000,
      (chn_inp_in_rsci_d_mxwt[405:396]), (IsZero_5U_10U_aelse_not_23_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_mux_4_nl = MUX_v_10_2_2(z_out_16, (FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_mx0w1 =
      MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_mux_4_nl), 10'b1111111111, IsInf_5U_10U_land_1_lpi_1_dfm);
  assign IsZero_5U_10U_aelse_not_22_nl = ~ IsZero_5U_10U_land_2_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_3_nl =
      MUX_v_10_2_2(10'b0000000000, (chn_inp_in_rsci_d_mxwt[421:412]), (IsZero_5U_10U_aelse_not_22_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_mux_36_nl = MUX_v_10_2_2(inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_itm,
      (FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_3_nl), FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_1_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_4_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_mux_36_nl), 10'b1111111111,
      IsInf_5U_10U_land_2_lpi_1_dfm);
  assign IsZero_5U_10U_aelse_not_21_nl = ~ IsZero_5U_10U_land_3_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_6_nl =
      MUX_v_10_2_2(10'b0000000000, (chn_inp_in_rsci_d_mxwt[437:428]), (IsZero_5U_10U_aelse_not_21_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_mux_37_nl = MUX_v_10_2_2(z_out_17, (FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_6_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_2_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_8_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_mux_37_nl), 10'b1111111111,
      IsInf_5U_10U_land_3_lpi_1_dfm);
  assign IsZero_5U_10U_aelse_not_20_nl = ~ IsZero_5U_10U_land_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_9_nl =
      MUX_v_10_2_2(10'b0000000000, (chn_inp_in_rsci_d_mxwt[453:444]), (IsZero_5U_10U_aelse_not_20_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_mux_38_nl = MUX_v_10_2_2(inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_lshift_itm,
      (FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_and_9_nl), FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_3_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_12_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_mux_38_nl), 10'b1111111111,
      IsInf_5U_10U_land_lpi_1_dfm);
  assign IsNaN_6U_10U_2_land_1_lpi_1_dfm_mx0w0 = ((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_1_lpi_1_dfm_3_mx0!=10'b0000000000))
      & (chn_inp_in_rsci_d_mxwt[282]) & FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_3_0_mx0w0
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_6U_10U_2_land_2_lpi_1_dfm_mx0w0 = ((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_2_lpi_1_dfm_3_mx0!=10'b0000000000))
      & (chn_inp_in_rsci_d_mxwt[298]) & FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_3_0_mx0w0
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_6U_10U_2_land_3_lpi_1_dfm_mx0w0 = ((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_3_mx1!=10'b0000000000))
      & (chn_inp_in_rsci_d_mxwt[314]) & FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_3_0_mx0w0
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsNaN_6U_10U_2_land_lpi_1_dfm_mx0w0 = ((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_lpi_1_dfm_3_mx0!=10'b0000000000))
      & (chn_inp_in_rsci_d_mxwt[330]) & FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_3_0_mx0w0
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_3_mx0w0==4'b1111);
  assign IsZero_5U_10U_1_aelse_not_23_nl = ~ IsZero_5U_10U_2_land_1_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_18_nl
      = MUX_v_10_2_2(10'b0000000000, (chn_inp_in_rsci_d_mxwt[277:268]), (IsZero_5U_10U_1_aelse_not_23_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux_43_nl = MUX_v_10_2_2(inp_lookup_1_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_itm,
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_18_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_or_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux_43_nl), 10'b1111111111,
      IsInf_5U_10U_1_land_1_lpi_1_dfm);
  assign IsZero_5U_10U_1_aelse_not_22_nl = ~ IsZero_5U_10U_2_land_2_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_22_nl
      = MUX_v_10_2_2(10'b0000000000, (chn_inp_in_rsci_d_mxwt[293:284]), (IsZero_5U_10U_1_aelse_not_22_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux_45_nl = MUX_v_10_2_2(inp_lookup_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_itm,
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_22_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_1_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_or_4_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux_45_nl), 10'b1111111111,
      IsInf_5U_10U_1_land_2_lpi_1_dfm);
  assign IsZero_5U_10U_1_aelse_not_20_nl = ~ IsZero_5U_10U_2_land_lpi_1_dfm;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_30_nl
      = MUX_v_10_2_2(10'b0000000000, (chn_inp_in_rsci_d_mxwt[325:316]), (IsZero_5U_10U_1_aelse_not_20_nl));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux_49_nl = MUX_v_10_2_2(inp_lookup_4_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_lshift_itm,
      (FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_and_30_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_3_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_or_12_mx0w1
      = MUX_v_10_2_2((FpExpoWidthInc_5U_6U_10U_1U_1U_2_mux_49_nl), 10'b1111111111,
      IsInf_5U_10U_1_land_lpi_1_dfm);
  assign FpAdd_8U_23U_mux_1_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_1_739_395_1[244]),
      (chn_inp_in_crt_sva_1_739_395_1[116]), FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_5);
  assign FpAdd_8U_23U_else_6_mux_mx0w1 = MUX_s_1_2_2((FpAdd_8U_23U_mux_1_nl), (chn_inp_in_crt_sva_1_739_395_1[244]),
      nor_1869_cse);
  assign FpAdd_8U_23U_mux_17_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_1_739_395_1[276]),
      (chn_inp_in_crt_sva_1_739_395_1[148]), FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_5);
  assign FpAdd_8U_23U_else_6_mux_3_mx0w1 = MUX_s_1_2_2((FpAdd_8U_23U_mux_17_nl),
      (chn_inp_in_crt_sva_1_739_395_1[276]), IsNaN_8U_23U_1_land_2_lpi_1_dfm_4);
  assign FpAdd_8U_23U_mux_33_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_1_739_395_1[308]),
      (chn_inp_in_crt_sva_1_739_395_1[180]), FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_5);
  assign FpAdd_8U_23U_else_6_mux_6_mx0w1 = MUX_s_1_2_2((FpAdd_8U_23U_mux_33_nl),
      (chn_inp_in_crt_sva_1_739_395_1[308]), IsNaN_8U_23U_1_land_3_lpi_1_dfm_4);
  assign FpAdd_8U_23U_mux_49_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_1_739_395_1[340]),
      (chn_inp_in_crt_sva_1_739_395_1[212]), FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2);
  assign FpAdd_8U_23U_else_6_mux_9_mx0w1 = MUX_s_1_2_2((FpAdd_8U_23U_mux_49_nl),
      (chn_inp_in_crt_sva_1_739_395_1[340]), IsNaN_8U_23U_1_land_lpi_1_dfm_4);
  assign FpMul_6U_10U_2_o_sign_lpi_1_dfm_mx0w0 = chn_inp_in_crt_sva_2_395_1 & (~
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_14);
  assign FpMul_6U_10U_2_o_sign_3_lpi_1_dfm_mx0w0 = chn_inp_in_crt_sva_2_379_1 & (~
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_14);
  assign FpMul_6U_10U_2_o_sign_2_lpi_1_dfm_mx0w0 = chn_inp_in_crt_sva_2_363_1 & (~
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_14);
  assign FpMul_6U_10U_2_o_sign_1_lpi_1_dfm_mx0w0 = chn_inp_in_crt_sva_2_347_1 & (~
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_14);
  assign FpMul_6U_10U_1_o_sign_lpi_1_dfm_mx0w0 = (chn_inp_in_crt_sva_2_331_268_1[63])
      & (~ IsNaN_6U_10U_4_land_lpi_1_dfm_mx0w1);
  assign FpMul_6U_10U_1_o_sign_3_lpi_1_dfm_mx0w0 = (chn_inp_in_crt_sva_2_331_268_1[47])
      & (~ IsNaN_6U_10U_4_land_3_lpi_1_dfm_mx0w1);
  assign FpMul_6U_10U_1_o_sign_2_lpi_1_dfm_mx0w0 = (chn_inp_in_crt_sva_2_331_268_1[31])
      & (~ IsNaN_6U_10U_4_land_2_lpi_1_dfm_mx0w1);
  assign FpMul_6U_10U_1_o_sign_1_lpi_1_dfm_mx0w0 = (chn_inp_in_crt_sva_2_331_268_1[15])
      & (~ IsNaN_6U_10U_4_land_1_lpi_1_dfm_mx0w1);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_3_mx1 = MUX_v_10_2_2((chn_inp_in_rsci_d_mxwt[405:396]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_mx0w1, or_dcpl_985);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_3_mx1 = MUX_v_10_2_2((chn_inp_in_rsci_d_mxwt[421:412]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_4_mx0w1, or_dcpl_990);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_3_mx1 = MUX_v_10_2_2((chn_inp_in_rsci_d_mxwt[437:428]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_8_mx0w1, or_dcpl_995);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_3_mx1 = MUX_v_10_2_2((chn_inp_in_rsci_d_mxwt[453:444]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_12_mx0w1,
      or_dcpl_1000);
  assign inp_lookup_2_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_mx0w0 = ~((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_2_lpi_1_dfm_3_mx0!=10'b0000000000));
  assign inp_lookup_4_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_mx0w0 = ~((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_lpi_1_dfm_3_mx0!=10'b0000000000));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_3_mx1 = MUX_v_10_2_2((chn_inp_in_rsci_d_mxwt[309:300]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_or_8_mx0w1,
      or_dcpl_818);
  assign IsDenorm_5U_10U_2_land_1_lpi_1_dfm = IsDenorm_5U_10U_2_or_tmp & IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_1_sva;
  assign IsDenorm_5U_10U_2_or_tmp = (chn_inp_in_rsci_d_mxwt[277:268]!=10'b0000000000);
  assign IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_1_sva = ~((chn_inp_in_rsci_d_mxwt[282:278]!=5'b00000));
  assign IsDenorm_5U_10U_land_1_lpi_1_dfm = IsDenorm_5U_10U_or_tmp & IsZero_5U_10U_IsZero_5U_10U_nor_cse_1_sva;
  assign IsDenorm_5U_10U_or_tmp = (chn_inp_in_rsci_d_mxwt[405:396]!=10'b0000000000);
  assign IsZero_5U_10U_IsZero_5U_10U_nor_cse_1_sva = ~((chn_inp_in_rsci_d_mxwt[410:406]!=5'b00000));
  assign FpMantRNE_36U_11U_1_else_carry_1_sva = (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[24])
      & ((inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[0])
      | (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[1])
      | (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[2])
      | (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[3])
      | (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[4])
      | (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[5])
      | (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[6])
      | (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[7])
      | (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[8])
      | (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[9])
      | (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[10])
      | (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[11])
      | (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[12])
      | (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[13])
      | (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[14])
      | (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[15])
      | (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[16])
      | (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[17])
      | (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[18])
      | (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[19])
      | (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[20])
      | (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[21])
      | (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[22])
      | (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[23])
      | (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[25]));
  assign IsDenorm_5U_10U_3_land_1_lpi_1_dfm = IsDenorm_5U_10U_3_or_tmp & IsZero_5U_10U_3_IsZero_5U_10U_3_nor_cse_1_sva;
  assign IsDenorm_5U_10U_3_or_tmp = (chn_inp_in_rsci_d_mxwt[341:332]!=10'b0000000000);
  assign IsZero_5U_10U_3_IsZero_5U_10U_3_nor_cse_1_sva = ~((chn_inp_in_rsci_d_mxwt[346:342]!=5'b00000));
  assign IsDenorm_5U_10U_2_land_2_lpi_1_dfm = IsDenorm_5U_10U_2_or_1_tmp & IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_2_sva;
  assign IsDenorm_5U_10U_2_or_1_tmp = (chn_inp_in_rsci_d_mxwt[293:284]!=10'b0000000000);
  assign IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_2_sva = ~((chn_inp_in_rsci_d_mxwt[298:294]!=5'b00000));
  assign IsDenorm_5U_10U_land_2_lpi_1_dfm = IsDenorm_5U_10U_or_1_tmp & IsZero_5U_10U_IsZero_5U_10U_nor_cse_2_sva;
  assign IsDenorm_5U_10U_or_1_tmp = (chn_inp_in_rsci_d_mxwt[421:412]!=10'b0000000000);
  assign IsZero_5U_10U_IsZero_5U_10U_nor_cse_2_sva = ~((chn_inp_in_rsci_d_mxwt[426:422]!=5'b00000));
  assign FpMantRNE_36U_11U_1_else_carry_2_sva = (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[24])
      & ((inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[0])
      | (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[1])
      | (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[2])
      | (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[3])
      | (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[4])
      | (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[5])
      | (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[6])
      | (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[7])
      | (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[8])
      | (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[9])
      | (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[10])
      | (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[11])
      | (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[12])
      | (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[13])
      | (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[14])
      | (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[15])
      | (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[16])
      | (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[17])
      | (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[18])
      | (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[19])
      | (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[20])
      | (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[21])
      | (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[22])
      | (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[23])
      | (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[25]));
  assign IsDenorm_5U_10U_3_land_2_lpi_1_dfm = IsDenorm_5U_10U_3_or_1_tmp & IsZero_5U_10U_3_IsZero_5U_10U_3_nor_cse_2_sva;
  assign IsDenorm_5U_10U_3_or_1_tmp = (chn_inp_in_rsci_d_mxwt[357:348]!=10'b0000000000);
  assign IsZero_5U_10U_3_IsZero_5U_10U_3_nor_cse_2_sva = ~((chn_inp_in_rsci_d_mxwt[362:358]!=5'b00000));
  assign IsDenorm_5U_10U_2_land_3_lpi_1_dfm = IsDenorm_5U_10U_2_or_2_tmp & IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_3_sva;
  assign IsDenorm_5U_10U_2_or_2_tmp = (chn_inp_in_rsci_d_mxwt[309:300]!=10'b0000000000);
  assign IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_3_sva = ~((chn_inp_in_rsci_d_mxwt[314:310]!=5'b00000));
  assign IsDenorm_5U_10U_land_3_lpi_1_dfm = IsDenorm_5U_10U_or_2_tmp & IsZero_5U_10U_IsZero_5U_10U_nor_cse_3_sva;
  assign IsDenorm_5U_10U_or_2_tmp = (chn_inp_in_rsci_d_mxwt[437:428]!=10'b0000000000);
  assign IsZero_5U_10U_IsZero_5U_10U_nor_cse_3_sva = ~((chn_inp_in_rsci_d_mxwt[442:438]!=5'b00000));
  assign FpMantRNE_36U_11U_1_else_carry_3_sva = (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[24])
      & ((inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[0])
      | (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[1])
      | (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[2])
      | (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[3])
      | (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[4])
      | (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[5])
      | (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[6])
      | (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[7])
      | (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[8])
      | (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[9])
      | (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[10])
      | (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[11])
      | (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[12])
      | (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[13])
      | (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[14])
      | (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[15])
      | (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[16])
      | (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[17])
      | (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[18])
      | (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[19])
      | (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[20])
      | (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[21])
      | (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[22])
      | (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[23])
      | (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[25]));
  assign IsDenorm_5U_10U_3_land_3_lpi_1_dfm = IsDenorm_5U_10U_3_or_2_tmp & IsZero_5U_10U_3_IsZero_5U_10U_3_nor_cse_3_sva;
  assign IsDenorm_5U_10U_3_or_2_tmp = (chn_inp_in_rsci_d_mxwt[373:364]!=10'b0000000000);
  assign IsZero_5U_10U_3_IsZero_5U_10U_3_nor_cse_3_sva = ~((chn_inp_in_rsci_d_mxwt[378:374]!=5'b00000));
  assign IsDenorm_5U_10U_2_land_lpi_1_dfm = IsDenorm_5U_10U_2_or_3_tmp & IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_sva;
  assign IsDenorm_5U_10U_2_or_3_tmp = (chn_inp_in_rsci_d_mxwt[325:316]!=10'b0000000000);
  assign IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_sva = ~((chn_inp_in_rsci_d_mxwt[330:326]!=5'b00000));
  assign IsDenorm_5U_10U_land_lpi_1_dfm = IsDenorm_5U_10U_or_3_tmp & IsZero_5U_10U_IsZero_5U_10U_nor_cse_sva;
  assign IsDenorm_5U_10U_or_3_tmp = (chn_inp_in_rsci_d_mxwt[453:444]!=10'b0000000000);
  assign IsZero_5U_10U_IsZero_5U_10U_nor_cse_sva = ~((chn_inp_in_rsci_d_mxwt[458:454]!=5'b00000));
  assign FpMantRNE_36U_11U_1_else_carry_sva = (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[24])
      & ((inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[0])
      | (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[1])
      | (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[2])
      | (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[3])
      | (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[4])
      | (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[5])
      | (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[6])
      | (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[7])
      | (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[8])
      | (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[9])
      | (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[10])
      | (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[11])
      | (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[12])
      | (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[13])
      | (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[14])
      | (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[15])
      | (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[16])
      | (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[17])
      | (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[18])
      | (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[19])
      | (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[20])
      | (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[21])
      | (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[22])
      | (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[23])
      | (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[25]));
  assign IsDenorm_5U_10U_3_land_lpi_1_dfm = IsDenorm_5U_10U_3_or_3_tmp & IsZero_5U_10U_3_IsZero_5U_10U_3_nor_cse_sva;
  assign IsDenorm_5U_10U_3_or_3_tmp = (chn_inp_in_rsci_d_mxwt[389:380]!=10'b0000000000);
  assign IsZero_5U_10U_3_IsZero_5U_10U_3_nor_cse_sva = ~((chn_inp_in_rsci_d_mxwt[394:390]!=5'b00000));
  assign nl_inp_lookup_1_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_nl = conv_u2u_5_6(IntLeadZero_35U_leading_sign_35_0_rtn_1_sva_2[5:1])
      + 6'b110001;
  assign inp_lookup_1_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_nl = nl_inp_lookup_1_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_nl[5:0];
  assign inp_lookup_1_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_itm_5_1 =
      readslicef_6_1_5((inp_lookup_1_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_nl));
  assign inp_lookup_1_FpMantRNE_36U_11U_else_and_tmp = FpMantRNE_36U_11U_else_carry_1_sva
      & (FpMantRNE_36U_11U_i_data_2_sva[35:25]==11'b11111111111);
  assign FpMantRNE_36U_11U_else_carry_1_sva = (FpMantRNE_36U_11U_i_data_2_sva[24])
      & ((FpMantRNE_36U_11U_i_data_2_sva[0]) | (FpMantRNE_36U_11U_i_data_2_sva[1])
      | (FpMantRNE_36U_11U_i_data_2_sva[2]) | (FpMantRNE_36U_11U_i_data_2_sva[3])
      | (FpMantRNE_36U_11U_i_data_2_sva[4]) | (FpMantRNE_36U_11U_i_data_2_sva[5])
      | (FpMantRNE_36U_11U_i_data_2_sva[6]) | (FpMantRNE_36U_11U_i_data_2_sva[7])
      | (FpMantRNE_36U_11U_i_data_2_sva[8]) | (FpMantRNE_36U_11U_i_data_2_sva[9])
      | (FpMantRNE_36U_11U_i_data_2_sva[10]) | (FpMantRNE_36U_11U_i_data_2_sva[11])
      | (FpMantRNE_36U_11U_i_data_2_sva[12]) | (FpMantRNE_36U_11U_i_data_2_sva[13])
      | (FpMantRNE_36U_11U_i_data_2_sva[14]) | (FpMantRNE_36U_11U_i_data_2_sva[15])
      | (FpMantRNE_36U_11U_i_data_2_sva[16]) | (FpMantRNE_36U_11U_i_data_2_sva[17])
      | (FpMantRNE_36U_11U_i_data_2_sva[18]) | (FpMantRNE_36U_11U_i_data_2_sva[19])
      | (FpMantRNE_36U_11U_i_data_2_sva[20]) | (FpMantRNE_36U_11U_i_data_2_sva[21])
      | (FpMantRNE_36U_11U_i_data_2_sva[22]) | (FpMantRNE_36U_11U_i_data_2_sva[23])
      | (FpMantRNE_36U_11U_i_data_2_sva[25]));
  assign FpFractionToFloat_35U_6U_10U_1_is_zero_1_lpi_1_dfm_1 = ~((FpFractionToFloat_35U_6U_10U_1_if_else_else_if_slc_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_5_mdf_1_sva_2
      | inp_lookup_1_FpMantRNE_36U_11U_1_else_and_svs_2) & FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_st_2);
  assign nl_inp_lookup_2_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_nl = conv_u2u_5_6(IntLeadZero_35U_leading_sign_35_0_rtn_2_sva_2[5:1])
      + 6'b110001;
  assign inp_lookup_2_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_nl = nl_inp_lookup_2_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_nl[5:0];
  assign inp_lookup_2_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_itm_5_1 =
      readslicef_6_1_5((inp_lookup_2_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_nl));
  assign inp_lookup_2_FpMantRNE_36U_11U_else_and_tmp = FpMantRNE_36U_11U_else_carry_2_sva
      & (FpMantRNE_36U_11U_i_data_3_sva[35:25]==11'b11111111111);
  assign FpMantRNE_36U_11U_else_carry_2_sva = (FpMantRNE_36U_11U_i_data_3_sva[24])
      & ((FpMantRNE_36U_11U_i_data_3_sva[0]) | (FpMantRNE_36U_11U_i_data_3_sva[1])
      | (FpMantRNE_36U_11U_i_data_3_sva[2]) | (FpMantRNE_36U_11U_i_data_3_sva[3])
      | (FpMantRNE_36U_11U_i_data_3_sva[4]) | (FpMantRNE_36U_11U_i_data_3_sva[5])
      | (FpMantRNE_36U_11U_i_data_3_sva[6]) | (FpMantRNE_36U_11U_i_data_3_sva[7])
      | (FpMantRNE_36U_11U_i_data_3_sva[8]) | (FpMantRNE_36U_11U_i_data_3_sva[9])
      | (FpMantRNE_36U_11U_i_data_3_sva[10]) | (FpMantRNE_36U_11U_i_data_3_sva[11])
      | (FpMantRNE_36U_11U_i_data_3_sva[12]) | (FpMantRNE_36U_11U_i_data_3_sva[13])
      | (FpMantRNE_36U_11U_i_data_3_sva[14]) | (FpMantRNE_36U_11U_i_data_3_sva[15])
      | (FpMantRNE_36U_11U_i_data_3_sva[16]) | (FpMantRNE_36U_11U_i_data_3_sva[17])
      | (FpMantRNE_36U_11U_i_data_3_sva[18]) | (FpMantRNE_36U_11U_i_data_3_sva[19])
      | (FpMantRNE_36U_11U_i_data_3_sva[20]) | (FpMantRNE_36U_11U_i_data_3_sva[21])
      | (FpMantRNE_36U_11U_i_data_3_sva[22]) | (FpMantRNE_36U_11U_i_data_3_sva[23])
      | (FpMantRNE_36U_11U_i_data_3_sva[25]));
  assign FpFractionToFloat_35U_6U_10U_1_is_zero_2_lpi_1_dfm_1 = ~((FpFractionToFloat_35U_6U_10U_1_if_else_else_if_slc_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_5_mdf_2_sva_2
      | inp_lookup_2_FpMantRNE_36U_11U_1_else_and_svs_2) & FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_st_2);
  assign nl_inp_lookup_3_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_nl = conv_u2u_5_6(IntLeadZero_35U_leading_sign_35_0_rtn_3_sva_2[5:1])
      + 6'b110001;
  assign inp_lookup_3_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_nl = nl_inp_lookup_3_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_nl[5:0];
  assign inp_lookup_3_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_itm_5_1 =
      readslicef_6_1_5((inp_lookup_3_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_nl));
  assign inp_lookup_3_FpMantRNE_36U_11U_else_and_tmp = FpMantRNE_36U_11U_else_carry_3_sva
      & (FpMantRNE_36U_11U_i_data_4_sva[35:25]==11'b11111111111);
  assign FpMantRNE_36U_11U_else_carry_3_sva = (FpMantRNE_36U_11U_i_data_4_sva[24])
      & ((FpMantRNE_36U_11U_i_data_4_sva[0]) | (FpMantRNE_36U_11U_i_data_4_sva[1])
      | (FpMantRNE_36U_11U_i_data_4_sva[2]) | (FpMantRNE_36U_11U_i_data_4_sva[3])
      | (FpMantRNE_36U_11U_i_data_4_sva[4]) | (FpMantRNE_36U_11U_i_data_4_sva[5])
      | (FpMantRNE_36U_11U_i_data_4_sva[6]) | (FpMantRNE_36U_11U_i_data_4_sva[7])
      | (FpMantRNE_36U_11U_i_data_4_sva[8]) | (FpMantRNE_36U_11U_i_data_4_sva[9])
      | (FpMantRNE_36U_11U_i_data_4_sva[10]) | (FpMantRNE_36U_11U_i_data_4_sva[11])
      | (FpMantRNE_36U_11U_i_data_4_sva[12]) | (FpMantRNE_36U_11U_i_data_4_sva[13])
      | (FpMantRNE_36U_11U_i_data_4_sva[14]) | (FpMantRNE_36U_11U_i_data_4_sva[15])
      | (FpMantRNE_36U_11U_i_data_4_sva[16]) | (FpMantRNE_36U_11U_i_data_4_sva[17])
      | (FpMantRNE_36U_11U_i_data_4_sva[18]) | (FpMantRNE_36U_11U_i_data_4_sva[19])
      | (FpMantRNE_36U_11U_i_data_4_sva[20]) | (FpMantRNE_36U_11U_i_data_4_sva[21])
      | (FpMantRNE_36U_11U_i_data_4_sva[22]) | (FpMantRNE_36U_11U_i_data_4_sva[23])
      | (FpMantRNE_36U_11U_i_data_4_sva[25]));
  assign FpFractionToFloat_35U_6U_10U_1_is_zero_3_lpi_1_dfm_1 = ~((FpFractionToFloat_35U_6U_10U_1_if_else_else_if_slc_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_5_mdf_3_sva_2
      | inp_lookup_3_FpMantRNE_36U_11U_1_else_and_svs_2) & FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_st_2);
  assign nl_inp_lookup_4_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_nl = conv_u2u_5_6(IntLeadZero_35U_leading_sign_35_0_rtn_sva_2[5:1])
      + 6'b110001;
  assign inp_lookup_4_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_nl = nl_inp_lookup_4_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_nl[5:0];
  assign inp_lookup_4_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_itm_5_1 =
      readslicef_6_1_5((inp_lookup_4_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_nl));
  assign inp_lookup_4_FpMantRNE_36U_11U_else_and_tmp = FpMantRNE_36U_11U_else_carry_sva
      & (FpMantRNE_36U_11U_i_data_sva[35:25]==11'b11111111111);
  assign FpMantRNE_36U_11U_else_carry_sva = (FpMantRNE_36U_11U_i_data_sva[24]) &
      ((FpMantRNE_36U_11U_i_data_sva[0]) | (FpMantRNE_36U_11U_i_data_sva[1]) | (FpMantRNE_36U_11U_i_data_sva[2])
      | (FpMantRNE_36U_11U_i_data_sva[3]) | (FpMantRNE_36U_11U_i_data_sva[4]) | (FpMantRNE_36U_11U_i_data_sva[5])
      | (FpMantRNE_36U_11U_i_data_sva[6]) | (FpMantRNE_36U_11U_i_data_sva[7]) | (FpMantRNE_36U_11U_i_data_sva[8])
      | (FpMantRNE_36U_11U_i_data_sva[9]) | (FpMantRNE_36U_11U_i_data_sva[10]) |
      (FpMantRNE_36U_11U_i_data_sva[11]) | (FpMantRNE_36U_11U_i_data_sva[12]) | (FpMantRNE_36U_11U_i_data_sva[13])
      | (FpMantRNE_36U_11U_i_data_sva[14]) | (FpMantRNE_36U_11U_i_data_sva[15]) |
      (FpMantRNE_36U_11U_i_data_sva[16]) | (FpMantRNE_36U_11U_i_data_sva[17]) | (FpMantRNE_36U_11U_i_data_sva[18])
      | (FpMantRNE_36U_11U_i_data_sva[19]) | (FpMantRNE_36U_11U_i_data_sva[20]) |
      (FpMantRNE_36U_11U_i_data_sva[21]) | (FpMantRNE_36U_11U_i_data_sva[22]) | (FpMantRNE_36U_11U_i_data_sva[23])
      | (FpMantRNE_36U_11U_i_data_sva[25]));
  assign FpFractionToFloat_35U_6U_10U_1_is_zero_lpi_1_dfm_1 = ~((FpFractionToFloat_35U_6U_10U_1_if_else_else_if_slc_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_5_mdf_sva_2
      | inp_lookup_4_FpMantRNE_36U_11U_1_else_and_svs_2) & FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2);
  assign nl_FpMul_6U_10U_1_oelse_1_acc_nl = conv_u2s_6_7({FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_7_1_1
      , FpAdd_8U_23U_o_sign_1_lpi_1_dfm_7 , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_9})
      + 7'b1100001;
  assign FpMul_6U_10U_1_oelse_1_acc_nl = nl_FpMul_6U_10U_1_oelse_1_acc_nl[6:0];
  assign nl_inp_lookup_1_FpMul_6U_10U_1_oelse_1_acc_nl = conv_s2s_7_8(FpMul_6U_10U_1_oelse_1_acc_nl)
      + conv_u2s_6_8({inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_3_5_mx0w1 , inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_3_4_0_mx0w0});
  assign inp_lookup_1_FpMul_6U_10U_1_oelse_1_acc_nl = nl_inp_lookup_1_FpMul_6U_10U_1_oelse_1_acc_nl[7:0];
  assign inp_lookup_1_FpMul_6U_10U_1_oelse_1_acc_itm_7_1 = readslicef_8_1_7((inp_lookup_1_FpMul_6U_10U_1_oelse_1_acc_nl));
  assign FpMul_6U_10U_1_if_2_FpMul_6U_10U_1_if_2_or_tmp = IsZero_6U_10U_1_IsZero_6U_10U_1_and_itm_8
      | (~((inp_lookup_else_if_a0_9_0_1_lpi_1_dfm_3_mx0w0!=10'b0000000000) | inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_3_5_mx0w1
      | (inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_3_4_0_mx0w0!=5'b00000)));
  assign nl_FpMul_6U_10U_1_oelse_1_acc_1_nl = conv_u2s_6_7({FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_7_1_1
      , FpAdd_8U_23U_o_sign_2_lpi_1_dfm_7 , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_9})
      + 7'b1100001;
  assign FpMul_6U_10U_1_oelse_1_acc_1_nl = nl_FpMul_6U_10U_1_oelse_1_acc_1_nl[6:0];
  assign nl_inp_lookup_2_FpMul_6U_10U_1_oelse_1_acc_nl = conv_s2s_7_8(FpMul_6U_10U_1_oelse_1_acc_1_nl)
      + conv_u2s_6_8({inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_3_5_mx0w1 , inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_3_4_0_mx0w0});
  assign inp_lookup_2_FpMul_6U_10U_1_oelse_1_acc_nl = nl_inp_lookup_2_FpMul_6U_10U_1_oelse_1_acc_nl[7:0];
  assign inp_lookup_2_FpMul_6U_10U_1_oelse_1_acc_itm_7_1 = readslicef_8_1_7((inp_lookup_2_FpMul_6U_10U_1_oelse_1_acc_nl));
  assign FpMul_6U_10U_1_if_2_FpMul_6U_10U_1_if_2_or_2_tmp = IsZero_6U_10U_1_IsZero_6U_10U_1_and_1_itm_6
      | (~((inp_lookup_else_if_a0_9_0_2_lpi_1_dfm_3_mx0w0!=10'b0000000000) | inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_3_5_mx0w1
      | (inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_3_4_0_mx0w0!=5'b00000)));
  assign nl_FpMul_6U_10U_1_oelse_1_acc_2_nl = conv_u2s_6_7({FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_7_1_1
      , FpAdd_8U_23U_o_sign_3_lpi_1_dfm_7 , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_9})
      + 7'b1100001;
  assign FpMul_6U_10U_1_oelse_1_acc_2_nl = nl_FpMul_6U_10U_1_oelse_1_acc_2_nl[6:0];
  assign nl_inp_lookup_3_FpMul_6U_10U_1_oelse_1_acc_nl = conv_s2s_7_8(FpMul_6U_10U_1_oelse_1_acc_2_nl)
      + conv_u2s_6_8({inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_3_5_mx0w1 , inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_3_4_0_mx0w0});
  assign inp_lookup_3_FpMul_6U_10U_1_oelse_1_acc_nl = nl_inp_lookup_3_FpMul_6U_10U_1_oelse_1_acc_nl[7:0];
  assign inp_lookup_3_FpMul_6U_10U_1_oelse_1_acc_itm_7_1 = readslicef_8_1_7((inp_lookup_3_FpMul_6U_10U_1_oelse_1_acc_nl));
  assign FpMul_6U_10U_1_if_2_FpMul_6U_10U_1_if_2_or_4_tmp = IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_itm_8
      | (~((inp_lookup_else_if_a0_9_0_3_lpi_1_dfm_3_mx0w0!=10'b0000000000) | inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_3_5_mx0w1
      | (inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_3_4_0_mx0w0!=5'b00000)));
  assign nl_FpMul_6U_10U_1_oelse_1_acc_3_nl = conv_u2s_6_7({FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_7_1_1
      , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_7_0_1 , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_9})
      + 7'b1100001;
  assign FpMul_6U_10U_1_oelse_1_acc_3_nl = nl_FpMul_6U_10U_1_oelse_1_acc_3_nl[6:0];
  assign nl_inp_lookup_4_FpMul_6U_10U_1_oelse_1_acc_nl = conv_s2s_7_8(FpMul_6U_10U_1_oelse_1_acc_3_nl)
      + conv_u2s_6_8({inp_lookup_else_if_a0_15_10_lpi_1_dfm_3_5_mx0w1 , inp_lookup_else_if_a0_15_10_lpi_1_dfm_3_4_0_mx0w0});
  assign inp_lookup_4_FpMul_6U_10U_1_oelse_1_acc_nl = nl_inp_lookup_4_FpMul_6U_10U_1_oelse_1_acc_nl[7:0];
  assign inp_lookup_4_FpMul_6U_10U_1_oelse_1_acc_itm_7_1 = readslicef_8_1_7((inp_lookup_4_FpMul_6U_10U_1_oelse_1_acc_nl));
  assign FpMul_6U_10U_1_if_2_FpMul_6U_10U_1_if_2_or_6_tmp = IsZero_6U_10U_1_IsZero_6U_10U_1_and_3_itm_6
      | (~((inp_lookup_else_if_a0_9_0_lpi_1_dfm_3_mx0w0!=10'b0000000000) | inp_lookup_else_if_a0_15_10_lpi_1_dfm_3_5_mx0w1
      | (inp_lookup_else_if_a0_15_10_lpi_1_dfm_3_4_0_mx0w0!=5'b00000)));
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_nl = FpAdd_8U_23U_is_inf_1_lpi_1_dfm
      | (~ inp_lookup_1_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1);
  assign FpAdd_8U_23U_is_inf_1_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_is_inf_1_lpi_1_dfm,
      (FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_nl), inp_lookup_1_FpMantRNE_49U_24U_else_and_tmp);
  assign nl_inp_lookup_1_FpAdd_8U_23U_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_8U_23U_o_expo_1_lpi_1_dfm_10[7:1])})
      + 8'b1;
  assign inp_lookup_1_FpAdd_8U_23U_if_4_if_acc_1_nl = nl_inp_lookup_1_FpAdd_8U_23U_if_4_if_acc_1_nl[7:0];
  assign inp_lookup_1_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1 = readslicef_8_1_7((inp_lookup_1_FpAdd_8U_23U_if_4_if_acc_1_nl));
  assign FpAdd_8U_23U_is_inf_1_lpi_1_dfm = ~(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_2
      | (~ (FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_3_49_1_1[48])));
  assign nl_FpAdd_8U_23U_1_is_a_greater_acc_nl = ({1'b1 , FpAdd_8U_23U_o_expo_1_lpi_1_dfm_7_mx1w1})
      + conv_u2u_8_9(~ (chn_inp_in_crt_sva_3_127_0_1[30:23])) + 9'b1;
  assign FpAdd_8U_23U_1_is_a_greater_acc_nl = nl_FpAdd_8U_23U_1_is_a_greater_acc_nl[8:0];
  assign FpAdd_8U_23U_1_is_a_greater_acc_itm_8_1 = readslicef_9_1_8((FpAdd_8U_23U_1_is_a_greater_acc_nl));
  assign FpAdd_8U_23U_and_tmp = inp_lookup_1_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1 &
      inp_lookup_1_FpMantRNE_49U_24U_else_and_tmp;
  assign FpMul_6U_10U_2_FpMul_6U_10U_2_nor_ssc = ~(IsNaN_6U_10U_7_land_1_lpi_1_dfm_6
      | IsNaN_6U_10U_6_land_1_lpi_1_dfm_5);
  assign inp_lookup_1_FpMantRNE_49U_24U_else_and_tmp = FpMantRNE_49U_24U_else_carry_1_sva
      & (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign FpMantRNE_49U_24U_else_carry_1_sva = (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0[25]));
  assign FpNormalize_8U_49U_oelse_not_nl = ~ FpMul_6U_10U_1_lor_6_lpi_1_dfm_5;
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_1_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      FpAdd_8U_23U_int_mant_2_sva_5, (FpNormalize_8U_49U_oelse_not_nl));
  assign FpAdd_8U_23U_int_mant_2_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_1_nl),
      FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_3_49_1_1, FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_3_49_1_1[48]);
  assign nl_inp_lookup_1_IntSaturation_51U_32U_if_acc_nl = conv_s2u_2_3(~ (inp_lookup_if_else_o_acc_psp_1_sva[32:31]))
      + 3'b1;
  assign inp_lookup_1_IntSaturation_51U_32U_if_acc_nl = nl_inp_lookup_1_IntSaturation_51U_32U_if_acc_nl[2:0];
  assign inp_lookup_1_IntSaturation_51U_32U_if_acc_itm_2_1 = readslicef_3_1_2((inp_lookup_1_IntSaturation_51U_32U_if_acc_nl));
  assign nl_inp_lookup_if_else_o_acc_psp_1_sva = conv_s2s_16_33(chn_inp_in_crt_sva_3_331_268_1[15:0])
      + conv_s2s_32_33({inp_lookup_1_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_itm_2
      , inp_lookup_1_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_itm_2
      , inp_lookup_1_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_itm_2});
  assign inp_lookup_if_else_o_acc_psp_1_sva = nl_inp_lookup_if_else_o_acc_psp_1_sva[32:0];
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_1_nl = FpAdd_8U_23U_is_inf_2_lpi_1_dfm
      | (~ inp_lookup_2_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1);
  assign FpAdd_8U_23U_is_inf_2_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_is_inf_2_lpi_1_dfm,
      (FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_1_nl), inp_lookup_2_FpMantRNE_49U_24U_else_and_tmp);
  assign nl_inp_lookup_2_FpAdd_8U_23U_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_8U_23U_o_expo_2_lpi_1_dfm_10[7:1])})
      + 8'b1;
  assign inp_lookup_2_FpAdd_8U_23U_if_4_if_acc_1_nl = nl_inp_lookup_2_FpAdd_8U_23U_if_4_if_acc_1_nl[7:0];
  assign inp_lookup_2_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1 = readslicef_8_1_7((inp_lookup_2_FpAdd_8U_23U_if_4_if_acc_1_nl));
  assign FpAdd_8U_23U_is_inf_2_lpi_1_dfm = ~(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_2
      | (~ (FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_3_49_1_1[48])));
  assign nl_FpAdd_8U_23U_1_is_a_greater_acc_1_nl = ({1'b1 , FpAdd_8U_23U_o_expo_2_lpi_1_dfm_7_mx1w1})
      + conv_u2u_8_9(~ (chn_inp_in_crt_sva_3_127_0_1[62:55])) + 9'b1;
  assign FpAdd_8U_23U_1_is_a_greater_acc_1_nl = nl_FpAdd_8U_23U_1_is_a_greater_acc_1_nl[8:0];
  assign FpAdd_8U_23U_1_is_a_greater_acc_1_itm_8_1 = readslicef_9_1_8((FpAdd_8U_23U_1_is_a_greater_acc_1_nl));
  assign FpAdd_8U_23U_and_1_tmp = inp_lookup_2_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1
      & inp_lookup_2_FpMantRNE_49U_24U_else_and_tmp;
  assign FpMul_6U_10U_2_FpMul_6U_10U_2_nor_1_ssc = ~(IsNaN_6U_10U_7_land_2_lpi_1_dfm_6
      | IsNaN_6U_10U_6_land_2_lpi_1_dfm_5);
  assign inp_lookup_2_FpMantRNE_49U_24U_else_and_tmp = FpMantRNE_49U_24U_else_carry_2_sva
      & (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign FpMantRNE_49U_24U_else_carry_2_sva = (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0[25]));
  assign FpNormalize_8U_49U_oelse_not_1_nl = ~ FpMul_6U_10U_1_lor_7_lpi_1_dfm_5;
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_3_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      FpAdd_8U_23U_int_mant_3_sva_5, (FpNormalize_8U_49U_oelse_not_1_nl));
  assign FpAdd_8U_23U_int_mant_3_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_3_nl),
      FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_3_49_1_1, FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_3_49_1_1[48]);
  assign nl_inp_lookup_2_IntSaturation_51U_32U_if_acc_nl = conv_s2u_2_3(~ (inp_lookup_if_else_o_acc_psp_2_sva[32:31]))
      + 3'b1;
  assign inp_lookup_2_IntSaturation_51U_32U_if_acc_nl = nl_inp_lookup_2_IntSaturation_51U_32U_if_acc_nl[2:0];
  assign inp_lookup_2_IntSaturation_51U_32U_if_acc_itm_2_1 = readslicef_3_1_2((inp_lookup_2_IntSaturation_51U_32U_if_acc_nl));
  assign nl_inp_lookup_if_else_o_acc_psp_2_sva = conv_s2s_16_33(chn_inp_in_crt_sva_3_331_268_1[31:16])
      + conv_s2s_32_33({inp_lookup_2_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_itm_2
      , inp_lookup_2_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_itm_2
      , inp_lookup_2_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_itm_2});
  assign inp_lookup_if_else_o_acc_psp_2_sva = nl_inp_lookup_if_else_o_acc_psp_2_sva[32:0];
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_2_nl = FpAdd_8U_23U_is_inf_3_lpi_1_dfm
      | (~ inp_lookup_3_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1);
  assign FpAdd_8U_23U_is_inf_3_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_is_inf_3_lpi_1_dfm,
      (FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_2_nl), inp_lookup_3_FpMantRNE_49U_24U_else_and_tmp);
  assign nl_inp_lookup_3_FpAdd_8U_23U_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_8U_23U_o_expo_3_lpi_1_dfm_10[7:1])})
      + 8'b1;
  assign inp_lookup_3_FpAdd_8U_23U_if_4_if_acc_1_nl = nl_inp_lookup_3_FpAdd_8U_23U_if_4_if_acc_1_nl[7:0];
  assign inp_lookup_3_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1 = readslicef_8_1_7((inp_lookup_3_FpAdd_8U_23U_if_4_if_acc_1_nl));
  assign FpAdd_8U_23U_is_inf_3_lpi_1_dfm = ~(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_2
      | (~ (FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_3_49_1_1[48])));
  assign nl_FpAdd_8U_23U_1_is_a_greater_acc_2_nl = ({1'b1 , FpAdd_8U_23U_o_expo_3_lpi_1_dfm_7_mx1w1})
      + conv_u2u_8_9(~ (chn_inp_in_crt_sva_3_127_0_1[94:87])) + 9'b1;
  assign FpAdd_8U_23U_1_is_a_greater_acc_2_nl = nl_FpAdd_8U_23U_1_is_a_greater_acc_2_nl[8:0];
  assign FpAdd_8U_23U_1_is_a_greater_acc_2_itm_8_1 = readslicef_9_1_8((FpAdd_8U_23U_1_is_a_greater_acc_2_nl));
  assign FpAdd_8U_23U_and_2_tmp = inp_lookup_3_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1
      & inp_lookup_3_FpMantRNE_49U_24U_else_and_tmp;
  assign FpMul_6U_10U_2_FpMul_6U_10U_2_nor_2_ssc = ~(IsNaN_6U_10U_7_land_3_lpi_1_dfm_6
      | IsNaN_6U_10U_6_land_3_lpi_1_dfm_5);
  assign inp_lookup_3_FpMantRNE_49U_24U_else_and_tmp = FpMantRNE_49U_24U_else_carry_3_sva
      & (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign FpMantRNE_49U_24U_else_carry_3_sva = (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0[25]));
  assign FpNormalize_8U_49U_oelse_not_2_nl = ~ FpMul_6U_10U_1_lor_8_lpi_1_dfm_5;
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_5_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      FpAdd_8U_23U_int_mant_4_sva_5, (FpNormalize_8U_49U_oelse_not_2_nl));
  assign FpAdd_8U_23U_int_mant_4_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_5_nl),
      FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_3_49_1_1, FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_3_49_1_1[48]);
  assign nl_inp_lookup_3_IntSaturation_51U_32U_if_acc_nl = conv_s2u_2_3(~ (inp_lookup_if_else_o_acc_psp_3_sva[32:31]))
      + 3'b1;
  assign inp_lookup_3_IntSaturation_51U_32U_if_acc_nl = nl_inp_lookup_3_IntSaturation_51U_32U_if_acc_nl[2:0];
  assign inp_lookup_3_IntSaturation_51U_32U_if_acc_itm_2_1 = readslicef_3_1_2((inp_lookup_3_IntSaturation_51U_32U_if_acc_nl));
  assign nl_inp_lookup_if_else_o_acc_psp_3_sva = conv_s2s_16_33(chn_inp_in_crt_sva_3_331_268_1[47:32])
      + conv_s2s_32_33({inp_lookup_3_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_itm_2
      , inp_lookup_3_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_itm_2
      , inp_lookup_3_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_itm_2});
  assign inp_lookup_if_else_o_acc_psp_3_sva = nl_inp_lookup_if_else_o_acc_psp_3_sva[32:0];
  assign FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_3_nl = FpAdd_8U_23U_is_inf_lpi_1_dfm
      | (~ inp_lookup_4_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1);
  assign FpAdd_8U_23U_is_inf_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_8U_23U_is_inf_lpi_1_dfm,
      (FpAdd_8U_23U_if_4_FpAdd_8U_23U_if_4_or_3_nl), inp_lookup_4_FpMantRNE_49U_24U_else_and_tmp);
  assign nl_inp_lookup_4_FpAdd_8U_23U_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_8U_23U_o_expo_lpi_1_dfm_10[7:1])})
      + 8'b1;
  assign inp_lookup_4_FpAdd_8U_23U_if_4_if_acc_1_nl = nl_inp_lookup_4_FpAdd_8U_23U_if_4_if_acc_1_nl[7:0];
  assign inp_lookup_4_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1 = readslicef_8_1_7((inp_lookup_4_FpAdd_8U_23U_if_4_if_acc_1_nl));
  assign FpAdd_8U_23U_is_inf_lpi_1_dfm = ~(FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_sva_2
      | (~ (FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_3_49_1_1[48])));
  assign nl_FpAdd_8U_23U_1_is_a_greater_acc_3_nl = ({1'b1 , FpAdd_8U_23U_o_expo_lpi_1_dfm_7_mx1w1})
      + conv_u2u_8_9(~ (chn_inp_in_crt_sva_3_127_0_1[126:119])) + 9'b1;
  assign FpAdd_8U_23U_1_is_a_greater_acc_3_nl = nl_FpAdd_8U_23U_1_is_a_greater_acc_3_nl[8:0];
  assign FpAdd_8U_23U_1_is_a_greater_acc_3_itm_8_1 = readslicef_9_1_8((FpAdd_8U_23U_1_is_a_greater_acc_3_nl));
  assign FpAdd_8U_23U_and_3_tmp = inp_lookup_4_FpAdd_8U_23U_if_4_if_acc_1_itm_7_1
      & inp_lookup_4_FpMantRNE_49U_24U_else_and_tmp;
  assign FpMul_6U_10U_2_FpMul_6U_10U_2_nor_3_ssc = ~(IsNaN_6U_10U_7_land_lpi_1_dfm_6
      | IsNaN_6U_10U_6_land_lpi_1_dfm_5);
  assign inp_lookup_4_FpMantRNE_49U_24U_else_and_tmp = FpMantRNE_49U_24U_else_carry_sva
      & (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[48:25]==24'b111111111111111111111111);
  assign FpMantRNE_49U_24U_else_carry_sva = (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[24])
      & ((FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[0]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[1])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[2]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[3])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[4]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[5])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[6]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[7])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[8]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[9])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[10]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[11])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[12]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[13])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[14]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[15])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[16]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[17])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[18]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[19])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[20]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[21])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[22]) | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[23])
      | (FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0[25]));
  assign FpNormalize_8U_49U_oelse_not_3_nl = ~ FpMul_6U_10U_1_lor_1_lpi_1_dfm_5;
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_7_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      FpAdd_8U_23U_int_mant_1_sva_5, (FpNormalize_8U_49U_oelse_not_3_nl));
  assign FpAdd_8U_23U_int_mant_1_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_7_nl),
      FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_3_49_1_1, FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_3_49_1_1[48]);
  assign nl_inp_lookup_4_IntSaturation_51U_32U_if_acc_nl = conv_s2u_2_3(~ (inp_lookup_if_else_o_acc_psp_sva[32:31]))
      + 3'b1;
  assign inp_lookup_4_IntSaturation_51U_32U_if_acc_nl = nl_inp_lookup_4_IntSaturation_51U_32U_if_acc_nl[2:0];
  assign inp_lookup_4_IntSaturation_51U_32U_if_acc_itm_2_1 = readslicef_3_1_2((inp_lookup_4_IntSaturation_51U_32U_if_acc_nl));
  assign nl_inp_lookup_if_else_o_acc_psp_sva = conv_s2s_16_33(chn_inp_in_crt_sva_3_331_268_1[63:48])
      + conv_s2s_32_33({inp_lookup_4_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_itm_2
      , inp_lookup_4_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_itm_2
      , inp_lookup_4_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_itm_2});
  assign inp_lookup_if_else_o_acc_psp_sva = nl_inp_lookup_if_else_o_acc_psp_sva[32:0];
  assign nl_inp_lookup_1_FpMul_6U_10U_1_else_2_else_if_if_acc_nl = reg_FpAdd_8U_23U_o_expo_1_lpi_1_dfm_11_1_reg
      + 6'b1;
  assign inp_lookup_1_FpMul_6U_10U_1_else_2_else_if_if_acc_nl = nl_inp_lookup_1_FpMul_6U_10U_1_else_2_else_if_if_acc_nl[5:0];
  assign FpMul_6U_10U_1_p_expo_1_lpi_1_dfm_1_mx0 = MUX_v_6_2_2(reg_FpAdd_8U_23U_o_expo_1_lpi_1_dfm_11_1_reg,
      (inp_lookup_1_FpMul_6U_10U_1_else_2_else_if_if_acc_nl), FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5);
  assign FpMantWidthDec_6U_21U_10U_0U_0U_1_if_1_unequal_tmp = ~((FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_1_sva_1==6'b111111));
  assign nl_FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_1_sva_1 = FpMul_6U_10U_1_p_expo_1_lpi_1_dfm_1_mx0
      + 6'b1;
  assign FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_1_sva_1 = nl_FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_1_sva_1[5:0];
  assign FpMul_6U_10U_1_lor_9_lpi_1_dfm = (~((FpMul_6U_10U_1_o_expo_1_lpi_1_dfm!=6'b000000)))
      | FpMul_6U_10U_1_lor_6_lpi_1_dfm_6;
  assign FpMul_6U_10U_1_FpMul_6U_10U_1_nor_ssc = ~(IsNaN_6U_10U_5_land_1_lpi_1_dfm_6
      | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_16);
  assign FpMul_6U_10U_1_and_ssc = IsNaN_6U_10U_5_land_1_lpi_1_dfm_6 & (~ IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_16);
  assign FpMul_6U_10U_1_or_4_nl = ((~ FpMantWidthDec_6U_21U_10U_0U_0U_1_if_1_unequal_tmp)
      & FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_9_1) | nor_1225_cse;
  assign FpMantWidthDec_6U_21U_10U_0U_0U_1_and_1_nl = FpMantWidthDec_6U_21U_10U_0U_0U_1_if_1_unequal_tmp
      & FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_9_1 & (~ nor_1225_cse);
  assign FpMul_6U_10U_1_o_expo_1_lpi_1_dfm = MUX1HOT_v_6_3_2(FpMul_6U_10U_1_p_expo_1_lpi_1_dfm_1_mx0,
      6'b111110, FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_1_sva_1, {nor_1224_cse
      , (FpMul_6U_10U_1_or_4_nl) , (FpMantWidthDec_6U_21U_10U_0U_0U_1_and_1_nl)});
  assign nl_inp_lookup_2_FpMul_6U_10U_1_else_2_else_if_if_acc_nl = reg_FpAdd_8U_23U_o_expo_2_lpi_1_dfm_11_1_reg
      + 6'b1;
  assign inp_lookup_2_FpMul_6U_10U_1_else_2_else_if_if_acc_nl = nl_inp_lookup_2_FpMul_6U_10U_1_else_2_else_if_if_acc_nl[5:0];
  assign FpMul_6U_10U_1_p_expo_2_lpi_1_dfm_1_mx0 = MUX_v_6_2_2(reg_FpAdd_8U_23U_o_expo_2_lpi_1_dfm_11_1_reg,
      (inp_lookup_2_FpMul_6U_10U_1_else_2_else_if_if_acc_nl), FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5);
  assign FpMantWidthDec_6U_21U_10U_0U_0U_1_if_1_unequal_tmp_1 = ~((FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_2_sva_1==6'b111111));
  assign nl_FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_2_sva_1 = FpMul_6U_10U_1_p_expo_2_lpi_1_dfm_1_mx0
      + 6'b1;
  assign FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_2_sva_1 = nl_FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_2_sva_1[5:0];
  assign FpMul_6U_10U_1_lor_10_lpi_1_dfm = (~((FpMul_6U_10U_1_o_expo_2_lpi_1_dfm!=6'b000000)))
      | FpMul_6U_10U_1_lor_7_lpi_1_dfm_6;
  assign FpMul_6U_10U_1_FpMul_6U_10U_1_nor_1_ssc = ~(IsNaN_6U_10U_5_land_2_lpi_1_dfm_6
      | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_16);
  assign FpMul_6U_10U_1_and_2_ssc = IsNaN_6U_10U_5_land_2_lpi_1_dfm_6 & (~ IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_16);
  assign FpMul_6U_10U_1_or_5_nl = ((~ FpMantWidthDec_6U_21U_10U_0U_0U_1_if_1_unequal_tmp_1)
      & FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_9_1) | nor_1208_cse;
  assign FpMantWidthDec_6U_21U_10U_0U_0U_1_and_3_nl = FpMantWidthDec_6U_21U_10U_0U_0U_1_if_1_unequal_tmp_1
      & FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_9_1 & (~ nor_1208_cse);
  assign FpMul_6U_10U_1_o_expo_2_lpi_1_dfm = MUX1HOT_v_6_3_2(FpMul_6U_10U_1_p_expo_2_lpi_1_dfm_1_mx0,
      6'b111110, FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_2_sva_1, {nor_1207_cse
      , (FpMul_6U_10U_1_or_5_nl) , (FpMantWidthDec_6U_21U_10U_0U_0U_1_and_3_nl)});
  assign nl_inp_lookup_3_FpMul_6U_10U_1_else_2_else_if_if_acc_nl = reg_FpAdd_8U_23U_o_expo_3_lpi_1_dfm_11_1_reg
      + 6'b1;
  assign inp_lookup_3_FpMul_6U_10U_1_else_2_else_if_if_acc_nl = nl_inp_lookup_3_FpMul_6U_10U_1_else_2_else_if_if_acc_nl[5:0];
  assign FpMul_6U_10U_1_p_expo_3_lpi_1_dfm_1_mx0 = MUX_v_6_2_2(reg_FpAdd_8U_23U_o_expo_3_lpi_1_dfm_11_1_reg,
      (inp_lookup_3_FpMul_6U_10U_1_else_2_else_if_if_acc_nl), FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5);
  assign FpMantWidthDec_6U_21U_10U_0U_0U_1_if_1_unequal_tmp_2 = ~((FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_3_sva_1==6'b111111));
  assign nl_FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_3_sva_1 = FpMul_6U_10U_1_p_expo_3_lpi_1_dfm_1_mx0
      + 6'b1;
  assign FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_3_sva_1 = nl_FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_3_sva_1[5:0];
  assign FpMul_6U_10U_1_lor_11_lpi_1_dfm = (~((FpMul_6U_10U_1_o_expo_3_lpi_1_dfm!=6'b000000)))
      | FpMul_6U_10U_1_lor_8_lpi_1_dfm_6;
  assign FpMul_6U_10U_1_FpMul_6U_10U_1_nor_2_ssc = ~(IsNaN_6U_10U_5_land_3_lpi_1_dfm_6
      | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_16);
  assign FpMul_6U_10U_1_and_4_ssc = IsNaN_6U_10U_5_land_3_lpi_1_dfm_6 & (~ IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_16);
  assign FpMul_6U_10U_1_or_6_nl = ((~ FpMantWidthDec_6U_21U_10U_0U_0U_1_if_1_unequal_tmp_2)
      & FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_9_1) | nor_1191_cse;
  assign FpMantWidthDec_6U_21U_10U_0U_0U_1_and_5_nl = FpMantWidthDec_6U_21U_10U_0U_0U_1_if_1_unequal_tmp_2
      & FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_9_1 & (~ nor_1191_cse);
  assign FpMul_6U_10U_1_o_expo_3_lpi_1_dfm = MUX1HOT_v_6_3_2(FpMul_6U_10U_1_p_expo_3_lpi_1_dfm_1_mx0,
      6'b111110, FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_3_sva_1, {nor_1190_cse
      , (FpMul_6U_10U_1_or_6_nl) , (FpMantWidthDec_6U_21U_10U_0U_0U_1_and_5_nl)});
  assign nl_inp_lookup_4_FpMul_6U_10U_1_else_2_else_if_if_acc_nl = reg_FpAdd_8U_23U_o_expo_lpi_1_dfm_11_1_reg
      + 6'b1;
  assign inp_lookup_4_FpMul_6U_10U_1_else_2_else_if_if_acc_nl = nl_inp_lookup_4_FpMul_6U_10U_1_else_2_else_if_if_acc_nl[5:0];
  assign FpMul_6U_10U_1_p_expo_lpi_1_dfm_1_mx0 = MUX_v_6_2_2(reg_FpAdd_8U_23U_o_expo_lpi_1_dfm_11_1_reg,
      (inp_lookup_4_FpMul_6U_10U_1_else_2_else_if_if_acc_nl), FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5);
  assign FpMantWidthDec_6U_21U_10U_0U_0U_1_if_1_unequal_tmp_3 = ~((FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_sva_1==6'b111111));
  assign nl_FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_sva_1 = FpMul_6U_10U_1_p_expo_lpi_1_dfm_1_mx0
      + 6'b1;
  assign FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_sva_1 = nl_FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_sva_1[5:0];
  assign FpMul_6U_10U_1_lor_2_lpi_1_dfm = (~((FpMul_6U_10U_1_o_expo_lpi_1_dfm!=6'b000000)))
      | FpMul_6U_10U_1_lor_1_lpi_1_dfm_6;
  assign FpMul_6U_10U_1_and_6_ssc = IsNaN_6U_10U_5_land_lpi_1_dfm_6 & (~ IsNaN_6U_10U_4_land_lpi_1_dfm_5);
  assign FpMul_6U_10U_1_FpMul_6U_10U_1_nor_11_nl = ~(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_9_1
      | nor_1180_cse);
  assign FpMul_6U_10U_1_or_7_nl = ((~ FpMantWidthDec_6U_21U_10U_0U_0U_1_if_1_unequal_tmp_3)
      & FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_9_1) | nor_1180_cse;
  assign FpMantWidthDec_6U_21U_10U_0U_0U_1_and_7_nl = FpMantWidthDec_6U_21U_10U_0U_0U_1_if_1_unequal_tmp_3
      & FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_9_1 & (~ nor_1180_cse);
  assign FpMul_6U_10U_1_o_expo_lpi_1_dfm = MUX1HOT_v_6_3_2(FpMul_6U_10U_1_p_expo_lpi_1_dfm_1_mx0,
      6'b111110, FpMantWidthDec_6U_21U_10U_0U_0U_1_o_expo_sva_1, {(FpMul_6U_10U_1_FpMul_6U_10U_1_nor_11_nl)
      , (FpMul_6U_10U_1_or_7_nl) , (FpMantWidthDec_6U_21U_10U_0U_0U_1_and_7_nl)});
  assign nl_inp_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_1_nl = ({1'b1 , (reg_FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_7_1_itm[7:1])})
      + 8'b1;
  assign inp_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_1_nl = nl_inp_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_1_nl[7:0];
  assign inp_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_1_itm_7_1 = readslicef_8_1_7((inp_lookup_1_FpAdd_8U_23U_1_if_3_if_acc_1_nl));
  assign FpNormalize_8U_49U_1_FpNormalize_8U_49U_1_and_1_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      inp_lookup_1_FpNormalize_8U_49U_1_else_lshift_itm, FpNormalize_8U_49U_1_oelse_not_9);
  assign FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_1_FpNormalize_8U_49U_1_and_1_nl),
      (FpAdd_8U_23U_1_int_mant_p1_1_sva_3[49:1]), FpAdd_8U_23U_1_int_mant_p1_1_sva_3[49]);
  assign nl_FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_22})
      + conv_u2u_10_11({(~ reg_FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_7_itm) , (~ reg_FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_7_1_itm)})
      + 11'b1;
  assign FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_nl = nl_FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_nl[10:0];
  assign FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_itm_10 = readslicef_11_1_10((FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_nl));
  assign nl_inp_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_1_nl = ({1'b1 , (reg_FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_7_1_itm[7:1])})
      + 8'b1;
  assign inp_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_1_nl = nl_inp_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_1_nl[7:0];
  assign inp_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_1_itm_7_1 = readslicef_8_1_7((inp_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_1_nl));
  assign FpNormalize_8U_49U_1_FpNormalize_8U_49U_1_and_3_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      inp_lookup_2_FpNormalize_8U_49U_1_else_lshift_itm, FpNormalize_8U_49U_1_oelse_not_11);
  assign FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_1_FpNormalize_8U_49U_1_and_3_nl),
      (FpAdd_8U_23U_1_int_mant_p1_2_sva_3[49:1]), FpAdd_8U_23U_1_int_mant_p1_2_sva_3[49]);
  assign nl_FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_1_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_22})
      + conv_u2u_10_11({(~ reg_FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_7_itm) , (~ reg_FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_7_1_itm)})
      + 11'b1;
  assign FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_1_nl = nl_FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_1_nl[10:0];
  assign FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_1_itm_10 = readslicef_11_1_10((FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_1_nl));
  assign nl_inp_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_1_nl = ({1'b1 , (reg_FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_7_1_itm[7:1])})
      + 8'b1;
  assign inp_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_1_nl = nl_inp_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_1_nl[7:0];
  assign inp_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_1_itm_7 = readslicef_8_1_7((inp_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_1_nl));
  assign FpNormalize_8U_49U_1_FpNormalize_8U_49U_1_and_5_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      inp_lookup_3_FpNormalize_8U_49U_1_else_lshift_itm, FpNormalize_8U_49U_1_oelse_not_13);
  assign FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_1_FpNormalize_8U_49U_1_and_5_nl),
      (FpAdd_8U_23U_1_int_mant_p1_3_sva_3[49:1]), FpAdd_8U_23U_1_int_mant_p1_3_sva_3[49]);
  assign nl_FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_2_nl = ({1'b1 , reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_6_itm
      , reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_6_1_itm}) + conv_u2u_10_11({(~ reg_FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_7_itm)
      , (~ reg_FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_7_1_itm)}) + 11'b1;
  assign FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_2_nl = nl_FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_2_nl[10:0];
  assign FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_2_itm_10 = readslicef_11_1_10((FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_2_nl));
  assign nl_inp_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_1_nl = ({1'b1 , (reg_FpMul_6U_10U_2_o_mant_lpi_1_dfm_7_1_reg[7:1])})
      + 8'b1;
  assign inp_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_1_nl = nl_inp_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_1_nl[7:0];
  assign inp_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_1_itm_7_1 = readslicef_8_1_7((inp_lookup_4_FpAdd_8U_23U_1_if_3_if_acc_1_nl));
  assign FpNormalize_8U_49U_1_FpNormalize_8U_49U_1_and_7_nl = MUX_v_49_2_2(49'b0000000000000000000000000000000000000000000000000,
      inp_lookup_4_FpNormalize_8U_49U_1_else_lshift_itm, FpNormalize_8U_49U_1_oelse_not_15);
  assign FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0 = MUX_v_49_2_2((FpNormalize_8U_49U_1_FpNormalize_8U_49U_1_and_7_nl),
      (FpAdd_8U_23U_1_int_mant_p1_sva_3[49:1]), FpAdd_8U_23U_1_int_mant_p1_sva_3[49]);
  assign nl_FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_3_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_22})
      + conv_u2u_10_11({(~ reg_FpMul_6U_10U_2_o_mant_lpi_1_dfm_7_reg) , (~ reg_FpMul_6U_10U_2_o_mant_lpi_1_dfm_7_1_reg)})
      + 11'b1;
  assign FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_3_nl = nl_FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_3_nl[10:0];
  assign FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_3_itm_10 = readslicef_11_1_10((FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_3_nl));
  assign FpAdd_8U_23U_1_and_tmp = FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_7_4_1 & inp_lookup_1_FpMantRNE_49U_24U_1_else_and_svs_2;
  assign FpAdd_8U_23U_1_if_4_FpAdd_8U_23U_1_if_4_or_4_nl = FpAdd_6U_10U_1_is_a_greater_lor_1_lpi_1_dfm_5
      | (~ FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_7_4_1);
  assign FpAdd_8U_23U_1_is_inf_1_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_1_is_a_greater_lor_1_lpi_1_dfm_5,
      (FpAdd_8U_23U_1_if_4_FpAdd_8U_23U_1_if_4_or_4_nl), inp_lookup_1_FpMantRNE_49U_24U_1_else_and_svs_2);
  assign FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_5_m1c = ~(IsNaN_8U_23U_3_land_1_lpi_1_dfm_7
      | IsNaN_6U_10U_8_land_1_lpi_1_dfm_st_3);
  assign nl_FpAdd_6U_10U_1_int_mant_p1_1_sva = conv_u2u_23_24(FpAdd_6U_10U_1_addend_larger_qr_1_lpi_1_dfm_mx0)
      + conv_u2u_23_24(FpAdd_6U_10U_1_addend_smaller_qr_1_lpi_1_dfm_mx0);
  assign FpAdd_6U_10U_1_int_mant_p1_1_sva = nl_FpAdd_6U_10U_1_int_mant_p1_1_sva[23:0];
  assign FpAdd_6U_10U_1_addend_larger_qr_1_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_1_b_int_mant_p1_1_sva_2,
      reg_chn_inp_in_crt_sva_6_30_0_1_reg, FpAdd_6U_10U_1_is_a_greater_lor_1_lpi_1_dfm_5);
  assign FpAdd_6U_10U_1_addend_smaller_qr_1_lpi_1_dfm_mx0 = MUX_v_23_2_2(reg_chn_inp_in_crt_sva_6_30_0_1_reg,
      FpAdd_6U_10U_1_b_int_mant_p1_1_sva_2, FpAdd_6U_10U_1_is_a_greater_lor_1_lpi_1_dfm_5);
  assign nl_FpAdd_6U_10U_1_int_mant_p1_1_sva_1 = ({1'b1 , (~ FpAdd_6U_10U_1_addend_smaller_qr_1_lpi_1_dfm_mx0)})
      + conv_u2u_23_24(FpAdd_6U_10U_1_addend_larger_qr_1_lpi_1_dfm_mx0) + 24'b1;
  assign FpAdd_6U_10U_1_int_mant_p1_1_sva_1 = nl_FpAdd_6U_10U_1_int_mant_p1_1_sva_1[23:0];
  assign FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_mx0 = MUX_v_24_2_2(FpAdd_6U_10U_1_int_mant_p1_1_sva_1,
      FpAdd_6U_10U_1_int_mant_p1_1_sva, IsNaN_8U_23U_3_land_1_lpi_1_dfm_7);
  assign nl_inp_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_nl = FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_13
      + 8'b1;
  assign inp_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_nl = nl_inp_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_nl[7:0];
  assign FpAdd_8U_23U_1_or_1_nl = ((~(FpAdd_8U_23U_1_and_1_tmp | FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_2_mx0))
      & FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_7_m1c) | (IsNaN_8U_23U_3_land_2_lpi_1_dfm_7
      & (~ IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_4));
  assign FpAdd_8U_23U_1_and_13_nl = FpAdd_8U_23U_1_and_1_tmp & (~ FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_2_mx0)
      & FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_7_m1c;
  assign FpAdd_8U_23U_1_and_30_nl = FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_2_mx0 & FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_7_m1c;
  assign FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_7 = MUX1HOT_v_8_4_2(FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_13,
      (inp_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_nl), 8'b11111110, reg_chn_inp_in_crt_sva_6_62_32_reg,
      {(FpAdd_8U_23U_1_or_1_nl) , (FpAdd_8U_23U_1_and_13_nl) , (FpAdd_8U_23U_1_and_30_nl)
      , IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_4});
  assign FpAdd_8U_23U_1_and_1_tmp = FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_7_4_1 & inp_lookup_2_FpMantRNE_49U_24U_1_else_and_svs_2;
  assign FpAdd_8U_23U_1_if_4_FpAdd_8U_23U_1_if_4_or_5_nl = FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_5
      | (~ FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_7_4_1);
  assign FpAdd_8U_23U_1_is_inf_2_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_5,
      (FpAdd_8U_23U_1_if_4_FpAdd_8U_23U_1_if_4_or_5_nl), inp_lookup_2_FpMantRNE_49U_24U_1_else_and_svs_2);
  assign FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_7_m1c = ~(IsNaN_8U_23U_3_land_2_lpi_1_dfm_7
      | IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_4);
  assign nl_FpAdd_6U_10U_1_int_mant_p1_2_sva = conv_u2u_23_24(FpAdd_6U_10U_1_addend_larger_qr_2_lpi_1_dfm_mx0)
      + conv_u2u_23_24(FpAdd_6U_10U_1_addend_smaller_qr_2_lpi_1_dfm_mx0);
  assign FpAdd_6U_10U_1_int_mant_p1_2_sva = nl_FpAdd_6U_10U_1_int_mant_p1_2_sva[23:0];
  assign FpAdd_6U_10U_1_addend_larger_qr_2_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_1_b_int_mant_p1_2_sva_2,
      reg_chn_inp_in_crt_sva_6_62_32_1_reg, FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_5);
  assign FpAdd_6U_10U_1_addend_smaller_qr_2_lpi_1_dfm_mx0 = MUX_v_23_2_2(reg_chn_inp_in_crt_sva_6_62_32_1_reg,
      FpAdd_6U_10U_1_b_int_mant_p1_2_sva_2, FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_5);
  assign nl_FpAdd_6U_10U_1_int_mant_p1_2_sva_1 = ({1'b1 , (~ FpAdd_6U_10U_1_addend_smaller_qr_2_lpi_1_dfm_mx0)})
      + conv_u2u_23_24(FpAdd_6U_10U_1_addend_larger_qr_2_lpi_1_dfm_mx0) + 24'b1;
  assign FpAdd_6U_10U_1_int_mant_p1_2_sva_1 = nl_FpAdd_6U_10U_1_int_mant_p1_2_sva_1[23:0];
  assign FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_mx0 = MUX_v_24_2_2(FpAdd_6U_10U_1_int_mant_p1_2_sva_1,
      FpAdd_6U_10U_1_int_mant_p1_2_sva, IsNaN_8U_23U_3_land_2_lpi_1_dfm_7);
  assign nl_inp_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_nl = reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_7_1_itm
      + 8'b1;
  assign inp_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_nl = nl_inp_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_nl[7:0];
  assign FpAdd_8U_23U_1_or_2_nl = ((~(FpAdd_8U_23U_1_and_2_tmp | FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_2_mx0))
      & FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_9_m1c) | (IsNaN_8U_23U_3_land_3_lpi_1_dfm_7
      & (~ IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_4));
  assign FpAdd_8U_23U_1_and_19_nl = FpAdd_8U_23U_1_and_2_tmp & (~ FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_2_mx0)
      & FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_9_m1c;
  assign FpAdd_8U_23U_1_and_32_nl = FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_2_mx0 & FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_9_m1c;
  assign FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_7 = MUX1HOT_v_8_4_2(reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_7_1_itm,
      (inp_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_nl), 8'b11111110, reg_chn_inp_in_crt_sva_6_94_64_reg,
      {(FpAdd_8U_23U_1_or_2_nl) , (FpAdd_8U_23U_1_and_19_nl) , (FpAdd_8U_23U_1_and_32_nl)
      , IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_4});
  assign FpAdd_8U_23U_1_and_2_tmp = FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_7_4_1 & reg_inp_lookup_3_FpMantRNE_49U_24U_1_else_and_svs_1_cse;
  assign FpAdd_8U_23U_1_if_4_FpAdd_8U_23U_1_if_4_or_6_nl = FpAdd_6U_10U_1_is_a_greater_lor_3_lpi_1_dfm_5
      | (~ FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_7_4_1);
  assign FpAdd_8U_23U_1_is_inf_3_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_1_is_a_greater_lor_3_lpi_1_dfm_5,
      (FpAdd_8U_23U_1_if_4_FpAdd_8U_23U_1_if_4_or_6_nl), reg_inp_lookup_3_FpMantRNE_49U_24U_1_else_and_svs_1_cse);
  assign FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_9_m1c = ~(IsNaN_8U_23U_3_land_3_lpi_1_dfm_7
      | IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_4);
  assign nl_FpAdd_6U_10U_1_int_mant_p1_3_sva = conv_u2u_23_24(FpAdd_6U_10U_1_addend_larger_qr_3_lpi_1_dfm_mx0)
      + conv_u2u_23_24(FpAdd_6U_10U_1_addend_smaller_qr_3_lpi_1_dfm_mx0);
  assign FpAdd_6U_10U_1_int_mant_p1_3_sva = nl_FpAdd_6U_10U_1_int_mant_p1_3_sva[23:0];
  assign FpAdd_6U_10U_1_addend_larger_qr_3_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_1_b_int_mant_p1_3_sva_2,
      reg_chn_inp_in_crt_sva_6_94_64_1_reg, FpAdd_6U_10U_1_is_a_greater_lor_3_lpi_1_dfm_5);
  assign FpAdd_6U_10U_1_addend_smaller_qr_3_lpi_1_dfm_mx0 = MUX_v_23_2_2(reg_chn_inp_in_crt_sva_6_94_64_1_reg,
      FpAdd_6U_10U_1_b_int_mant_p1_3_sva_2, FpAdd_6U_10U_1_is_a_greater_lor_3_lpi_1_dfm_5);
  assign nl_FpAdd_6U_10U_1_int_mant_p1_3_sva_1 = ({1'b1 , (~ FpAdd_6U_10U_1_addend_smaller_qr_3_lpi_1_dfm_mx0)})
      + conv_u2u_23_24(FpAdd_6U_10U_1_addend_larger_qr_3_lpi_1_dfm_mx0) + 24'b1;
  assign FpAdd_6U_10U_1_int_mant_p1_3_sva_1 = nl_FpAdd_6U_10U_1_int_mant_p1_3_sva_1[23:0];
  assign FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_mx0 = MUX_v_24_2_2(FpAdd_6U_10U_1_int_mant_p1_3_sva_1,
      FpAdd_6U_10U_1_int_mant_p1_3_sva, IsNaN_8U_23U_3_land_3_lpi_1_dfm_7);
  assign nl_inp_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_nl = FpAdd_8U_23U_1_o_expo_lpi_1_dfm_13
      + 8'b1;
  assign inp_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_nl = nl_inp_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_nl[7:0];
  assign FpAdd_8U_23U_1_or_3_nl = ((~(FpAdd_8U_23U_1_and_3_tmp | FpAdd_8U_23U_1_is_inf_lpi_1_dfm_2_mx0))
      & FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_11_m1c) | (IsNaN_8U_23U_3_land_lpi_1_dfm_6
      & (~ IsNaN_6U_10U_8_land_lpi_1_dfm_st_4));
  assign FpAdd_8U_23U_1_and_25_nl = FpAdd_8U_23U_1_and_3_tmp & (~ FpAdd_8U_23U_1_is_inf_lpi_1_dfm_2_mx0)
      & FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_11_m1c;
  assign FpAdd_8U_23U_1_and_34_nl = FpAdd_8U_23U_1_is_inf_lpi_1_dfm_2_mx0 & FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_11_m1c;
  assign FpAdd_8U_23U_1_o_expo_lpi_1_dfm_7 = MUX1HOT_v_8_4_2(FpAdd_8U_23U_1_o_expo_lpi_1_dfm_13,
      (inp_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_nl), 8'b11111110, reg_chn_inp_in_crt_sva_6_126_96_reg,
      {(FpAdd_8U_23U_1_or_3_nl) , (FpAdd_8U_23U_1_and_25_nl) , (FpAdd_8U_23U_1_and_34_nl)
      , IsNaN_6U_10U_8_land_lpi_1_dfm_st_4});
  assign FpAdd_8U_23U_1_and_3_tmp = FpMul_6U_10U_1_o_expo_lpi_1_dfm_7_4_1 & inp_lookup_4_FpMantRNE_49U_24U_1_else_and_svs_2;
  assign FpAdd_8U_23U_1_if_4_FpAdd_8U_23U_1_if_4_or_7_nl = FpAdd_6U_10U_1_is_a_greater_lor_lpi_1_dfm_5
      | (~ FpMul_6U_10U_1_o_expo_lpi_1_dfm_7_4_1);
  assign FpAdd_8U_23U_1_is_inf_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_1_is_a_greater_lor_lpi_1_dfm_5,
      (FpAdd_8U_23U_1_if_4_FpAdd_8U_23U_1_if_4_or_7_nl), inp_lookup_4_FpMantRNE_49U_24U_1_else_and_svs_2);
  assign FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_11_m1c = ~(IsNaN_8U_23U_3_land_lpi_1_dfm_6
      | IsNaN_6U_10U_8_land_lpi_1_dfm_st_4);
  assign nl_FpAdd_6U_10U_1_int_mant_p1_sva = conv_u2u_23_24(FpAdd_6U_10U_1_addend_larger_qr_lpi_1_dfm_mx0)
      + conv_u2u_23_24(FpAdd_6U_10U_1_addend_smaller_qr_lpi_1_dfm_mx0);
  assign FpAdd_6U_10U_1_int_mant_p1_sva = nl_FpAdd_6U_10U_1_int_mant_p1_sva[23:0];
  assign FpAdd_6U_10U_1_addend_larger_qr_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_1_b_int_mant_p1_sva_2,
      reg_chn_inp_in_crt_sva_6_126_96_1_reg, FpAdd_6U_10U_1_is_a_greater_lor_lpi_1_dfm_5);
  assign FpAdd_6U_10U_1_addend_smaller_qr_lpi_1_dfm_mx0 = MUX_v_23_2_2(reg_chn_inp_in_crt_sva_6_126_96_1_reg,
      FpAdd_6U_10U_1_b_int_mant_p1_sva_2, FpAdd_6U_10U_1_is_a_greater_lor_lpi_1_dfm_5);
  assign nl_FpAdd_6U_10U_1_int_mant_p1_sva_1 = ({1'b1 , (~ FpAdd_6U_10U_1_addend_smaller_qr_lpi_1_dfm_mx0)})
      + conv_u2u_23_24(FpAdd_6U_10U_1_addend_larger_qr_lpi_1_dfm_mx0) + 24'b1;
  assign FpAdd_6U_10U_1_int_mant_p1_sva_1 = nl_FpAdd_6U_10U_1_int_mant_p1_sva_1[23:0];
  assign FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_mx0 = MUX_v_24_2_2(FpAdd_6U_10U_1_int_mant_p1_sva_1,
      FpAdd_6U_10U_1_int_mant_p1_sva, IsNaN_8U_23U_3_land_lpi_1_dfm_6);
  assign inp_lookup_1_FpMantDecShiftRight_23U_8U_10U_carry_and_nl = ((FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_1_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_guard_mask_1_sva[23])) & ((FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_1_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_1_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_mask_1_sva[23]));
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_1_sva = (inp_lookup_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_itm[23:13])
      + conv_u2u_1_11(inp_lookup_1_FpMantDecShiftRight_23U_8U_10U_carry_and_nl);
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_1_sva = nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_1_sva[10:0];
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_1_lpi_1_dfm_3 = ~((~((FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_sva_3==6'b111111)
      & inp_lookup_1_FpMantRNE_24U_11U_else_and_svs_2 & inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_2
      & (~ inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2)))
      & inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_nor_ssc =
      ~(FpWidthDec_8U_23U_6U_10U_0U_1U_else_and_tmp | FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_1_lpi_1_dfm_3);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_and_1_m1c = FpWidthDec_8U_23U_6U_10U_0U_1U_else_and_tmp
      & (~ FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_1_lpi_1_dfm_3);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_and_tmp = inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_2
      & (~ inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2);
  assign nl_FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_sva_3 = ({(~ (FpAdd_6U_10U_1_qr_2_lpi_1_dfm_5[5]))
      , (FpAdd_6U_10U_1_qr_2_lpi_1_dfm_5[4:0])}) + 6'b1;
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_sva_3 = nl_FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_sva_3[5:0];
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_1_sva = FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_6
      & (FpMantDecShiftRight_23U_8U_10U_guard_mask_1_sva[22:0]);
  assign nl_inp_lookup_1_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl = (FpMantDecShiftRight_23U_8U_10U_guard_mask_1_sva[22:0])
      + 23'b11111111111111111111111;
  assign inp_lookup_1_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl = nl_inp_lookup_1_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_1_sva = FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_6
      & (inp_lookup_1_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl);
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_1_sva = FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_6
      & (FpMantDecShiftRight_23U_8U_10U_least_mask_1_sva[22:0]);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_1_lpi_1_dfm_2 = ((~((FpMantDecShiftRight_23U_8U_10U_o_mant_sum_1_sva[10])
      | inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_2))
      | inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2)
      & inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2;
  assign nl_FpAdd_6U_10U_1_o_expo_1_sva_1 = FpAdd_6U_10U_1_qr_2_lpi_1_dfm_5 + 6'b1;
  assign FpAdd_6U_10U_1_o_expo_1_sva_1 = nl_FpAdd_6U_10U_1_o_expo_1_sva_1[5:0];
  assign nl_inp_lookup_1_FpAdd_6U_10U_1_if_3_if_acc_1_nl = ({1'b1 , (FpAdd_6U_10U_1_qr_2_lpi_1_dfm_5[5:1])})
      + 6'b1;
  assign inp_lookup_1_FpAdd_6U_10U_1_if_3_if_acc_1_nl = nl_inp_lookup_1_FpAdd_6U_10U_1_if_3_if_acc_1_nl[5:0];
  assign inp_lookup_1_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((inp_lookup_1_FpAdd_6U_10U_1_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      inp_lookup_1_FpNormalize_6U_23U_1_else_lshift_itm, FpNormalize_6U_23U_1_oelse_not_9);
  assign nl_inp_lookup_1_FpNormalize_6U_23U_1_else_acc_nl = FpAdd_6U_10U_1_qr_2_lpi_1_dfm_5
      + ({1'b1 , (~ libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_8)})
      + 6'b1;
  assign inp_lookup_1_FpNormalize_6U_23U_1_else_acc_nl = nl_inp_lookup_1_FpNormalize_6U_23U_1_else_acc_nl[5:0];
  assign FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000, (inp_lookup_1_FpNormalize_6U_23U_1_else_acc_nl),
      FpNormalize_6U_23U_1_oelse_not_9);
  assign FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_5 = MUX1HOT_s_1_3_2((FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_1[5]),
      (FpAdd_6U_10U_1_qr_2_lpi_1_dfm_5[5]), (FpAdd_6U_10U_1_o_expo_1_sva_1[5]), {(~
      (FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_4[23])) , FpAdd_6U_10U_1_and_4_ssc
      , FpAdd_6U_10U_1_asn_124});
  assign FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_4 = MUX1HOT_s_1_3_2((FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_1[4]),
      (FpAdd_6U_10U_1_qr_2_lpi_1_dfm_5[4]), (FpAdd_6U_10U_1_o_expo_1_sva_1[4]), {(~
      (FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_4[23])) , FpAdd_6U_10U_1_and_4_ssc
      , FpAdd_6U_10U_1_asn_124});
  assign FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_3_0 = MUX1HOT_v_4_3_2((FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_1[3:0]),
      (FpAdd_6U_10U_1_qr_2_lpi_1_dfm_5[3:0]), (FpAdd_6U_10U_1_o_expo_1_sva_1[3:0]),
      {(~ (FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_4[23])) , FpAdd_6U_10U_1_and_4_ssc
      , FpAdd_6U_10U_1_asn_124});
  assign inp_lookup_1_FpMantRNE_23U_11U_1_else_and_tmp = FpMantRNE_23U_11U_1_else_carry_1_sva
      & (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_4[23]));
  assign FpMantRNE_23U_11U_1_else_carry_1_sva = (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_1_int_mant_2_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_4[22:1]), FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_4[23]);
  assign FpAdd_6U_10U_1_and_4_ssc = (~ inp_lookup_1_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1)
      & (FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_4[23]);
  assign inp_lookup_2_FpMantDecShiftRight_23U_8U_10U_carry_and_nl = ((FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_2_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_guard_mask_2_sva[23])) & ((FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_2_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_2_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_mask_2_sva[23]));
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_2_sva = (inp_lookup_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_itm[23:13])
      + conv_u2u_1_11(inp_lookup_2_FpMantDecShiftRight_23U_8U_10U_carry_and_nl);
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_2_sva = nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_2_sva[10:0];
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_2_lpi_1_dfm_3 = ~((~((FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_sva_3==6'b111111)
      & inp_lookup_2_FpMantRNE_24U_11U_else_and_svs_2 & IsNaN_6U_10U_9_land_2_lpi_1_dfm_8
      & (~ inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2)))
      & inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_nor_1_ssc
      = ~(FpWidthDec_8U_23U_6U_10U_0U_1U_else_and_1_tmp | FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_2_lpi_1_dfm_3);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_and_3_m1c = FpWidthDec_8U_23U_6U_10U_0U_1U_else_and_1_tmp
      & (~ FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_2_lpi_1_dfm_3);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_and_1_tmp = IsNaN_6U_10U_9_land_2_lpi_1_dfm_8
      & (~ inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2);
  assign nl_FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_sva_3 = ({(~ (FpAdd_6U_10U_1_qr_3_lpi_1_dfm_5[5]))
      , (FpAdd_6U_10U_1_qr_3_lpi_1_dfm_5[4:0])}) + 6'b1;
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_sva_3 = nl_FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_sva_3[5:0];
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_2_sva = FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_6
      & (FpMantDecShiftRight_23U_8U_10U_guard_mask_2_sva[22:0]);
  assign nl_inp_lookup_2_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl = (FpMantDecShiftRight_23U_8U_10U_guard_mask_2_sva[22:0])
      + 23'b11111111111111111111111;
  assign inp_lookup_2_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl = nl_inp_lookup_2_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_2_sva = FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_6
      & (inp_lookup_2_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl);
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_2_sva = FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_6
      & (FpMantDecShiftRight_23U_8U_10U_least_mask_2_sva[22:0]);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_2_lpi_1_dfm_5_mx0 = MUX_v_10_2_2(FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_1_mx0w1,
      (FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_6[9:0]), IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_5);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_2_lpi_1_dfm_2 = ((~((FpMantDecShiftRight_23U_8U_10U_o_mant_sum_2_sva[10])
      | IsNaN_6U_10U_9_land_2_lpi_1_dfm_8)) | inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2)
      & inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2;
  assign nl_FpAdd_6U_10U_1_o_expo_2_sva_1 = FpAdd_6U_10U_1_qr_3_lpi_1_dfm_5 + 6'b1;
  assign FpAdd_6U_10U_1_o_expo_2_sva_1 = nl_FpAdd_6U_10U_1_o_expo_2_sva_1[5:0];
  assign nl_inp_lookup_2_FpAdd_6U_10U_1_if_3_if_acc_1_nl = ({1'b1 , (FpAdd_6U_10U_1_qr_3_lpi_1_dfm_5[5:1])})
      + 6'b1;
  assign inp_lookup_2_FpAdd_6U_10U_1_if_3_if_acc_1_nl = nl_inp_lookup_2_FpAdd_6U_10U_1_if_3_if_acc_1_nl[5:0];
  assign inp_lookup_2_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((inp_lookup_2_FpAdd_6U_10U_1_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      inp_lookup_2_FpNormalize_6U_23U_1_else_lshift_itm, FpNormalize_6U_23U_1_oelse_not_11);
  assign nl_inp_lookup_2_FpNormalize_6U_23U_1_else_acc_nl = FpAdd_6U_10U_1_qr_3_lpi_1_dfm_5
      + ({1'b1 , (~ libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_9)})
      + 6'b1;
  assign inp_lookup_2_FpNormalize_6U_23U_1_else_acc_nl = nl_inp_lookup_2_FpNormalize_6U_23U_1_else_acc_nl[5:0];
  assign FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000, (inp_lookup_2_FpNormalize_6U_23U_1_else_acc_nl),
      FpNormalize_6U_23U_1_oelse_not_11);
  assign FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_5 = MUX1HOT_s_1_3_2((FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_1[5]),
      (FpAdd_6U_10U_1_qr_3_lpi_1_dfm_5[5]), (FpAdd_6U_10U_1_o_expo_2_sva_1[5]), {(~
      (FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_4[23])) , FpAdd_6U_10U_1_and_10_ssc
      , FpAdd_6U_10U_1_asn_126});
  assign FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_4 = MUX1HOT_s_1_3_2((FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_1[4]),
      (FpAdd_6U_10U_1_qr_3_lpi_1_dfm_5[4]), (FpAdd_6U_10U_1_o_expo_2_sva_1[4]), {(~
      (FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_4[23])) , FpAdd_6U_10U_1_and_10_ssc
      , FpAdd_6U_10U_1_asn_126});
  assign FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_3_0 = MUX1HOT_v_4_3_2((FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_1[3:0]),
      (FpAdd_6U_10U_1_qr_3_lpi_1_dfm_5[3:0]), (FpAdd_6U_10U_1_o_expo_2_sva_1[3:0]),
      {(~ (FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_4[23])) , FpAdd_6U_10U_1_and_10_ssc
      , FpAdd_6U_10U_1_asn_126});
  assign inp_lookup_2_FpMantRNE_23U_11U_1_else_and_tmp = FpMantRNE_23U_11U_1_else_carry_2_sva
      & (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_4[23]));
  assign FpMantRNE_23U_11U_1_else_carry_2_sva = (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_1_int_mant_3_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_4[22:1]), FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_4[23]);
  assign FpAdd_6U_10U_1_and_10_ssc = (~ inp_lookup_2_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1)
      & (FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_4[23]);
  assign inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_carry_and_nl = ((FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_3_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_guard_mask_3_sva[23])) & ((FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_3_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_3_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_mask_3_sva[23]));
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_3_sva = (inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_itm[23:13])
      + conv_u2u_1_11(inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_carry_and_nl);
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_3_sva = nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_3_sva[10:0];
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_3_lpi_1_dfm_3 = ~((~((FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_sva_3==6'b111111)
      & inp_lookup_3_FpMantRNE_24U_11U_else_and_svs_2 & IsNaN_6U_10U_9_land_3_lpi_1_dfm_8
      & (~ inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2)))
      & inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_nor_2_ssc
      = ~(FpWidthDec_8U_23U_6U_10U_0U_1U_else_and_2_tmp | FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_3_lpi_1_dfm_3);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_and_5_m1c = FpWidthDec_8U_23U_6U_10U_0U_1U_else_and_2_tmp
      & (~ FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_3_lpi_1_dfm_3);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_and_2_tmp = IsNaN_6U_10U_9_land_3_lpi_1_dfm_8
      & (~ inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2);
  assign nl_FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_sva_3 = ({(~ (FpAdd_6U_10U_1_qr_4_lpi_1_dfm_5[5]))
      , (FpAdd_6U_10U_1_qr_4_lpi_1_dfm_5[4:0])}) + 6'b1;
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_sva_3 = nl_FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_sva_3[5:0];
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_3_sva = FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_6
      & (FpMantDecShiftRight_23U_8U_10U_guard_mask_3_sva[22:0]);
  assign nl_inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl = (FpMantDecShiftRight_23U_8U_10U_guard_mask_3_sva[22:0])
      + 23'b11111111111111111111111;
  assign inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl = nl_inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_3_sva = FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_6
      & (inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl);
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_3_sva = FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_6
      & (FpMantDecShiftRight_23U_8U_10U_least_mask_3_sva[22:0]);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_3_lpi_1_dfm_5_mx0 = MUX_v_10_2_2(FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_2_mx0w1,
      (FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_6[9:0]), IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_5);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_3_lpi_1_dfm_2 = ((~((FpMantDecShiftRight_23U_8U_10U_o_mant_sum_3_sva[10])
      | IsNaN_6U_10U_9_land_3_lpi_1_dfm_8)) | inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2)
      & inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2;
  assign nl_FpAdd_6U_10U_1_o_expo_3_sva_1 = FpAdd_6U_10U_1_qr_4_lpi_1_dfm_5 + 6'b1;
  assign FpAdd_6U_10U_1_o_expo_3_sva_1 = nl_FpAdd_6U_10U_1_o_expo_3_sva_1[5:0];
  assign nl_inp_lookup_3_FpAdd_6U_10U_1_if_3_if_acc_1_nl = ({1'b1 , (FpAdd_6U_10U_1_qr_4_lpi_1_dfm_5[5:1])})
      + 6'b1;
  assign inp_lookup_3_FpAdd_6U_10U_1_if_3_if_acc_1_nl = nl_inp_lookup_3_FpAdd_6U_10U_1_if_3_if_acc_1_nl[5:0];
  assign inp_lookup_3_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((inp_lookup_3_FpAdd_6U_10U_1_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      inp_lookup_3_FpNormalize_6U_23U_1_else_lshift_itm, FpNormalize_6U_23U_1_oelse_not_13);
  assign nl_inp_lookup_3_FpNormalize_6U_23U_1_else_acc_nl = FpAdd_6U_10U_1_qr_4_lpi_1_dfm_5
      + ({1'b1 , (~ libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_10)})
      + 6'b1;
  assign inp_lookup_3_FpNormalize_6U_23U_1_else_acc_nl = nl_inp_lookup_3_FpNormalize_6U_23U_1_else_acc_nl[5:0];
  assign FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000, (inp_lookup_3_FpNormalize_6U_23U_1_else_acc_nl),
      FpNormalize_6U_23U_1_oelse_not_13);
  assign FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_5 = MUX1HOT_s_1_3_2((FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_1[5]),
      (FpAdd_6U_10U_1_qr_4_lpi_1_dfm_5[5]), (FpAdd_6U_10U_1_o_expo_3_sva_1[5]), {(~
      (FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_4[23])) , FpAdd_6U_10U_1_and_16_ssc
      , FpAdd_6U_10U_1_asn_128});
  assign FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_4 = MUX1HOT_s_1_3_2((FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_1[4]),
      (FpAdd_6U_10U_1_qr_4_lpi_1_dfm_5[4]), (FpAdd_6U_10U_1_o_expo_3_sva_1[4]), {(~
      (FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_4[23])) , FpAdd_6U_10U_1_and_16_ssc
      , FpAdd_6U_10U_1_asn_128});
  assign FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_3_0 = MUX1HOT_v_4_3_2((FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_1[3:0]),
      (FpAdd_6U_10U_1_qr_4_lpi_1_dfm_5[3:0]), (FpAdd_6U_10U_1_o_expo_3_sva_1[3:0]),
      {(~ (FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_4[23])) , FpAdd_6U_10U_1_and_16_ssc
      , FpAdd_6U_10U_1_asn_128});
  assign inp_lookup_3_FpMantRNE_23U_11U_1_else_and_tmp = FpMantRNE_23U_11U_1_else_carry_3_sva
      & (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_4[23]));
  assign FpMantRNE_23U_11U_1_else_carry_3_sva = (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_1_int_mant_4_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_4[22:1]), FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_4[23]);
  assign FpAdd_6U_10U_1_and_16_ssc = (~ inp_lookup_3_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1)
      & (FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_4[23]);
  assign inp_lookup_4_FpMantDecShiftRight_23U_8U_10U_carry_and_nl = ((FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_guard_mask_sva[23])) & ((FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_mask_sva[23]));
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva = (inp_lookup_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_itm[23:13])
      + conv_u2u_1_11(inp_lookup_4_FpMantDecShiftRight_23U_8U_10U_carry_and_nl);
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva = nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva[10:0];
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_lpi_1_dfm_3 = ~((~((FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_sva_3==6'b111111)
      & inp_lookup_4_FpMantRNE_24U_11U_else_and_svs_2 & IsNaN_6U_10U_9_land_lpi_1_dfm_8
      & (~ inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2)))
      & inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_FpWidthDec_8U_23U_6U_10U_0U_1U_nor_3_ssc
      = ~(FpWidthDec_8U_23U_6U_10U_0U_1U_else_and_3_tmp | FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_lpi_1_dfm_3);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_and_7_m1c = FpWidthDec_8U_23U_6U_10U_0U_1U_else_and_3_tmp
      & (~ FpWidthDec_8U_23U_6U_10U_0U_1U_is_inf_lpi_1_dfm_3);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_else_and_3_tmp = IsNaN_6U_10U_9_land_lpi_1_dfm_8
      & (~ inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2);
  assign nl_FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_sva_3 = ({(~ (FpAdd_6U_10U_1_qr_lpi_1_dfm_5[5]))
      , (FpAdd_6U_10U_1_qr_lpi_1_dfm_5[4:0])}) + 6'b1;
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_sva_3 = nl_FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_sva_3[5:0];
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_sva = FpAdd_8U_23U_1_o_mant_lpi_1_dfm_6
      & (FpMantDecShiftRight_23U_8U_10U_guard_mask_sva[22:0]);
  assign nl_inp_lookup_4_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl = (FpMantDecShiftRight_23U_8U_10U_guard_mask_sva[22:0])
      + 23'b11111111111111111111111;
  assign inp_lookup_4_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl = nl_inp_lookup_4_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_sva = FpAdd_8U_23U_1_o_mant_lpi_1_dfm_6
      & (inp_lookup_4_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl);
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_sva = FpAdd_8U_23U_1_o_mant_lpi_1_dfm_6
      & (FpMantDecShiftRight_23U_8U_10U_least_mask_sva[22:0]);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_lpi_1_dfm_5_mx0 = MUX_v_10_2_2(FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_3_mx0w1,
      (FpAdd_8U_23U_1_o_mant_lpi_1_dfm_6[9:0]), IsNaN_6U_10U_8_land_lpi_1_dfm_st_5);
  assign FpWidthDec_8U_23U_6U_10U_0U_1U_is_zero_lpi_1_dfm_2 = ((~((FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva[10])
      | IsNaN_6U_10U_9_land_lpi_1_dfm_8)) | inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2)
      & inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2;
  assign nl_FpAdd_6U_10U_1_o_expo_sva_1 = FpAdd_6U_10U_1_qr_lpi_1_dfm_5 + 6'b1;
  assign FpAdd_6U_10U_1_o_expo_sva_1 = nl_FpAdd_6U_10U_1_o_expo_sva_1[5:0];
  assign nl_inp_lookup_4_FpAdd_6U_10U_1_if_3_if_acc_1_nl = ({1'b1 , (FpAdd_6U_10U_1_qr_lpi_1_dfm_5[5:1])})
      + 6'b1;
  assign inp_lookup_4_FpAdd_6U_10U_1_if_3_if_acc_1_nl = nl_inp_lookup_4_FpAdd_6U_10U_1_if_3_if_acc_1_nl[5:0];
  assign inp_lookup_4_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((inp_lookup_4_FpAdd_6U_10U_1_if_3_if_acc_1_nl));
  assign FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      inp_lookup_4_FpNormalize_6U_23U_1_else_lshift_itm, FpNormalize_6U_23U_1_oelse_not_15);
  assign nl_inp_lookup_4_FpNormalize_6U_23U_1_else_acc_nl = FpAdd_6U_10U_1_qr_lpi_1_dfm_5
      + ({1'b1 , (~ libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_11)})
      + 6'b1;
  assign inp_lookup_4_FpNormalize_6U_23U_1_else_acc_nl = nl_inp_lookup_4_FpNormalize_6U_23U_1_else_acc_nl[5:0];
  assign FpAdd_6U_10U_1_o_expo_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000, (inp_lookup_4_FpNormalize_6U_23U_1_else_acc_nl),
      FpNormalize_6U_23U_1_oelse_not_15);
  assign FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_5 = MUX1HOT_s_1_3_2((FpAdd_6U_10U_1_o_expo_lpi_1_dfm_1[5]),
      (FpAdd_6U_10U_1_qr_lpi_1_dfm_5[5]), (FpAdd_6U_10U_1_o_expo_sva_1[5]), {(~ (FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_4[23]))
      , FpAdd_6U_10U_1_and_22_ssc , FpAdd_6U_10U_1_asn_130});
  assign FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_4 = MUX1HOT_s_1_3_2((FpAdd_6U_10U_1_o_expo_lpi_1_dfm_1[4]),
      (FpAdd_6U_10U_1_qr_lpi_1_dfm_5[4]), (FpAdd_6U_10U_1_o_expo_sva_1[4]), {(~ (FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_4[23]))
      , FpAdd_6U_10U_1_and_22_ssc , FpAdd_6U_10U_1_asn_130});
  assign FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_3_0 = MUX1HOT_v_4_3_2((FpAdd_6U_10U_1_o_expo_lpi_1_dfm_1[3:0]),
      (FpAdd_6U_10U_1_qr_lpi_1_dfm_5[3:0]), (FpAdd_6U_10U_1_o_expo_sva_1[3:0]), {(~
      (FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_4[23])) , FpAdd_6U_10U_1_and_22_ssc ,
      FpAdd_6U_10U_1_asn_130});
  assign inp_lookup_4_FpMantRNE_23U_11U_1_else_and_tmp = FpMantRNE_23U_11U_1_else_carry_sva
      & (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) &
      ((FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_1[22]) | (FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_4[23]));
  assign FpMantRNE_23U_11U_1_else_carry_sva = (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_1_int_mant_1_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_4[22:1]), FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_4[23]);
  assign FpAdd_6U_10U_1_and_22_ssc = (~ inp_lookup_4_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1)
      & (FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_4[23]);
  assign nl_inp_lookup_1_FpMul_6U_10U_oelse_1_acc_nl = conv_s2s_7_8(FpMul_6U_10U_oelse_1_acc_itm_2)
      + conv_u2s_6_8({FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_10_5_1 ,
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_10_4_0_1});
  assign inp_lookup_1_FpMul_6U_10U_oelse_1_acc_nl = nl_inp_lookup_1_FpMul_6U_10U_oelse_1_acc_nl[7:0];
  assign inp_lookup_1_FpMul_6U_10U_oelse_1_acc_itm_7_1 = readslicef_8_1_7((inp_lookup_1_FpMul_6U_10U_oelse_1_acc_nl));
  assign FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_9_0_1_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_itm_2, IsNaN_6U_23U_2_land_1_lpi_1_dfm);
  assign IsNaN_6U_23U_2_land_1_lpi_1_dfm = ~((~((FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_itm_2!=10'b0000000000)))
      | IsNaN_6U_10U_land_1_lpi_1_dfm_5);
  assign nl_inp_lookup_2_FpMul_6U_10U_oelse_1_acc_nl = conv_s2s_7_8(FpMul_6U_10U_oelse_1_acc_1_itm_2)
      + conv_u2s_6_8({FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_10_5_1 ,
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_10_4_0_1});
  assign inp_lookup_2_FpMul_6U_10U_oelse_1_acc_nl = nl_inp_lookup_2_FpMul_6U_10U_oelse_1_acc_nl[7:0];
  assign inp_lookup_2_FpMul_6U_10U_oelse_1_acc_itm_7_1 = readslicef_8_1_7((inp_lookup_2_FpMul_6U_10U_oelse_1_acc_nl));
  assign FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_9_0_2_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_1_itm_2, IsNaN_6U_23U_2_land_2_lpi_1_dfm);
  assign IsNaN_6U_23U_2_land_2_lpi_1_dfm = ~((~((FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_1_itm_2!=10'b0000000000)))
      | IsNaN_6U_10U_land_2_lpi_1_dfm_5);
  assign nl_inp_lookup_3_FpMul_6U_10U_oelse_1_acc_nl = conv_s2s_7_8(FpMul_6U_10U_oelse_1_acc_2_itm_2)
      + conv_u2s_6_8({FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_10_5_1 ,
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_10_4_0_1});
  assign inp_lookup_3_FpMul_6U_10U_oelse_1_acc_nl = nl_inp_lookup_3_FpMul_6U_10U_oelse_1_acc_nl[7:0];
  assign inp_lookup_3_FpMul_6U_10U_oelse_1_acc_itm_7_1 = readslicef_8_1_7((inp_lookup_3_FpMul_6U_10U_oelse_1_acc_nl));
  assign FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_9_0_3_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_2_itm_2, IsNaN_6U_23U_2_land_3_lpi_1_dfm);
  assign IsNaN_6U_23U_2_land_3_lpi_1_dfm = ~((~((FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_2_itm_2!=10'b0000000000)))
      | IsNaN_6U_10U_land_3_lpi_1_dfm_5);
  assign nl_inp_lookup_4_FpMul_6U_10U_oelse_1_acc_nl = conv_s2s_7_8(FpMul_6U_10U_oelse_1_acc_3_itm_2)
      + conv_u2s_6_8({FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_10_5_1 , FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_10_4_0_1});
  assign inp_lookup_4_FpMul_6U_10U_oelse_1_acc_nl = nl_inp_lookup_4_FpMul_6U_10U_oelse_1_acc_nl[7:0];
  assign inp_lookup_4_FpMul_6U_10U_oelse_1_acc_itm_7_1 = readslicef_8_1_7((inp_lookup_4_FpMul_6U_10U_oelse_1_acc_nl));
  assign FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_9_0_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_3_itm_2, IsNaN_6U_23U_2_land_lpi_1_dfm);
  assign IsNaN_6U_23U_2_land_lpi_1_dfm = ~((~((FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_3_itm_2!=10'b0000000000)))
      | IsNaN_6U_10U_land_lpi_1_dfm_5);
  assign nl_inp_lookup_1_FpMul_6U_10U_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_6U_10U_else_2_else_ac_int_cctor_1_sva_2[5:1])})
      + 6'b1;
  assign inp_lookup_1_FpMul_6U_10U_else_2_else_if_if_acc_1_nl = nl_inp_lookup_1_FpMul_6U_10U_else_2_else_if_if_acc_1_nl[5:0];
  assign inp_lookup_1_FpMul_6U_10U_else_2_else_if_if_acc_1_itm_5_1 = readslicef_6_1_5((inp_lookup_1_FpMul_6U_10U_else_2_else_if_if_acc_1_nl));
  assign inp_lookup_1_FpMantRNE_22U_11U_else_and_svs = FpMantRNE_22U_11U_else_carry_1_sva
      & (FpMul_6U_10U_p_mant_20_1_1_lpi_1_dfm_3_mx0[19:10]==10'b1111111111);
  assign FpMantRNE_22U_11U_else_carry_1_sva = (FpMul_6U_10U_p_mant_20_1_1_lpi_1_dfm_3_mx0[9])
      & (((FpMul_6U_10U_p_mant_p1_1_sva_2[0]) & (FpMul_6U_10U_p_mant_p1_1_sva_2[21]))
      | (FpMul_6U_10U_p_mant_20_1_1_lpi_1_dfm_3_mx0[0]) | (FpMul_6U_10U_p_mant_20_1_1_lpi_1_dfm_3_mx0[1])
      | (FpMul_6U_10U_p_mant_20_1_1_lpi_1_dfm_3_mx0[2]) | (FpMul_6U_10U_p_mant_20_1_1_lpi_1_dfm_3_mx0[3])
      | (FpMul_6U_10U_p_mant_20_1_1_lpi_1_dfm_3_mx0[4]) | (FpMul_6U_10U_p_mant_20_1_1_lpi_1_dfm_3_mx0[5])
      | (FpMul_6U_10U_p_mant_20_1_1_lpi_1_dfm_3_mx0[6]) | (FpMul_6U_10U_p_mant_20_1_1_lpi_1_dfm_3_mx0[7])
      | (FpMul_6U_10U_p_mant_20_1_1_lpi_1_dfm_3_mx0[8]) | (FpMul_6U_10U_p_mant_20_1_1_lpi_1_dfm_3_mx0[10]));
  assign FpMul_6U_10U_p_mant_20_1_1_lpi_1_dfm_3_mx0 = MUX_v_20_2_2((FpMul_6U_10U_p_mant_p1_1_sva_2[19:0]),
      (FpMul_6U_10U_p_mant_p1_1_sva_2[20:1]), FpMul_6U_10U_p_mant_p1_1_sva_2[21]);
  assign nl_inp_lookup_2_FpMul_6U_10U_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_6U_10U_else_2_else_ac_int_cctor_2_sva_2[5:1])})
      + 6'b1;
  assign inp_lookup_2_FpMul_6U_10U_else_2_else_if_if_acc_1_nl = nl_inp_lookup_2_FpMul_6U_10U_else_2_else_if_if_acc_1_nl[5:0];
  assign inp_lookup_2_FpMul_6U_10U_else_2_else_if_if_acc_1_itm_5_1 = readslicef_6_1_5((inp_lookup_2_FpMul_6U_10U_else_2_else_if_if_acc_1_nl));
  assign inp_lookup_2_FpMantRNE_22U_11U_else_and_svs = FpMantRNE_22U_11U_else_carry_2_sva
      & (FpMul_6U_10U_p_mant_20_1_2_lpi_1_dfm_3_mx0[19:10]==10'b1111111111);
  assign FpMantRNE_22U_11U_else_carry_2_sva = (FpMul_6U_10U_p_mant_20_1_2_lpi_1_dfm_3_mx0[9])
      & (((FpMul_6U_10U_p_mant_p1_2_sva_2[0]) & (FpMul_6U_10U_p_mant_p1_2_sva_2[21]))
      | (FpMul_6U_10U_p_mant_20_1_2_lpi_1_dfm_3_mx0[0]) | (FpMul_6U_10U_p_mant_20_1_2_lpi_1_dfm_3_mx0[1])
      | (FpMul_6U_10U_p_mant_20_1_2_lpi_1_dfm_3_mx0[2]) | (FpMul_6U_10U_p_mant_20_1_2_lpi_1_dfm_3_mx0[3])
      | (FpMul_6U_10U_p_mant_20_1_2_lpi_1_dfm_3_mx0[4]) | (FpMul_6U_10U_p_mant_20_1_2_lpi_1_dfm_3_mx0[5])
      | (FpMul_6U_10U_p_mant_20_1_2_lpi_1_dfm_3_mx0[6]) | (FpMul_6U_10U_p_mant_20_1_2_lpi_1_dfm_3_mx0[7])
      | (FpMul_6U_10U_p_mant_20_1_2_lpi_1_dfm_3_mx0[8]) | (FpMul_6U_10U_p_mant_20_1_2_lpi_1_dfm_3_mx0[10]));
  assign FpMul_6U_10U_p_mant_20_1_2_lpi_1_dfm_3_mx0 = MUX_v_20_2_2((FpMul_6U_10U_p_mant_p1_2_sva_2[19:0]),
      (FpMul_6U_10U_p_mant_p1_2_sva_2[20:1]), FpMul_6U_10U_p_mant_p1_2_sva_2[21]);
  assign nl_inp_lookup_3_FpMul_6U_10U_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_6U_10U_else_2_else_ac_int_cctor_3_sva_2[5:1])})
      + 6'b1;
  assign inp_lookup_3_FpMul_6U_10U_else_2_else_if_if_acc_1_nl = nl_inp_lookup_3_FpMul_6U_10U_else_2_else_if_if_acc_1_nl[5:0];
  assign inp_lookup_3_FpMul_6U_10U_else_2_else_if_if_acc_1_itm_5_1 = readslicef_6_1_5((inp_lookup_3_FpMul_6U_10U_else_2_else_if_if_acc_1_nl));
  assign inp_lookup_3_FpMantRNE_22U_11U_else_and_svs = FpMantRNE_22U_11U_else_carry_3_sva
      & (FpMul_6U_10U_p_mant_20_1_3_lpi_1_dfm_3_mx0[19:10]==10'b1111111111);
  assign FpMantRNE_22U_11U_else_carry_3_sva = (FpMul_6U_10U_p_mant_20_1_3_lpi_1_dfm_3_mx0[9])
      & (((FpMul_6U_10U_p_mant_p1_3_sva_2[0]) & (FpMul_6U_10U_p_mant_p1_3_sva_2[21]))
      | (FpMul_6U_10U_p_mant_20_1_3_lpi_1_dfm_3_mx0[0]) | (FpMul_6U_10U_p_mant_20_1_3_lpi_1_dfm_3_mx0[1])
      | (FpMul_6U_10U_p_mant_20_1_3_lpi_1_dfm_3_mx0[2]) | (FpMul_6U_10U_p_mant_20_1_3_lpi_1_dfm_3_mx0[3])
      | (FpMul_6U_10U_p_mant_20_1_3_lpi_1_dfm_3_mx0[4]) | (FpMul_6U_10U_p_mant_20_1_3_lpi_1_dfm_3_mx0[5])
      | (FpMul_6U_10U_p_mant_20_1_3_lpi_1_dfm_3_mx0[6]) | (FpMul_6U_10U_p_mant_20_1_3_lpi_1_dfm_3_mx0[7])
      | (FpMul_6U_10U_p_mant_20_1_3_lpi_1_dfm_3_mx0[8]) | (FpMul_6U_10U_p_mant_20_1_3_lpi_1_dfm_3_mx0[10]));
  assign FpMul_6U_10U_p_mant_20_1_3_lpi_1_dfm_3_mx0 = MUX_v_20_2_2((FpMul_6U_10U_p_mant_p1_3_sva_2[19:0]),
      (FpMul_6U_10U_p_mant_p1_3_sva_2[20:1]), FpMul_6U_10U_p_mant_p1_3_sva_2[21]);
  assign nl_inp_lookup_4_FpMul_6U_10U_else_2_else_if_if_acc_1_nl = ({1'b1 , (FpMul_6U_10U_else_2_else_ac_int_cctor_sva_2[5:1])})
      + 6'b1;
  assign inp_lookup_4_FpMul_6U_10U_else_2_else_if_if_acc_1_nl = nl_inp_lookup_4_FpMul_6U_10U_else_2_else_if_if_acc_1_nl[5:0];
  assign inp_lookup_4_FpMul_6U_10U_else_2_else_if_if_acc_1_itm_5_1 = readslicef_6_1_5((inp_lookup_4_FpMul_6U_10U_else_2_else_if_if_acc_1_nl));
  assign inp_lookup_4_FpMantRNE_22U_11U_else_and_svs = FpMantRNE_22U_11U_else_carry_sva
      & (FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0[19:10]==10'b1111111111);
  assign FpMantRNE_22U_11U_else_carry_sva = (FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0[9])
      & (((FpMul_6U_10U_p_mant_p1_sva_2[0]) & (FpMul_6U_10U_p_mant_p1_sva_2[21]))
      | (FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0[0]) | (FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0[1])
      | (FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0[2]) | (FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0[3])
      | (FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0[4]) | (FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0[5])
      | (FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0[6]) | (FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0[7])
      | (FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0[8]) | (FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0[10]));
  assign FpMul_6U_10U_p_mant_20_1_lpi_1_dfm_3_mx0 = MUX_v_20_2_2((FpMul_6U_10U_p_mant_p1_sva_2[19:0]),
      (FpMul_6U_10U_p_mant_p1_sva_2[20:1]), FpMul_6U_10U_p_mant_p1_sva_2[21]);
  assign nl_FpAdd_6U_10U_int_mant_p1_1_sva = conv_u2u_23_24(FpAdd_6U_10U_addend_larger_qr_1_lpi_1_dfm_mx0)
      + conv_u2u_23_24(FpAdd_6U_10U_addend_smaller_qr_1_lpi_1_dfm_mx0);
  assign FpAdd_6U_10U_int_mant_p1_1_sva = nl_FpAdd_6U_10U_int_mant_p1_1_sva[23:0];
  assign FpAdd_6U_10U_addend_larger_qr_1_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_b_int_mant_p1_1_sva_2,
      FpAdd_6U_10U_a_int_mant_p1_1_sva_2, FpAdd_6U_10U_is_a_greater_lor_1_lpi_1_dfm_5);
  assign FpAdd_6U_10U_addend_smaller_qr_1_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_a_int_mant_p1_1_sva_2,
      FpAdd_6U_10U_b_int_mant_p1_1_sva_2, FpAdd_6U_10U_is_a_greater_lor_1_lpi_1_dfm_5);
  assign FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_mx0 = MUX_v_24_2_2(FpAdd_6U_10U_asn_23_mx0w1,
      FpAdd_6U_10U_int_mant_p1_1_sva, reg_inp_lookup_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse);
  assign nl_FpAdd_6U_10U_int_mant_p1_2_sva = conv_u2u_23_24(FpAdd_6U_10U_addend_larger_qr_2_lpi_1_dfm_mx0)
      + conv_u2u_23_24(FpAdd_6U_10U_addend_smaller_qr_2_lpi_1_dfm_mx0);
  assign FpAdd_6U_10U_int_mant_p1_2_sva = nl_FpAdd_6U_10U_int_mant_p1_2_sva[23:0];
  assign FpAdd_6U_10U_addend_larger_qr_2_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_b_int_mant_p1_2_sva_2,
      FpAdd_6U_10U_a_int_mant_p1_2_sva_2, FpAdd_6U_10U_is_a_greater_lor_2_lpi_1_dfm_5);
  assign FpAdd_6U_10U_addend_smaller_qr_2_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_a_int_mant_p1_2_sva_2,
      FpAdd_6U_10U_b_int_mant_p1_2_sva_2, FpAdd_6U_10U_is_a_greater_lor_2_lpi_1_dfm_5);
  assign FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_mx0 = MUX_v_24_2_2(FpAdd_6U_10U_asn_20_mx0w1,
      FpAdd_6U_10U_int_mant_p1_2_sva, reg_inp_lookup_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse);
  assign nl_FpAdd_6U_10U_int_mant_p1_3_sva = conv_u2u_23_24(FpAdd_6U_10U_addend_larger_qr_3_lpi_1_dfm_mx0)
      + conv_u2u_23_24(FpAdd_6U_10U_addend_smaller_qr_3_lpi_1_dfm_mx0);
  assign FpAdd_6U_10U_int_mant_p1_3_sva = nl_FpAdd_6U_10U_int_mant_p1_3_sva[23:0];
  assign FpAdd_6U_10U_addend_larger_qr_3_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_b_int_mant_p1_3_sva_2,
      FpAdd_6U_10U_a_int_mant_p1_3_sva_2, FpAdd_6U_10U_is_a_greater_lor_3_lpi_1_dfm_5);
  assign FpAdd_6U_10U_addend_smaller_qr_3_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_a_int_mant_p1_3_sva_2,
      FpAdd_6U_10U_b_int_mant_p1_3_sva_2, FpAdd_6U_10U_is_a_greater_lor_3_lpi_1_dfm_5);
  assign FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_mx0 = MUX_v_24_2_2(FpAdd_6U_10U_asn_17_mx0w1,
      FpAdd_6U_10U_int_mant_p1_3_sva, reg_inp_lookup_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse);
  assign nl_FpAdd_6U_10U_int_mant_p1_sva = conv_u2u_23_24(FpAdd_6U_10U_addend_larger_qr_lpi_1_dfm_mx0)
      + conv_u2u_23_24(FpAdd_6U_10U_addend_smaller_qr_lpi_1_dfm_mx0);
  assign FpAdd_6U_10U_int_mant_p1_sva = nl_FpAdd_6U_10U_int_mant_p1_sva[23:0];
  assign FpAdd_6U_10U_addend_larger_qr_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_b_int_mant_p1_sva_2,
      FpAdd_6U_10U_a_int_mant_p1_sva_2, FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_5);
  assign FpAdd_6U_10U_addend_smaller_qr_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_a_int_mant_p1_sva_2,
      FpAdd_6U_10U_b_int_mant_p1_sva_2, FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_5);
  assign FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_mx0 = MUX_v_24_2_2(FpAdd_6U_10U_asn_mx0w1,
      FpAdd_6U_10U_int_mant_p1_sva, reg_inp_lookup_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse);
  assign or_5860_nl = (~ IsInf_6U_23U_land_1_lpi_1_dfm_mx0w0) | IsNaN_6U_23U_IsNaN_6U_23U_nor_tmp;
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_o_mant_9_0_1_lpi_1_dfm_2_mx0 = MUX_v_10_2_2(({{9{IsInf_6U_23U_land_1_lpi_1_dfm_mx0w0}},
      IsInf_6U_23U_land_1_lpi_1_dfm_mx0w0}), FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_9_0_1_lpi_1_dfm,
      or_5860_nl);
  assign IsNaN_6U_23U_aelse_not_8_nl = ~ IsNaN_6U_23U_IsNaN_6U_23U_nor_tmp;
  assign FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_22_13_1_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      FpAdd_6U_10U_o_mant_1_lpi_1_dfm_2_mx0, (IsNaN_6U_23U_aelse_not_8_nl));
  assign nl_FpAdd_6U_10U_o_expo_1_sva_1 = ({reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_4_5_4_tmp
      , reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_4_5_4_tmp_1 , FpAdd_6U_10U_qr_2_lpi_1_dfm_4_3_0_1})
      + 6'b1;
  assign FpAdd_6U_10U_o_expo_1_sva_1 = nl_FpAdd_6U_10U_o_expo_1_sva_1[5:0];
  assign FpNormalize_6U_23U_oelse_not_16_nl = ~ reg_FpNormalize_6U_23U_lor_1_lpi_1_dfm_4_cse;
  assign FpAdd_6U_10U_int_mant_2_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      inp_lookup_1_FpNormalize_6U_23U_else_lshift_itm, (FpNormalize_6U_23U_oelse_not_16_nl));
  assign nl_inp_lookup_1_FpNormalize_6U_23U_else_acc_nl = ({reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_4_5_4_tmp
      , reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_4_5_4_tmp_1 , FpAdd_6U_10U_qr_2_lpi_1_dfm_4_3_0_1})
      + ({1'b1 , (~ IntLeadZero_23U_leading_sign_23_0_rtn_1_sva_2)}) + 6'b1;
  assign inp_lookup_1_FpNormalize_6U_23U_else_acc_nl = nl_inp_lookup_1_FpNormalize_6U_23U_else_acc_nl[5:0];
  assign FpNormalize_6U_23U_oelse_not_8_nl = ~ reg_FpNormalize_6U_23U_lor_1_lpi_1_dfm_4_cse;
  assign FpAdd_6U_10U_o_expo_1_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000, (inp_lookup_1_FpNormalize_6U_23U_else_acc_nl),
      (FpNormalize_6U_23U_oelse_not_8_nl));
  assign nl_FpAdd_6U_10U_o_expo_1_sva_4 = ({FpAdd_6U_10U_o_expo_1_lpi_1_dfm_2_5_4
      , FpAdd_6U_10U_o_expo_1_lpi_1_dfm_2_3_0}) + 6'b1;
  assign FpAdd_6U_10U_o_expo_1_sva_4 = nl_FpAdd_6U_10U_o_expo_1_sva_4[5:0];
  assign FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_int_mant_2_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_4[22:1]), FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_4[23]);
  assign FpMantRNE_23U_11U_else_carry_1_sva = (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_nl = FpAdd_6U_10U_and_4_ssc | (~
      inp_lookup_1_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_is_inf_1_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_and_4_ssc,
      (FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_nl), inp_lookup_1_FpMantRNE_23U_11U_else_and_tmp);
  assign nl_inp_lookup_1_FpAdd_6U_10U_if_4_if_acc_1_nl = ({1'b1 , FpAdd_6U_10U_o_expo_1_lpi_1_dfm_2_5_4
      , (FpAdd_6U_10U_o_expo_1_lpi_1_dfm_2_3_0[3:1])}) + 6'b1;
  assign inp_lookup_1_FpAdd_6U_10U_if_4_if_acc_1_nl = nl_inp_lookup_1_FpAdd_6U_10U_if_4_if_acc_1_nl[5:0];
  assign inp_lookup_1_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((inp_lookup_1_FpAdd_6U_10U_if_4_if_acc_1_nl));
  assign FpAdd_6U_10U_o_expo_1_lpi_1_dfm_2_5_4 = MUX1HOT_v_2_3_2((FpAdd_6U_10U_o_expo_1_lpi_1_dfm_1[5:4]),
      ({reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_4_5_4_tmp , reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_4_5_4_tmp_1}),
      (FpAdd_6U_10U_o_expo_1_sva_1[5:4]), {(~ (FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_4[23]))
      , FpAdd_6U_10U_and_4_ssc , FpAdd_6U_10U_asn_87});
  assign FpAdd_6U_10U_o_expo_1_lpi_1_dfm_2_3_0 = MUX1HOT_v_4_3_2((FpAdd_6U_10U_o_expo_1_lpi_1_dfm_1[3:0]),
      FpAdd_6U_10U_qr_2_lpi_1_dfm_4_3_0_1, (FpAdd_6U_10U_o_expo_1_sva_1[3:0]), {(~
      (FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_4[23])) , FpAdd_6U_10U_and_4_ssc , FpAdd_6U_10U_asn_87});
  assign FpAdd_6U_10U_and_4_ssc = (~ FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_1_sva_2)
      & (FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_4[23]);
  assign FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_9_0_1_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      FpAdd_6U_10U_o_mant_1_lpi_1_dfm_2_mx0, IsNaN_6U_23U_IsNaN_6U_23U_nor_tmp);
  assign FpAdd_6U_10U_o_expo_1_lpi_1_dfm_7_3_0 = MUX1HOT_v_4_4_2(FpAdd_6U_10U_o_expo_1_lpi_1_dfm_2_3_0,
      (FpAdd_6U_10U_o_expo_1_sva_4[3:0]), 4'b1110, FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_29,
      {FpAdd_6U_10U_and_ssc , FpAdd_6U_10U_and_6_ssc , FpAdd_6U_10U_and_28_ssc ,
      FpAdd_6U_10U_or_16_cse});
  assign IsNaN_6U_23U_IsNaN_6U_23U_nand_cse = ~((FpAdd_6U_10U_o_expo_1_lpi_1_dfm_7_5_4==2'b11)
      & (FpAdd_6U_10U_o_expo_1_lpi_1_dfm_7_3_0==4'b1111));
  assign nl_inp_lookup_1_FpMantRNE_23U_11U_else_acc_nl = (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_else_carry_1_sva);
  assign inp_lookup_1_FpMantRNE_23U_11U_else_acc_nl = nl_inp_lookup_1_FpMantRNE_23U_11U_else_acc_nl[9:0];
  assign FpAdd_6U_10U_FpAdd_6U_10U_or_4_nl = MUX_v_10_2_2((inp_lookup_1_FpMantRNE_23U_11U_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_is_inf_1_lpi_1_dfm_2_mx0);
  assign FpAdd_6U_10U_o_mant_1_lpi_1_dfm_2_mx0 = MUX_v_10_2_2((FpAdd_6U_10U_FpAdd_6U_10U_or_4_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_26, FpAdd_6U_10U_or_16_cse);
  assign FpAdd_6U_10U_and_ssc = (~(FpAdd_6U_10U_and_tmp | FpAdd_6U_10U_is_inf_1_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_FpAdd_6U_10U_nor_5_m1c;
  assign FpAdd_6U_10U_and_6_ssc = FpAdd_6U_10U_and_tmp & (~ FpAdd_6U_10U_is_inf_1_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_FpAdd_6U_10U_nor_5_m1c;
  assign FpAdd_6U_10U_and_28_ssc = FpAdd_6U_10U_is_inf_1_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_FpAdd_6U_10U_nor_5_m1c;
  assign FpAdd_6U_10U_FpAdd_6U_10U_nor_5_m1c = ~(IsNaN_6U_10U_3_land_1_lpi_1_dfm_8
      | IsNaN_6U_10U_2_land_1_lpi_1_dfm_26);
  assign FpAdd_6U_10U_and_tmp = inp_lookup_1_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1 &
      inp_lookup_1_FpMantRNE_23U_11U_else_and_tmp;
  assign inp_lookup_1_FpMantRNE_23U_11U_else_and_tmp = FpMantRNE_23U_11U_else_carry_1_sva
      & (FpAdd_6U_10U_int_mant_2_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) & ((FpAdd_6U_10U_int_mant_2_lpi_1_dfm_1[22])
      | (FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_4[23]));
  assign or_5861_nl = (~ IsInf_6U_23U_land_2_lpi_1_dfm_mx0w0) | IsNaN_6U_23U_IsNaN_6U_23U_nor_1_tmp;
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_o_mant_9_0_2_lpi_1_dfm_2_mx0 = MUX_v_10_2_2(({{9{IsInf_6U_23U_land_2_lpi_1_dfm_mx0w0}},
      IsInf_6U_23U_land_2_lpi_1_dfm_mx0w0}), FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_9_0_2_lpi_1_dfm,
      or_5861_nl);
  assign IsNaN_6U_23U_aelse_not_9_nl = ~ IsNaN_6U_23U_IsNaN_6U_23U_nor_1_tmp;
  assign FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_22_13_2_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      FpAdd_6U_10U_o_mant_2_lpi_1_dfm_2_mx0, (IsNaN_6U_23U_aelse_not_9_nl));
  assign nl_FpAdd_6U_10U_o_expo_2_sva_1 = ({reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_4_5_4_tmp
      , reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_4_5_4_tmp_1 , FpAdd_6U_10U_qr_3_lpi_1_dfm_4_3_0_1})
      + 6'b1;
  assign FpAdd_6U_10U_o_expo_2_sva_1 = nl_FpAdd_6U_10U_o_expo_2_sva_1[5:0];
  assign FpNormalize_6U_23U_oelse_not_17_nl = ~ reg_FpNormalize_6U_23U_lor_2_lpi_1_dfm_4_cse;
  assign FpAdd_6U_10U_int_mant_3_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      inp_lookup_2_FpNormalize_6U_23U_else_lshift_itm, (FpNormalize_6U_23U_oelse_not_17_nl));
  assign nl_inp_lookup_2_FpNormalize_6U_23U_else_acc_nl = ({reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_4_5_4_tmp
      , reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_4_5_4_tmp_1 , FpAdd_6U_10U_qr_3_lpi_1_dfm_4_3_0_1})
      + ({1'b1 , (~ IntLeadZero_23U_leading_sign_23_0_rtn_2_sva_2)}) + 6'b1;
  assign inp_lookup_2_FpNormalize_6U_23U_else_acc_nl = nl_inp_lookup_2_FpNormalize_6U_23U_else_acc_nl[5:0];
  assign FpNormalize_6U_23U_oelse_not_10_nl = ~ reg_FpNormalize_6U_23U_lor_2_lpi_1_dfm_4_cse;
  assign FpAdd_6U_10U_o_expo_2_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000, (inp_lookup_2_FpNormalize_6U_23U_else_acc_nl),
      (FpNormalize_6U_23U_oelse_not_10_nl));
  assign nl_FpAdd_6U_10U_o_expo_2_sva_4 = ({FpAdd_6U_10U_o_expo_2_lpi_1_dfm_2_5_4
      , FpAdd_6U_10U_o_expo_2_lpi_1_dfm_2_3_0}) + 6'b1;
  assign FpAdd_6U_10U_o_expo_2_sva_4 = nl_FpAdd_6U_10U_o_expo_2_sva_4[5:0];
  assign FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_int_mant_3_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_4[22:1]), FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_4[23]);
  assign FpMantRNE_23U_11U_else_carry_2_sva = (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_1_nl = FpAdd_6U_10U_and_10_ssc |
      (~ inp_lookup_2_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_is_inf_2_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_and_10_ssc,
      (FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_1_nl), inp_lookup_2_FpMantRNE_23U_11U_else_and_tmp);
  assign nl_inp_lookup_2_FpAdd_6U_10U_if_4_if_acc_1_nl = ({1'b1 , FpAdd_6U_10U_o_expo_2_lpi_1_dfm_2_5_4
      , (FpAdd_6U_10U_o_expo_2_lpi_1_dfm_2_3_0[3:1])}) + 6'b1;
  assign inp_lookup_2_FpAdd_6U_10U_if_4_if_acc_1_nl = nl_inp_lookup_2_FpAdd_6U_10U_if_4_if_acc_1_nl[5:0];
  assign inp_lookup_2_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((inp_lookup_2_FpAdd_6U_10U_if_4_if_acc_1_nl));
  assign FpAdd_6U_10U_o_expo_2_lpi_1_dfm_2_5_4 = MUX1HOT_v_2_3_2((FpAdd_6U_10U_o_expo_2_lpi_1_dfm_1[5:4]),
      ({reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_4_5_4_tmp , reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_4_5_4_tmp_1}),
      (FpAdd_6U_10U_o_expo_2_sva_1[5:4]), {(~ (FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_4[23]))
      , FpAdd_6U_10U_and_10_ssc , FpAdd_6U_10U_asn_89});
  assign FpAdd_6U_10U_o_expo_2_lpi_1_dfm_2_3_0 = MUX1HOT_v_4_3_2((FpAdd_6U_10U_o_expo_2_lpi_1_dfm_1[3:0]),
      FpAdd_6U_10U_qr_3_lpi_1_dfm_4_3_0_1, (FpAdd_6U_10U_o_expo_2_sva_1[3:0]), {(~
      (FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_4[23])) , FpAdd_6U_10U_and_10_ssc , FpAdd_6U_10U_asn_89});
  assign FpAdd_6U_10U_and_10_ssc = (~ FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_2_sva_2)
      & (FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_4[23]);
  assign FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_9_0_2_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      FpAdd_6U_10U_o_mant_2_lpi_1_dfm_2_mx0, IsNaN_6U_23U_IsNaN_6U_23U_nor_1_tmp);
  assign FpAdd_6U_10U_o_expo_2_lpi_1_dfm_7_3_0 = MUX1HOT_v_4_4_2(FpAdd_6U_10U_o_expo_2_lpi_1_dfm_2_3_0,
      (FpAdd_6U_10U_o_expo_2_sva_4[3:0]), 4'b1110, FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_29,
      {FpAdd_6U_10U_and_29_ssc , FpAdd_6U_10U_and_13_ssc , FpAdd_6U_10U_and_30_ssc
      , FpAdd_6U_10U_or_17_cse});
  assign IsNaN_6U_23U_IsNaN_6U_23U_nand_1_cse = ~((FpAdd_6U_10U_o_expo_2_lpi_1_dfm_7_5_4==2'b11)
      & (FpAdd_6U_10U_o_expo_2_lpi_1_dfm_7_3_0==4'b1111));
  assign nl_inp_lookup_2_FpMantRNE_23U_11U_else_acc_nl = (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_else_carry_2_sva);
  assign inp_lookup_2_FpMantRNE_23U_11U_else_acc_nl = nl_inp_lookup_2_FpMantRNE_23U_11U_else_acc_nl[9:0];
  assign FpAdd_6U_10U_FpAdd_6U_10U_or_6_nl = MUX_v_10_2_2((inp_lookup_2_FpMantRNE_23U_11U_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_is_inf_2_lpi_1_dfm_2_mx0);
  assign FpAdd_6U_10U_o_mant_2_lpi_1_dfm_2_mx0 = MUX_v_10_2_2((FpAdd_6U_10U_FpAdd_6U_10U_or_6_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_26, FpAdd_6U_10U_or_17_cse);
  assign FpAdd_6U_10U_and_29_ssc = (~(FpAdd_6U_10U_and_1_tmp | FpAdd_6U_10U_is_inf_2_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_FpAdd_6U_10U_nor_7_m1c;
  assign FpAdd_6U_10U_and_13_ssc = FpAdd_6U_10U_and_1_tmp & (~ FpAdd_6U_10U_is_inf_2_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_FpAdd_6U_10U_nor_7_m1c;
  assign FpAdd_6U_10U_and_30_ssc = FpAdd_6U_10U_is_inf_2_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_FpAdd_6U_10U_nor_7_m1c;
  assign FpAdd_6U_10U_FpAdd_6U_10U_nor_7_m1c = ~(IsNaN_6U_10U_3_land_2_lpi_1_dfm_8
      | IsNaN_6U_10U_2_land_2_lpi_1_dfm_26);
  assign FpAdd_6U_10U_and_1_tmp = inp_lookup_2_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1
      & inp_lookup_2_FpMantRNE_23U_11U_else_and_tmp;
  assign inp_lookup_2_FpMantRNE_23U_11U_else_and_tmp = FpMantRNE_23U_11U_else_carry_2_sva
      & (FpAdd_6U_10U_int_mant_3_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) & ((FpAdd_6U_10U_int_mant_3_lpi_1_dfm_1[22])
      | (FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_4[23]));
  assign or_5862_nl = (~ IsInf_6U_23U_land_3_lpi_1_dfm_mx0w0) | IsNaN_6U_23U_IsNaN_6U_23U_nor_2_tmp;
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_o_mant_9_0_3_lpi_1_dfm_2_mx0 = MUX_v_10_2_2(({{9{IsInf_6U_23U_land_3_lpi_1_dfm_mx0w0}},
      IsInf_6U_23U_land_3_lpi_1_dfm_mx0w0}), FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_9_0_3_lpi_1_dfm,
      or_5862_nl);
  assign IsNaN_6U_23U_aelse_not_10_nl = ~ IsNaN_6U_23U_IsNaN_6U_23U_nor_2_tmp;
  assign FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_22_13_3_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      FpAdd_6U_10U_o_mant_3_lpi_1_dfm_2_mx0, (IsNaN_6U_23U_aelse_not_10_nl));
  assign nl_FpAdd_6U_10U_o_expo_3_sva_1 = ({reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_4_5_4_tmp
      , reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_4_5_4_tmp_1 , FpAdd_6U_10U_qr_4_lpi_1_dfm_4_3_0_1})
      + 6'b1;
  assign FpAdd_6U_10U_o_expo_3_sva_1 = nl_FpAdd_6U_10U_o_expo_3_sva_1[5:0];
  assign FpNormalize_6U_23U_oelse_not_18_nl = ~ FpNormalize_6U_23U_lor_3_lpi_1_dfm_5;
  assign FpAdd_6U_10U_int_mant_4_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      inp_lookup_3_FpNormalize_6U_23U_else_lshift_itm, (FpNormalize_6U_23U_oelse_not_18_nl));
  assign nl_inp_lookup_3_FpNormalize_6U_23U_else_acc_nl = ({reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_4_5_4_tmp
      , reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_4_5_4_tmp_1 , FpAdd_6U_10U_qr_4_lpi_1_dfm_4_3_0_1})
      + ({1'b1 , (~ IntLeadZero_23U_leading_sign_23_0_rtn_3_sva_2)}) + 6'b1;
  assign inp_lookup_3_FpNormalize_6U_23U_else_acc_nl = nl_inp_lookup_3_FpNormalize_6U_23U_else_acc_nl[5:0];
  assign FpNormalize_6U_23U_oelse_not_12_nl = ~ FpNormalize_6U_23U_lor_3_lpi_1_dfm_5;
  assign FpAdd_6U_10U_o_expo_3_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000, (inp_lookup_3_FpNormalize_6U_23U_else_acc_nl),
      (FpNormalize_6U_23U_oelse_not_12_nl));
  assign nl_FpAdd_6U_10U_o_expo_3_sva_4 = ({FpAdd_6U_10U_o_expo_3_lpi_1_dfm_2_5_4
      , FpAdd_6U_10U_o_expo_3_lpi_1_dfm_2_3_0}) + 6'b1;
  assign FpAdd_6U_10U_o_expo_3_sva_4 = nl_FpAdd_6U_10U_o_expo_3_sva_4[5:0];
  assign FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_int_mant_4_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_4[22:1]), FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_4[23]);
  assign FpMantRNE_23U_11U_else_carry_3_sva = (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_2_nl = FpAdd_6U_10U_and_16_ssc |
      (~ inp_lookup_3_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_is_inf_3_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_and_16_ssc,
      (FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_2_nl), inp_lookup_3_FpMantRNE_23U_11U_else_and_tmp);
  assign nl_inp_lookup_3_FpAdd_6U_10U_if_4_if_acc_1_nl = ({1'b1 , FpAdd_6U_10U_o_expo_3_lpi_1_dfm_2_5_4
      , (FpAdd_6U_10U_o_expo_3_lpi_1_dfm_2_3_0[3:1])}) + 6'b1;
  assign inp_lookup_3_FpAdd_6U_10U_if_4_if_acc_1_nl = nl_inp_lookup_3_FpAdd_6U_10U_if_4_if_acc_1_nl[5:0];
  assign inp_lookup_3_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((inp_lookup_3_FpAdd_6U_10U_if_4_if_acc_1_nl));
  assign FpAdd_6U_10U_o_expo_3_lpi_1_dfm_2_5_4 = MUX1HOT_v_2_3_2((FpAdd_6U_10U_o_expo_3_lpi_1_dfm_1[5:4]),
      ({reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_4_5_4_tmp , reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_4_5_4_tmp_1}),
      (FpAdd_6U_10U_o_expo_3_sva_1[5:4]), {(~ (FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_4[23]))
      , FpAdd_6U_10U_and_16_ssc , FpAdd_6U_10U_asn_91});
  assign FpAdd_6U_10U_o_expo_3_lpi_1_dfm_2_3_0 = MUX1HOT_v_4_3_2((FpAdd_6U_10U_o_expo_3_lpi_1_dfm_1[3:0]),
      FpAdd_6U_10U_qr_4_lpi_1_dfm_4_3_0_1, (FpAdd_6U_10U_o_expo_3_sva_1[3:0]), {(~
      (FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_4[23])) , FpAdd_6U_10U_and_16_ssc , FpAdd_6U_10U_asn_91});
  assign FpAdd_6U_10U_and_16_ssc = (~ FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_3_sva_2)
      & (FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_4[23]);
  assign FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_9_0_3_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      FpAdd_6U_10U_o_mant_3_lpi_1_dfm_2_mx0, IsNaN_6U_23U_IsNaN_6U_23U_nor_2_tmp);
  assign FpAdd_6U_10U_o_expo_3_lpi_1_dfm_7_3_0 = MUX1HOT_v_4_4_2(FpAdd_6U_10U_o_expo_3_lpi_1_dfm_2_3_0,
      (FpAdd_6U_10U_o_expo_3_sva_4[3:0]), 4'b1110, FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_29,
      {FpAdd_6U_10U_and_31_ssc , FpAdd_6U_10U_and_19_ssc , FpAdd_6U_10U_and_32_ssc
      , FpAdd_6U_10U_or_18_cse});
  assign IsNaN_6U_23U_IsNaN_6U_23U_nand_2_cse = ~((FpAdd_6U_10U_o_expo_3_lpi_1_dfm_7_5_4==2'b11)
      & (FpAdd_6U_10U_o_expo_3_lpi_1_dfm_7_3_0==4'b1111));
  assign nl_inp_lookup_3_FpMantRNE_23U_11U_else_acc_nl = (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_else_carry_3_sva);
  assign inp_lookup_3_FpMantRNE_23U_11U_else_acc_nl = nl_inp_lookup_3_FpMantRNE_23U_11U_else_acc_nl[9:0];
  assign FpAdd_6U_10U_FpAdd_6U_10U_or_8_nl = MUX_v_10_2_2((inp_lookup_3_FpMantRNE_23U_11U_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_is_inf_3_lpi_1_dfm_2_mx0);
  assign FpAdd_6U_10U_o_mant_3_lpi_1_dfm_2_mx0 = MUX_v_10_2_2((FpAdd_6U_10U_FpAdd_6U_10U_or_8_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_29, FpAdd_6U_10U_or_18_cse);
  assign FpAdd_6U_10U_and_31_ssc = (~(FpAdd_6U_10U_and_2_tmp | FpAdd_6U_10U_is_inf_3_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_FpAdd_6U_10U_nor_9_m1c;
  assign FpAdd_6U_10U_and_19_ssc = FpAdd_6U_10U_and_2_tmp & (~ FpAdd_6U_10U_is_inf_3_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_FpAdd_6U_10U_nor_9_m1c;
  assign FpAdd_6U_10U_and_32_ssc = FpAdd_6U_10U_is_inf_3_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_FpAdd_6U_10U_nor_9_m1c;
  assign FpAdd_6U_10U_FpAdd_6U_10U_nor_9_m1c = ~(IsNaN_6U_10U_3_land_3_lpi_1_dfm_8
      | IsNaN_6U_10U_2_land_3_lpi_1_dfm_26);
  assign FpAdd_6U_10U_and_2_tmp = inp_lookup_3_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1
      & inp_lookup_3_FpMantRNE_23U_11U_else_and_tmp;
  assign inp_lookup_3_FpMantRNE_23U_11U_else_and_tmp = FpMantRNE_23U_11U_else_carry_3_sva
      & (FpAdd_6U_10U_int_mant_4_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) & ((FpAdd_6U_10U_int_mant_4_lpi_1_dfm_1[22])
      | (FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_4[23]));
  assign or_5863_nl = (~ IsInf_6U_23U_land_lpi_1_dfm_mx0w0) | IsNaN_6U_23U_IsNaN_6U_23U_nor_3_tmp;
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_o_mant_9_0_lpi_1_dfm_2_mx0 = MUX_v_10_2_2(({{9{IsInf_6U_23U_land_lpi_1_dfm_mx0w0}},
      IsInf_6U_23U_land_lpi_1_dfm_mx0w0}), FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_9_0_lpi_1_dfm,
      or_5863_nl);
  assign IsNaN_6U_23U_aelse_not_11_nl = ~ IsNaN_6U_23U_IsNaN_6U_23U_nor_3_tmp;
  assign FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_22_13_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      FpAdd_6U_10U_o_mant_lpi_1_dfm_2_mx0, (IsNaN_6U_23U_aelse_not_11_nl));
  assign nl_FpAdd_6U_10U_o_expo_sva_1 = ({reg_FpAdd_6U_10U_qr_lpi_1_dfm_4_5_4_tmp
      , reg_FpAdd_6U_10U_qr_lpi_1_dfm_4_5_4_tmp_1 , FpAdd_6U_10U_qr_lpi_1_dfm_4_3_0_1})
      + 6'b1;
  assign FpAdd_6U_10U_o_expo_sva_1 = nl_FpAdd_6U_10U_o_expo_sva_1[5:0];
  assign FpNormalize_6U_23U_oelse_not_19_nl = ~ reg_FpNormalize_6U_23U_lor_lpi_1_dfm_4_cse;
  assign FpAdd_6U_10U_int_mant_1_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      inp_lookup_4_FpNormalize_6U_23U_else_lshift_itm, (FpNormalize_6U_23U_oelse_not_19_nl));
  assign nl_inp_lookup_4_FpNormalize_6U_23U_else_acc_nl = ({reg_FpAdd_6U_10U_qr_lpi_1_dfm_4_5_4_tmp
      , reg_FpAdd_6U_10U_qr_lpi_1_dfm_4_5_4_tmp_1 , FpAdd_6U_10U_qr_lpi_1_dfm_4_3_0_1})
      + ({1'b1 , (~ IntLeadZero_23U_leading_sign_23_0_rtn_sva_2)}) + 6'b1;
  assign inp_lookup_4_FpNormalize_6U_23U_else_acc_nl = nl_inp_lookup_4_FpNormalize_6U_23U_else_acc_nl[5:0];
  assign FpNormalize_6U_23U_oelse_not_14_nl = ~ reg_FpNormalize_6U_23U_lor_lpi_1_dfm_4_cse;
  assign FpAdd_6U_10U_o_expo_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000, (inp_lookup_4_FpNormalize_6U_23U_else_acc_nl),
      (FpNormalize_6U_23U_oelse_not_14_nl));
  assign nl_FpAdd_6U_10U_o_expo_sva_4 = ({FpAdd_6U_10U_o_expo_lpi_1_dfm_2_5_4 , FpAdd_6U_10U_o_expo_lpi_1_dfm_2_3_0})
      + 6'b1;
  assign FpAdd_6U_10U_o_expo_sva_4 = nl_FpAdd_6U_10U_o_expo_sva_4[5:0];
  assign FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_int_mant_1_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_4[22:1]), FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_4[23]);
  assign FpMantRNE_23U_11U_else_carry_sva = (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_3_nl = FpAdd_6U_10U_and_22_ssc |
      (~ inp_lookup_4_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_is_inf_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_and_22_ssc,
      (FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_3_nl), inp_lookup_4_FpMantRNE_23U_11U_else_and_tmp);
  assign nl_inp_lookup_4_FpAdd_6U_10U_if_4_if_acc_1_nl = ({1'b1 , FpAdd_6U_10U_o_expo_lpi_1_dfm_2_5_4
      , (FpAdd_6U_10U_o_expo_lpi_1_dfm_2_3_0[3:1])}) + 6'b1;
  assign inp_lookup_4_FpAdd_6U_10U_if_4_if_acc_1_nl = nl_inp_lookup_4_FpAdd_6U_10U_if_4_if_acc_1_nl[5:0];
  assign inp_lookup_4_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((inp_lookup_4_FpAdd_6U_10U_if_4_if_acc_1_nl));
  assign FpAdd_6U_10U_o_expo_lpi_1_dfm_2_5_4 = MUX1HOT_v_2_3_2((FpAdd_6U_10U_o_expo_lpi_1_dfm_1[5:4]),
      ({reg_FpAdd_6U_10U_qr_lpi_1_dfm_4_5_4_tmp , reg_FpAdd_6U_10U_qr_lpi_1_dfm_4_5_4_tmp_1}),
      (FpAdd_6U_10U_o_expo_sva_1[5:4]), {(~ (FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_4[23]))
      , FpAdd_6U_10U_and_22_ssc , FpAdd_6U_10U_asn_93});
  assign FpAdd_6U_10U_o_expo_lpi_1_dfm_2_3_0 = MUX1HOT_v_4_3_2((FpAdd_6U_10U_o_expo_lpi_1_dfm_1[3:0]),
      FpAdd_6U_10U_qr_lpi_1_dfm_4_3_0_1, (FpAdd_6U_10U_o_expo_sva_1[3:0]), {(~ (FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_4[23]))
      , FpAdd_6U_10U_and_22_ssc , FpAdd_6U_10U_asn_93});
  assign FpAdd_6U_10U_and_22_ssc = (~ FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_sva_2)
      & (FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_4[23]);
  assign FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_9_0_lpi_1_dfm = MUX_v_10_2_2(10'b0000000000,
      FpAdd_6U_10U_o_mant_lpi_1_dfm_2_mx0, IsNaN_6U_23U_IsNaN_6U_23U_nor_3_tmp);
  assign FpAdd_6U_10U_o_expo_lpi_1_dfm_7_3_0 = MUX1HOT_v_4_4_2(FpAdd_6U_10U_o_expo_lpi_1_dfm_2_3_0,
      (FpAdd_6U_10U_o_expo_sva_4[3:0]), 4'b1110, FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_29,
      {FpAdd_6U_10U_and_33_ssc , FpAdd_6U_10U_and_25_ssc , FpAdd_6U_10U_and_34_ssc
      , FpAdd_6U_10U_or_19_cse});
  assign IsNaN_6U_23U_IsNaN_6U_23U_nand_3_cse = ~((FpAdd_6U_10U_o_expo_lpi_1_dfm_7_5_4==2'b11)
      & (FpAdd_6U_10U_o_expo_lpi_1_dfm_7_3_0==4'b1111));
  assign nl_inp_lookup_4_FpMantRNE_23U_11U_else_acc_nl = (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[21:12])
      + conv_u2u_1_10(FpMantRNE_23U_11U_else_carry_sva);
  assign inp_lookup_4_FpMantRNE_23U_11U_else_acc_nl = nl_inp_lookup_4_FpMantRNE_23U_11U_else_acc_nl[9:0];
  assign FpAdd_6U_10U_FpAdd_6U_10U_or_10_nl = MUX_v_10_2_2((inp_lookup_4_FpMantRNE_23U_11U_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_is_inf_lpi_1_dfm_2_mx0);
  assign FpAdd_6U_10U_o_mant_lpi_1_dfm_2_mx0 = MUX_v_10_2_2((FpAdd_6U_10U_FpAdd_6U_10U_or_10_nl),
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_26, FpAdd_6U_10U_or_19_cse);
  assign FpAdd_6U_10U_and_33_ssc = (~(FpAdd_6U_10U_and_3_tmp | FpAdd_6U_10U_is_inf_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_FpAdd_6U_10U_nor_11_m1c;
  assign FpAdd_6U_10U_and_25_ssc = FpAdd_6U_10U_and_3_tmp & (~ FpAdd_6U_10U_is_inf_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_FpAdd_6U_10U_nor_11_m1c;
  assign FpAdd_6U_10U_and_34_ssc = FpAdd_6U_10U_is_inf_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_FpAdd_6U_10U_nor_11_m1c;
  assign FpAdd_6U_10U_FpAdd_6U_10U_nor_11_m1c = ~(IsNaN_6U_10U_3_land_lpi_1_dfm_8
      | IsNaN_6U_10U_2_land_lpi_1_dfm_26);
  assign FpAdd_6U_10U_and_3_tmp = inp_lookup_4_FpAdd_6U_10U_if_4_if_acc_1_itm_5_1
      & inp_lookup_4_FpMantRNE_23U_11U_else_and_tmp;
  assign inp_lookup_4_FpMantRNE_23U_11U_else_and_tmp = FpMantRNE_23U_11U_else_carry_sva
      & (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) & ((FpAdd_6U_10U_int_mant_1_lpi_1_dfm_1[22])
      | (FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_4[23]));
  assign inp_lookup_and_68_m1c = ~(inp_lookup_else_unequal_tmp_38 | (chn_inp_in_crt_sva_12_739_736_1[3]));
  assign inp_lookup_and_70_m1c = (~ inp_lookup_if_unequal_tmp_19) & (chn_inp_in_crt_sva_12_739_736_1[3]);
  assign inp_lookup_and_8_m1c = ~(inp_lookup_else_unequal_tmp_38 | (chn_inp_in_crt_sva_12_739_736_1[0]));
  assign inp_lookup_and_10_m1c = (~ inp_lookup_if_unequal_tmp_19) & (chn_inp_in_crt_sva_12_739_736_1[0]);
  assign inp_lookup_and_48_m1c = ~(inp_lookup_else_unequal_tmp_38 | (chn_inp_in_crt_sva_12_739_736_1[2]));
  assign inp_lookup_and_50_m1c = (~ inp_lookup_if_unequal_tmp_19) & (chn_inp_in_crt_sva_12_739_736_1[2]);
  assign inp_lookup_and_28_m1c = ~(inp_lookup_else_unequal_tmp_38 | (chn_inp_in_crt_sva_12_739_736_1[1]));
  assign inp_lookup_and_30_m1c = (~ inp_lookup_if_unequal_tmp_19) & (chn_inp_in_crt_sva_12_739_736_1[1]);
  assign main_stage_en_1 = chn_inp_in_rsci_bawt & or_11_cse;
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_1_sva = ({1'b1 , (~
      libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_16)}) + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_1_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_1_sva[4:0];
  assign IsZero_5U_10U_3_land_1_lpi_1_dfm = ~((chn_inp_in_rsci_d_mxwt[341:332]!=10'b0000000000)
      | (~ IsZero_5U_10U_3_IsZero_5U_10U_3_nor_cse_1_sva));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_cse
      = ~(IsDenorm_5U_10U_3_land_1_lpi_1_dfm | IsInf_5U_10U_3_land_1_lpi_1_dfm);
  assign IsInf_5U_10U_3_land_1_lpi_1_dfm = ~((chn_inp_in_rsci_d_mxwt[341:332]!=10'b0000000000)
      | (~ IsInf_5U_10U_3_IsInf_5U_10U_3_and_cse_1_sva));
  assign IsNaN_5U_10U_3_land_1_lpi_1_dfm = IsDenorm_5U_10U_3_or_tmp & IsInf_5U_10U_3_IsInf_5U_10U_3_and_cse_1_sva;
  assign IsInf_5U_10U_3_IsInf_5U_10U_3_and_cse_1_sva = (chn_inp_in_rsci_d_mxwt[346:342]==5'b11111);
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_2_sva = ({1'b1 , (~
      libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_17)}) + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_2_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_2_sva[4:0];
  assign IsZero_5U_10U_3_land_2_lpi_1_dfm = ~((chn_inp_in_rsci_d_mxwt[357:348]!=10'b0000000000)
      | (~ IsZero_5U_10U_3_IsZero_5U_10U_3_nor_cse_2_sva));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_1_cse
      = ~(IsDenorm_5U_10U_3_land_2_lpi_1_dfm | IsInf_5U_10U_3_land_2_lpi_1_dfm);
  assign IsInf_5U_10U_3_land_2_lpi_1_dfm = ~((chn_inp_in_rsci_d_mxwt[357:348]!=10'b0000000000)
      | (~ IsInf_5U_10U_3_IsInf_5U_10U_3_and_cse_2_sva));
  assign IsNaN_5U_10U_3_land_2_lpi_1_dfm = IsDenorm_5U_10U_3_or_1_tmp & IsInf_5U_10U_3_IsInf_5U_10U_3_and_cse_2_sva;
  assign IsInf_5U_10U_3_IsInf_5U_10U_3_and_cse_2_sva = (chn_inp_in_rsci_d_mxwt[362:358]==5'b11111);
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_3_sva = ({1'b1 , (~
      libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_18)}) + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_3_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_3_sva[4:0];
  assign IsZero_5U_10U_3_land_3_lpi_1_dfm = ~((chn_inp_in_rsci_d_mxwt[373:364]!=10'b0000000000)
      | (~ IsZero_5U_10U_3_IsZero_5U_10U_3_nor_cse_3_sva));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_2_cse
      = ~(IsDenorm_5U_10U_3_land_3_lpi_1_dfm | IsInf_5U_10U_3_land_3_lpi_1_dfm);
  assign IsInf_5U_10U_3_land_3_lpi_1_dfm = ~((chn_inp_in_rsci_d_mxwt[373:364]!=10'b0000000000)
      | (~ IsInf_5U_10U_3_IsInf_5U_10U_3_and_cse_3_sva));
  assign IsNaN_5U_10U_3_land_3_lpi_1_dfm = IsDenorm_5U_10U_3_or_2_tmp & IsInf_5U_10U_3_IsInf_5U_10U_3_and_cse_3_sva;
  assign IsInf_5U_10U_3_IsInf_5U_10U_3_and_cse_3_sva = (chn_inp_in_rsci_d_mxwt[378:374]==5'b11111);
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_sva = ({1'b1 , (~ libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_19)})
      + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_3_if_1_if_acc_psp_sva[4:0];
  assign IsZero_5U_10U_3_land_lpi_1_dfm = ~((chn_inp_in_rsci_d_mxwt[389:380]!=10'b0000000000)
      | (~ IsZero_5U_10U_3_IsZero_5U_10U_3_nor_cse_sva));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_nor_3_cse
      = ~(IsDenorm_5U_10U_3_land_lpi_1_dfm | IsInf_5U_10U_3_land_lpi_1_dfm);
  assign IsInf_5U_10U_3_land_lpi_1_dfm = ~((chn_inp_in_rsci_d_mxwt[389:380]!=10'b0000000000)
      | (~ IsInf_5U_10U_3_IsInf_5U_10U_3_and_cse_sva));
  assign IsNaN_5U_10U_3_land_lpi_1_dfm = IsDenorm_5U_10U_3_or_3_tmp & IsInf_5U_10U_3_IsInf_5U_10U_3_and_cse_sva;
  assign IsInf_5U_10U_3_IsInf_5U_10U_3_and_cse_sva = (chn_inp_in_rsci_d_mxwt[394:390]==5'b11111);
  assign FpAdd_8U_23U_b_right_shift_qr_1_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_4,
      FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_5);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_23_nl = ~ FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_5;
  assign FpAdd_8U_23U_a_right_shift_qr_1_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_4,
      (FpAdd_8U_23U_is_a_greater_oelse_not_23_nl));
  assign nl_FpMantRNE_36U_11U_else_ac_int_cctor_2_sva = (FpMantRNE_36U_11U_i_data_2_sva[35:25])
      + conv_u2u_1_11(FpMantRNE_36U_11U_else_carry_1_sva);
  assign FpMantRNE_36U_11U_else_ac_int_cctor_2_sva = nl_FpMantRNE_36U_11U_else_ac_int_cctor_2_sva[10:0];
  assign FpAdd_8U_23U_b_right_shift_qr_2_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_6,
      FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_5);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_25_nl = ~ FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_5;
  assign FpAdd_8U_23U_a_right_shift_qr_2_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_6,
      (FpAdd_8U_23U_is_a_greater_oelse_not_25_nl));
  assign nl_FpMantRNE_36U_11U_else_ac_int_cctor_3_sva = (FpMantRNE_36U_11U_i_data_3_sva[35:25])
      + conv_u2u_1_11(FpMantRNE_36U_11U_else_carry_2_sva);
  assign FpMantRNE_36U_11U_else_ac_int_cctor_3_sva = nl_FpMantRNE_36U_11U_else_ac_int_cctor_3_sva[10:0];
  assign FpAdd_8U_23U_b_right_shift_qr_3_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_7,
      FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_5);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_27_nl = ~ FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_5;
  assign FpAdd_8U_23U_a_right_shift_qr_3_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_7,
      (FpAdd_8U_23U_is_a_greater_oelse_not_27_nl));
  assign nl_FpMantRNE_36U_11U_else_ac_int_cctor_4_sva = (FpMantRNE_36U_11U_i_data_4_sva[35:25])
      + conv_u2u_1_11(FpMantRNE_36U_11U_else_carry_3_sva);
  assign FpMantRNE_36U_11U_else_ac_int_cctor_4_sva = nl_FpMantRNE_36U_11U_else_ac_int_cctor_4_sva[10:0];
  assign FpAdd_8U_23U_b_right_shift_qr_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_5,
      FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2);
  assign FpAdd_8U_23U_is_a_greater_oelse_not_29_nl = ~ FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2;
  assign FpAdd_8U_23U_a_right_shift_qr_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, z_out_5,
      (FpAdd_8U_23U_is_a_greater_oelse_not_29_nl));
  assign nl_FpMantRNE_36U_11U_else_ac_int_cctor_sva = (FpMantRNE_36U_11U_i_data_sva[35:25])
      + conv_u2u_1_11(FpMantRNE_36U_11U_else_carry_sva);
  assign FpMantRNE_36U_11U_else_ac_int_cctor_sva = nl_FpMantRNE_36U_11U_else_ac_int_cctor_sva[10:0];
  assign inp_lookup_1_IntSignedShiftRight_50U_5U_32U_obits_fixed_and_nl = (IntSignedShiftRight_50U_5U_32U_mbits_fixed_1_sva_1_80_14_1[0])
      & inp_lookup_1_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2;
  assign nl_IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_1_sva = conv_s2s_66_67(IntSignedShiftRight_50U_5U_32U_mbits_fixed_1_sva_1_80_14_1[66:1])
      + conv_u2s_1_67(inp_lookup_1_IntSignedShiftRight_50U_5U_32U_obits_fixed_and_nl);
  assign IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_1_sva = nl_IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_1_sva[66:0];
  assign IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_ovfl_1_sva = ~((IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_1_sva[66])
      | (~((IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_1_sva[65:31]!=35'b00000000000000000000000000000000000))));
  assign IntSignedShiftRight_50U_5U_32U_obits_fixed_and_unfl_1_sva = (IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_1_sva[66])
      & (~((IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_1_sva[65:31]==35'b11111111111111111111111111111111111)));
  assign mux_1980_nl = MUX_s_1_2_2((FpMul_6U_10U_2_p_mant_p1_1_sva[21]), (inp_lookup_1_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21]),
      nor_44_cse);
  assign FpMul_6U_10U_2_p_mant_20_1_1_lpi_1_dfm_3_mx0 = MUX_v_20_2_2((FpMul_6U_10U_2_p_mant_p1_1_sva_mx1_20_0[19:0]),
      (FpMul_6U_10U_2_p_mant_p1_1_sva_mx1_20_0[20:1]), mux_1980_nl);
  assign inp_lookup_2_IntSignedShiftRight_50U_5U_32U_obits_fixed_and_nl = (IntSignedShiftRight_50U_5U_32U_mbits_fixed_2_sva_1_80_14_1[0])
      & inp_lookup_2_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2;
  assign nl_IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_2_sva = conv_s2s_66_67(IntSignedShiftRight_50U_5U_32U_mbits_fixed_2_sva_1_80_14_1[66:1])
      + conv_u2s_1_67(inp_lookup_2_IntSignedShiftRight_50U_5U_32U_obits_fixed_and_nl);
  assign IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_2_sva = nl_IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_2_sva[66:0];
  assign IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_ovfl_2_sva = ~((IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_2_sva[66])
      | (~((IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_2_sva[65:31]!=35'b00000000000000000000000000000000000))));
  assign IntSignedShiftRight_50U_5U_32U_obits_fixed_and_unfl_2_sva = (IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_2_sva[66])
      & (~((IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_2_sva[65:31]==35'b11111111111111111111111111111111111)));
  assign nor_707_nl = ~((inp_lookup_2_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21]) | (~
      inp_lookup_2_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs)
      | FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_3);
  assign or_5639_nl = (~ (inp_lookup_2_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21])) | (~
      inp_lookup_2_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs)
      | FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_3;
  assign mux_1981_nl = MUX_s_1_2_2((or_5639_nl), (nor_707_nl), FpMul_6U_10U_2_p_mant_p1_2_sva[21]);
  assign FpMul_6U_10U_2_p_mant_20_1_2_lpi_1_dfm_3_mx0 = MUX_v_20_2_2((FpMul_6U_10U_2_p_mant_p1_2_sva_mx1_20_0[20:1]),
      (FpMul_6U_10U_2_p_mant_p1_2_sva_mx1_20_0[19:0]), mux_1981_nl);
  assign inp_lookup_3_IntSignedShiftRight_50U_5U_32U_obits_fixed_and_nl = (IntSignedShiftRight_50U_5U_32U_mbits_fixed_3_sva_1_80_14_1[0])
      & inp_lookup_3_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2;
  assign nl_IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_3_sva = conv_s2s_66_67(IntSignedShiftRight_50U_5U_32U_mbits_fixed_3_sva_1_80_14_1[66:1])
      + conv_u2s_1_67(inp_lookup_3_IntSignedShiftRight_50U_5U_32U_obits_fixed_and_nl);
  assign IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_3_sva = nl_IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_3_sva[66:0];
  assign IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_ovfl_3_sva = ~((IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_3_sva[66])
      | (~((IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_3_sva[65:31]!=35'b00000000000000000000000000000000000))));
  assign IntSignedShiftRight_50U_5U_32U_obits_fixed_and_unfl_3_sva = (IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_3_sva[66])
      & (~((IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_3_sva[65:31]==35'b11111111111111111111111111111111111)));
  assign nor_706_nl = ~(FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_3 | (~ inp_lookup_3_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs)
      | (inp_lookup_3_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21]));
  assign or_5638_nl = FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_3 | (~(inp_lookup_3_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs
      & (inp_lookup_3_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21])));
  assign mux_1982_nl = MUX_s_1_2_2((or_5638_nl), (nor_706_nl), FpMul_6U_10U_2_p_mant_p1_3_sva[21]);
  assign FpMul_6U_10U_2_p_mant_20_1_3_lpi_1_dfm_3_mx0 = MUX_v_20_2_2((FpMul_6U_10U_2_p_mant_p1_3_sva_mx1_20_0[20:1]),
      (FpMul_6U_10U_2_p_mant_p1_3_sva_mx1_20_0[19:0]), mux_1982_nl);
  assign inp_lookup_4_IntSignedShiftRight_50U_5U_32U_obits_fixed_and_nl = (IntSignedShiftRight_50U_5U_32U_mbits_fixed_sva_1_80_14_1[0])
      & inp_lookup_4_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2;
  assign nl_IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_sva = conv_s2s_66_67(IntSignedShiftRight_50U_5U_32U_mbits_fixed_sva_1_80_14_1[66:1])
      + conv_u2s_1_67(inp_lookup_4_IntSignedShiftRight_50U_5U_32U_obits_fixed_and_nl);
  assign IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_sva = nl_IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_sva[66:0];
  assign IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_ovfl_sva = ~((IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_sva[66])
      | (~((IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_sva[65:31]!=35'b00000000000000000000000000000000000))));
  assign IntSignedShiftRight_50U_5U_32U_obits_fixed_and_unfl_sva = (IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_sva[66])
      & (~((IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_sva[65:31]==35'b11111111111111111111111111111111111)));
  assign nor_705_nl = ~((inp_lookup_4_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21]) | (~
      inp_lookup_4_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs)
      | FpMul_6U_10U_2_lor_1_lpi_1_dfm_st_3);
  assign or_5637_nl = (~ (inp_lookup_4_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21])) | (~
      inp_lookup_4_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs)
      | FpMul_6U_10U_2_lor_1_lpi_1_dfm_st_3;
  assign mux_1983_nl = MUX_s_1_2_2((or_5637_nl), (nor_705_nl), FpMul_6U_10U_2_p_mant_p1_sva[21]);
  assign FpMul_6U_10U_2_p_mant_20_1_lpi_1_dfm_3_mx0 = MUX_v_20_2_2((FpMul_6U_10U_2_p_mant_p1_sva_mx1_20_0[20:1]),
      (FpMul_6U_10U_2_p_mant_p1_sva_mx1_20_0[19:0]), mux_1983_nl);
  assign or_5369_cse = (~ inp_lookup_1_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs)
      | FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_3;
  assign mux_1984_nl = MUX_s_1_2_2((inp_lookup_1_FpMul_6U_10U_1_p_mant_p1_mul_tmp[21]),
      (FpMul_6U_10U_1_p_mant_p1_1_sva[21]), or_5369_cse);
  assign FpMul_6U_10U_1_p_mant_20_1_1_lpi_1_dfm_3_mx0 = MUX_v_20_2_2((FpMul_6U_10U_1_p_mant_p1_1_sva_mx1_20_0[19:0]),
      (FpMul_6U_10U_1_p_mant_p1_1_sva_mx1_20_0[20:1]), mux_1984_nl);
  assign nl_inp_lookup_1_FpMul_6U_10U_2_else_2_else_if_if_acc_nl = reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_8_1_reg
      + 6'b1;
  assign inp_lookup_1_FpMul_6U_10U_2_else_2_else_if_if_acc_nl = nl_inp_lookup_1_FpMul_6U_10U_2_else_2_else_if_if_acc_nl[5:0];
  assign FpMul_6U_10U_2_p_expo_1_lpi_1_dfm_1_mx0 = MUX_v_6_2_2(reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_8_1_reg,
      (inp_lookup_1_FpMul_6U_10U_2_else_2_else_if_if_acc_nl), FpMul_6U_10U_2_else_2_else_and_itm_2);
  assign nl_FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_1_sva_1 = FpMul_6U_10U_2_p_expo_1_lpi_1_dfm_1_mx0
      + 6'b1;
  assign FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_1_sva_1 = nl_FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_1_sva_1[5:0];
  assign FpMantWidthDec_6U_21U_10U_0U_0U_2_if_1_unequal_tmp = ~((FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_1_sva_1==6'b111111));
  assign FpMul_6U_10U_2_and_ssc = IsNaN_6U_10U_7_land_1_lpi_1_dfm_6 & (~ IsNaN_6U_10U_6_land_1_lpi_1_dfm_5);
  assign FpMul_6U_10U_2_or_4_nl = ((~ FpMantWidthDec_6U_21U_10U_0U_0U_2_if_1_unequal_tmp)
      & FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_2) | nor_1274_cse;
  assign FpMantWidthDec_6U_21U_10U_0U_0U_2_and_1_nl = FpMantWidthDec_6U_21U_10U_0U_0U_2_if_1_unequal_tmp
      & FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_2 & (~ nor_1274_cse);
  assign FpMul_6U_10U_2_o_expo_1_lpi_1_dfm = MUX1HOT_v_6_3_2(FpMul_6U_10U_2_p_expo_1_lpi_1_dfm_1_mx0,
      6'b111110, FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_1_sva_1, {nor_1273_cse
      , (FpMul_6U_10U_2_or_4_nl) , (FpMantWidthDec_6U_21U_10U_0U_0U_2_and_1_nl)});
  assign FpMul_6U_10U_2_lor_9_lpi_1_dfm = (~((FpMul_6U_10U_2_o_expo_1_lpi_1_dfm!=6'b000000)))
      | FpMul_6U_10U_2_lor_6_lpi_1_dfm_6;
  assign nor_704_nl = ~((inp_lookup_2_FpMul_6U_10U_1_p_mant_p1_mul_tmp[21]) | (~
      inp_lookup_2_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs)
      | FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_3);
  assign or_5636_nl = (~ (inp_lookup_2_FpMul_6U_10U_1_p_mant_p1_mul_tmp[21])) | (~
      inp_lookup_2_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs)
      | FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_3;
  assign mux_1985_nl = MUX_s_1_2_2((or_5636_nl), (nor_704_nl), FpMul_6U_10U_1_p_mant_p1_2_sva[21]);
  assign FpMul_6U_10U_1_p_mant_20_1_2_lpi_1_dfm_3_mx0 = MUX_v_20_2_2((FpMul_6U_10U_1_p_mant_p1_2_sva_mx1_20_0[20:1]),
      (FpMul_6U_10U_1_p_mant_p1_2_sva_mx1_20_0[19:0]), mux_1985_nl);
  assign nl_inp_lookup_2_FpMul_6U_10U_2_else_2_else_if_if_acc_nl = FpMul_6U_10U_2_else_2_else_ac_int_cctor_2_sva_2
      + 6'b1;
  assign inp_lookup_2_FpMul_6U_10U_2_else_2_else_if_if_acc_nl = nl_inp_lookup_2_FpMul_6U_10U_2_else_2_else_if_if_acc_nl[5:0];
  assign FpMul_6U_10U_2_p_expo_2_lpi_1_dfm_1_mx0 = MUX_v_6_2_2(FpMul_6U_10U_2_else_2_else_ac_int_cctor_2_sva_2,
      (inp_lookup_2_FpMul_6U_10U_2_else_2_else_if_if_acc_nl), FpMul_6U_10U_2_else_2_else_and_1_itm_2);
  assign nl_FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_2_sva_1 = FpMul_6U_10U_2_p_expo_2_lpi_1_dfm_1_mx0
      + 6'b1;
  assign FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_2_sva_1 = nl_FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_2_sva_1[5:0];
  assign FpMantWidthDec_6U_21U_10U_0U_0U_2_if_1_unequal_tmp_1 = ~((FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_2_sva_1==6'b111111));
  assign FpMul_6U_10U_2_and_2_ssc = IsNaN_6U_10U_7_land_2_lpi_1_dfm_6 & (~ IsNaN_6U_10U_6_land_2_lpi_1_dfm_5);
  assign FpMul_6U_10U_2_or_5_nl = ((~ FpMantWidthDec_6U_21U_10U_0U_0U_2_if_1_unequal_tmp_1)
      & FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_2) | nor_1790_cse;
  assign FpMantWidthDec_6U_21U_10U_0U_0U_2_and_3_nl = FpMantWidthDec_6U_21U_10U_0U_0U_2_if_1_unequal_tmp_1
      & FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_2 & (~ nor_1790_cse);
  assign FpMul_6U_10U_2_o_expo_2_lpi_1_dfm = MUX1HOT_v_6_3_2(FpMul_6U_10U_2_p_expo_2_lpi_1_dfm_1_mx0,
      6'b111110, FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_2_sva_1, {nor_1264_cse
      , (FpMul_6U_10U_2_or_5_nl) , (FpMantWidthDec_6U_21U_10U_0U_0U_2_and_3_nl)});
  assign FpMul_6U_10U_2_lor_10_lpi_1_dfm = (~((FpMul_6U_10U_2_o_expo_2_lpi_1_dfm!=6'b000000)))
      | FpMul_6U_10U_2_lor_7_lpi_1_dfm_6;
  assign or_5372_cse = (~ inp_lookup_3_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs)
      | FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_3;
  assign mux_1986_nl = MUX_s_1_2_2((inp_lookup_3_FpMul_6U_10U_1_p_mant_p1_mul_tmp[21]),
      (FpMul_6U_10U_1_p_mant_p1_3_sva[21]), or_5372_cse);
  assign FpMul_6U_10U_1_p_mant_20_1_3_lpi_1_dfm_3_mx0 = MUX_v_20_2_2((FpMul_6U_10U_1_p_mant_p1_3_sva_mx1_20_0[19:0]),
      (FpMul_6U_10U_1_p_mant_p1_3_sva_mx1_20_0[20:1]), mux_1986_nl);
  assign nl_inp_lookup_3_FpMul_6U_10U_2_else_2_else_if_if_acc_nl = FpMul_6U_10U_2_else_2_else_ac_int_cctor_3_sva_2
      + 6'b1;
  assign inp_lookup_3_FpMul_6U_10U_2_else_2_else_if_if_acc_nl = nl_inp_lookup_3_FpMul_6U_10U_2_else_2_else_if_if_acc_nl[5:0];
  assign FpMul_6U_10U_2_p_expo_3_lpi_1_dfm_1_mx0 = MUX_v_6_2_2(FpMul_6U_10U_2_else_2_else_ac_int_cctor_3_sva_2,
      (inp_lookup_3_FpMul_6U_10U_2_else_2_else_if_if_acc_nl), FpMul_6U_10U_2_else_2_else_and_2_itm_2);
  assign nl_FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_3_sva_1 = FpMul_6U_10U_2_p_expo_3_lpi_1_dfm_1_mx0
      + 6'b1;
  assign FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_3_sva_1 = nl_FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_3_sva_1[5:0];
  assign FpMantWidthDec_6U_21U_10U_0U_0U_2_if_1_unequal_tmp_2 = ~((FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_3_sva_1==6'b111111));
  assign FpMul_6U_10U_2_and_4_ssc = IsNaN_6U_10U_7_land_3_lpi_1_dfm_6 & (~ IsNaN_6U_10U_6_land_3_lpi_1_dfm_5);
  assign FpMul_6U_10U_2_or_6_nl = ((~ FpMantWidthDec_6U_21U_10U_0U_0U_2_if_1_unequal_tmp_2)
      & FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_2) | nor_1789_cse;
  assign FpMantWidthDec_6U_21U_10U_0U_0U_2_and_5_nl = FpMantWidthDec_6U_21U_10U_0U_0U_2_if_1_unequal_tmp_2
      & FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_2 & (~ nor_1789_cse);
  assign FpMul_6U_10U_2_o_expo_3_lpi_1_dfm = MUX1HOT_v_6_3_2(FpMul_6U_10U_2_p_expo_3_lpi_1_dfm_1_mx0,
      6'b111110, FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_3_sva_1, {nor_1251_cse
      , (FpMul_6U_10U_2_or_6_nl) , (FpMantWidthDec_6U_21U_10U_0U_0U_2_and_5_nl)});
  assign FpMul_6U_10U_2_lor_11_lpi_1_dfm = (~((FpMul_6U_10U_2_o_expo_3_lpi_1_dfm!=6'b000000)))
      | FpMul_6U_10U_2_lor_8_lpi_1_dfm_6;
  assign mux_1987_nl = MUX_s_1_2_2((inp_lookup_4_FpMul_6U_10U_1_p_mant_p1_mul_tmp[21]),
      (FpMul_6U_10U_1_p_mant_p1_sva[21]), or_3779_cse);
  assign FpMul_6U_10U_1_p_mant_20_1_lpi_1_dfm_3_mx0 = MUX_v_20_2_2((FpMul_6U_10U_1_p_mant_p1_sva_mx1_20_0[19:0]),
      (FpMul_6U_10U_1_p_mant_p1_sva_mx1_20_0[20:1]), mux_1987_nl);
  assign nl_inp_lookup_4_FpMul_6U_10U_2_else_2_else_if_if_acc_nl = reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_8_1_reg
      + 6'b1;
  assign inp_lookup_4_FpMul_6U_10U_2_else_2_else_if_if_acc_nl = nl_inp_lookup_4_FpMul_6U_10U_2_else_2_else_if_if_acc_nl[5:0];
  assign FpMul_6U_10U_2_p_expo_lpi_1_dfm_1_mx0 = MUX_v_6_2_2(reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_8_1_reg,
      (inp_lookup_4_FpMul_6U_10U_2_else_2_else_if_if_acc_nl), FpMul_6U_10U_2_else_2_else_and_3_itm_2);
  assign nl_FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_sva_1 = FpMul_6U_10U_2_p_expo_lpi_1_dfm_1_mx0
      + 6'b1;
  assign FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_sva_1 = nl_FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_sva_1[5:0];
  assign FpMantWidthDec_6U_21U_10U_0U_0U_2_if_1_unequal_tmp_3 = ~((FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_sva_1==6'b111111));
  assign FpMul_6U_10U_2_and_6_ssc = IsNaN_6U_10U_7_land_lpi_1_dfm_6 & (~ IsNaN_6U_10U_6_land_lpi_1_dfm_5);
  assign FpMul_6U_10U_2_or_7_nl = ((~ FpMantWidthDec_6U_21U_10U_0U_0U_2_if_1_unequal_tmp_3)
      & FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_sva_2) | nor_1238_cse;
  assign FpMantWidthDec_6U_21U_10U_0U_0U_2_and_7_nl = FpMantWidthDec_6U_21U_10U_0U_0U_2_if_1_unequal_tmp_3
      & FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_sva_2 & (~ nor_1238_cse);
  assign FpMul_6U_10U_2_o_expo_lpi_1_dfm = MUX1HOT_v_6_3_2(FpMul_6U_10U_2_p_expo_lpi_1_dfm_1_mx0,
      6'b111110, FpMantWidthDec_6U_21U_10U_0U_0U_2_o_expo_sva_1, {nor_1237_cse ,
      (FpMul_6U_10U_2_or_7_nl) , (FpMantWidthDec_6U_21U_10U_0U_0U_2_and_7_nl)});
  assign FpMul_6U_10U_2_lor_2_lpi_1_dfm = (~((FpMul_6U_10U_2_o_expo_lpi_1_dfm!=6'b000000)))
      | FpMul_6U_10U_2_lor_1_lpi_1_dfm_6;
  assign FpAdd_8U_23U_1_addend_larger_qr_1_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_1_addend_larger_asn_19_mx0w1,
      FpAdd_8U_23U_1_a_int_mant_p1_1_sva, FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5);
  assign FpAdd_8U_23U_1_addend_smaller_qr_1_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_1_a_int_mant_p1_1_sva,
      FpAdd_8U_23U_1_addend_larger_asn_19_mx0w1, FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5);
  assign nl_inp_lookup_1_FpAdd_8U_23U_1_b_right_shift_qif_acc_nl = (chn_inp_in_crt_sva_4_127_0_1[30:23])
      + ({(~ reg_FpAdd_8U_23U_o_expo_1_lpi_1_dfm_11_reg) , (~ reg_FpAdd_8U_23U_o_expo_1_lpi_1_dfm_11_1_reg)})
      + 8'b1;
  assign inp_lookup_1_FpAdd_8U_23U_1_b_right_shift_qif_acc_nl = nl_inp_lookup_1_FpAdd_8U_23U_1_b_right_shift_qif_acc_nl[7:0];
  assign FpAdd_8U_23U_1_b_right_shift_qr_1_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, (inp_lookup_1_FpAdd_8U_23U_1_b_right_shift_qif_acc_nl),
      FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5);
  assign nl_inp_lookup_1_FpAdd_8U_23U_1_a_right_shift_qelse_acc_nl = ({reg_FpAdd_8U_23U_o_expo_1_lpi_1_dfm_11_reg
      , reg_FpAdd_8U_23U_o_expo_1_lpi_1_dfm_11_1_reg}) - (chn_inp_in_crt_sva_4_127_0_1[30:23]);
  assign inp_lookup_1_FpAdd_8U_23U_1_a_right_shift_qelse_acc_nl = nl_inp_lookup_1_FpAdd_8U_23U_1_a_right_shift_qelse_acc_nl[7:0];
  assign FpAdd_8U_23U_1_is_a_greater_oelse_not_23_nl = ~ FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5;
  assign FpAdd_8U_23U_1_a_right_shift_qr_1_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, (inp_lookup_1_FpAdd_8U_23U_1_a_right_shift_qelse_acc_nl),
      (FpAdd_8U_23U_1_is_a_greater_oelse_not_23_nl));
  assign FpAdd_8U_23U_1_addend_larger_qr_2_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_1_addend_larger_asn_13_mx0w1,
      FpAdd_8U_23U_1_a_int_mant_p1_2_sva, FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5);
  assign FpAdd_8U_23U_1_addend_smaller_qr_2_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_1_a_int_mant_p1_2_sva,
      FpAdd_8U_23U_1_addend_larger_asn_13_mx0w1, FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5);
  assign nl_inp_lookup_2_FpAdd_8U_23U_1_b_right_shift_qif_acc_nl = (chn_inp_in_crt_sva_4_127_0_1[62:55])
      + ({(~ reg_FpAdd_8U_23U_o_expo_2_lpi_1_dfm_11_reg) , (~ reg_FpAdd_8U_23U_o_expo_2_lpi_1_dfm_11_1_reg)})
      + 8'b1;
  assign inp_lookup_2_FpAdd_8U_23U_1_b_right_shift_qif_acc_nl = nl_inp_lookup_2_FpAdd_8U_23U_1_b_right_shift_qif_acc_nl[7:0];
  assign FpAdd_8U_23U_1_b_right_shift_qr_2_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, (inp_lookup_2_FpAdd_8U_23U_1_b_right_shift_qif_acc_nl),
      FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5);
  assign nl_inp_lookup_2_FpAdd_8U_23U_1_a_right_shift_qelse_acc_nl = ({reg_FpAdd_8U_23U_o_expo_2_lpi_1_dfm_11_reg
      , reg_FpAdd_8U_23U_o_expo_2_lpi_1_dfm_11_1_reg}) - (chn_inp_in_crt_sva_4_127_0_1[62:55]);
  assign inp_lookup_2_FpAdd_8U_23U_1_a_right_shift_qelse_acc_nl = nl_inp_lookup_2_FpAdd_8U_23U_1_a_right_shift_qelse_acc_nl[7:0];
  assign FpAdd_8U_23U_1_is_a_greater_oelse_not_25_nl = ~ FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5;
  assign FpAdd_8U_23U_1_a_right_shift_qr_2_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, (inp_lookup_2_FpAdd_8U_23U_1_a_right_shift_qelse_acc_nl),
      (FpAdd_8U_23U_1_is_a_greater_oelse_not_25_nl));
  assign FpAdd_8U_23U_1_addend_larger_qr_3_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_1_addend_larger_asn_7_mx0w1,
      FpAdd_8U_23U_1_a_int_mant_p1_3_sva, FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5);
  assign FpAdd_8U_23U_1_addend_smaller_qr_3_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_1_a_int_mant_p1_3_sva,
      FpAdd_8U_23U_1_addend_larger_asn_7_mx0w1, FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5);
  assign nl_inp_lookup_3_FpAdd_8U_23U_1_b_right_shift_qif_acc_nl = (chn_inp_in_crt_sva_4_127_0_1[94:87])
      + ({(~ reg_FpAdd_8U_23U_o_expo_3_lpi_1_dfm_11_reg) , (~ reg_FpAdd_8U_23U_o_expo_3_lpi_1_dfm_11_1_reg)})
      + 8'b1;
  assign inp_lookup_3_FpAdd_8U_23U_1_b_right_shift_qif_acc_nl = nl_inp_lookup_3_FpAdd_8U_23U_1_b_right_shift_qif_acc_nl[7:0];
  assign FpAdd_8U_23U_1_b_right_shift_qr_3_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, (inp_lookup_3_FpAdd_8U_23U_1_b_right_shift_qif_acc_nl),
      FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5);
  assign nl_inp_lookup_3_FpAdd_8U_23U_1_a_right_shift_qelse_acc_nl = ({reg_FpAdd_8U_23U_o_expo_3_lpi_1_dfm_11_reg
      , reg_FpAdd_8U_23U_o_expo_3_lpi_1_dfm_11_1_reg}) - (chn_inp_in_crt_sva_4_127_0_1[94:87]);
  assign inp_lookup_3_FpAdd_8U_23U_1_a_right_shift_qelse_acc_nl = nl_inp_lookup_3_FpAdd_8U_23U_1_a_right_shift_qelse_acc_nl[7:0];
  assign FpAdd_8U_23U_1_is_a_greater_oelse_not_27_nl = ~ FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5;
  assign FpAdd_8U_23U_1_a_right_shift_qr_3_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, (inp_lookup_3_FpAdd_8U_23U_1_a_right_shift_qelse_acc_nl),
      (FpAdd_8U_23U_1_is_a_greater_oelse_not_27_nl));
  assign FpAdd_8U_23U_1_addend_larger_qr_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_1_addend_larger_asn_1_mx0w1,
      FpAdd_8U_23U_1_a_int_mant_p1_sva, FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5);
  assign FpAdd_8U_23U_1_addend_smaller_qr_lpi_1_dfm_mx0 = MUX_v_49_2_2(FpAdd_8U_23U_1_a_int_mant_p1_sva,
      FpAdd_8U_23U_1_addend_larger_asn_1_mx0w1, FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5);
  assign nl_inp_lookup_4_FpAdd_8U_23U_1_b_right_shift_qif_acc_nl = (chn_inp_in_crt_sva_4_127_0_1[126:119])
      + ({(~ reg_FpAdd_8U_23U_o_expo_lpi_1_dfm_11_reg) , (~ reg_FpAdd_8U_23U_o_expo_lpi_1_dfm_11_1_reg)})
      + 8'b1;
  assign inp_lookup_4_FpAdd_8U_23U_1_b_right_shift_qif_acc_nl = nl_inp_lookup_4_FpAdd_8U_23U_1_b_right_shift_qif_acc_nl[7:0];
  assign FpAdd_8U_23U_1_b_right_shift_qr_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, (inp_lookup_4_FpAdd_8U_23U_1_b_right_shift_qif_acc_nl),
      FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5);
  assign nl_inp_lookup_4_FpAdd_8U_23U_1_a_right_shift_qelse_acc_nl = ({reg_FpAdd_8U_23U_o_expo_lpi_1_dfm_11_reg
      , reg_FpAdd_8U_23U_o_expo_lpi_1_dfm_11_1_reg}) - (chn_inp_in_crt_sva_4_127_0_1[126:119]);
  assign inp_lookup_4_FpAdd_8U_23U_1_a_right_shift_qelse_acc_nl = nl_inp_lookup_4_FpAdd_8U_23U_1_a_right_shift_qelse_acc_nl[7:0];
  assign FpAdd_8U_23U_1_is_a_greater_oelse_not_29_nl = ~ FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5;
  assign FpAdd_8U_23U_1_a_right_shift_qr_lpi_1_dfm = MUX_v_8_2_2(8'b00000000, (inp_lookup_4_FpAdd_8U_23U_1_a_right_shift_qelse_acc_nl),
      (FpAdd_8U_23U_1_is_a_greater_oelse_not_29_nl));
  assign nl_FpAdd_6U_10U_1_o_expo_1_sva_4 = ({FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_5
      , FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_4 , FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_3_0})
      + 6'b1;
  assign FpAdd_6U_10U_1_o_expo_1_sva_4 = nl_FpAdd_6U_10U_1_o_expo_1_sva_4[5:0];
  assign FpAdd_6U_10U_1_if_4_FpAdd_6U_10U_1_if_4_or_nl = FpAdd_6U_10U_1_and_4_ssc
      | (~ (z_out_8[5]));
  assign FpAdd_6U_10U_1_is_inf_1_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_1_and_4_ssc,
      (FpAdd_6U_10U_1_if_4_FpAdd_6U_10U_1_if_4_or_nl), inp_lookup_1_FpMantRNE_23U_11U_1_else_and_tmp);
  assign FpAdd_6U_10U_1_and_ssc = (~(FpAdd_6U_10U_1_and_tmp | FpAdd_6U_10U_1_is_inf_1_lpi_1_dfm_2_mx0))
      & nor_1727_cse;
  assign FpAdd_6U_10U_1_and_6_ssc = FpAdd_6U_10U_1_and_tmp & (~ FpAdd_6U_10U_1_is_inf_1_lpi_1_dfm_2_mx0)
      & nor_1727_cse;
  assign FpAdd_6U_10U_1_and_28_ssc = FpAdd_6U_10U_1_is_inf_1_lpi_1_dfm_2_mx0 & nor_1727_cse;
  assign FpAdd_6U_10U_1_and_tmp = (z_out_8[5]) & inp_lookup_1_FpMantRNE_23U_11U_1_else_and_tmp;
  assign nl_FpAdd_6U_10U_1_o_expo_2_sva_4 = ({FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_5
      , FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_4 , FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_3_0})
      + 6'b1;
  assign FpAdd_6U_10U_1_o_expo_2_sva_4 = nl_FpAdd_6U_10U_1_o_expo_2_sva_4[5:0];
  assign FpAdd_6U_10U_1_if_4_FpAdd_6U_10U_1_if_4_or_1_nl = FpAdd_6U_10U_1_and_10_ssc
      | (~ (z_out_9[5]));
  assign FpAdd_6U_10U_1_is_inf_2_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_1_and_10_ssc,
      (FpAdd_6U_10U_1_if_4_FpAdd_6U_10U_1_if_4_or_1_nl), inp_lookup_2_FpMantRNE_23U_11U_1_else_and_tmp);
  assign FpAdd_6U_10U_1_and_29_ssc = (~(FpAdd_6U_10U_1_and_1_tmp | FpAdd_6U_10U_1_is_inf_2_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_7_m1c;
  assign FpAdd_6U_10U_1_and_13_ssc = FpAdd_6U_10U_1_and_1_tmp & (~ FpAdd_6U_10U_1_is_inf_2_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_7_m1c;
  assign FpAdd_6U_10U_1_and_30_ssc = FpAdd_6U_10U_1_is_inf_2_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_7_m1c;
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_7_m1c = ~(IsNaN_6U_10U_9_land_2_lpi_1_dfm_8
      | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_19);
  assign FpAdd_6U_10U_1_and_1_tmp = (z_out_9[5]) & inp_lookup_2_FpMantRNE_23U_11U_1_else_and_tmp;
  assign nl_FpAdd_6U_10U_1_o_expo_3_sva_4 = ({FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_5
      , FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_4 , FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_3_0})
      + 6'b1;
  assign FpAdd_6U_10U_1_o_expo_3_sva_4 = nl_FpAdd_6U_10U_1_o_expo_3_sva_4[5:0];
  assign FpAdd_6U_10U_1_if_4_FpAdd_6U_10U_1_if_4_or_2_nl = FpAdd_6U_10U_1_and_16_ssc
      | (~ (z_out_10[5]));
  assign FpAdd_6U_10U_1_is_inf_3_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_1_and_16_ssc,
      (FpAdd_6U_10U_1_if_4_FpAdd_6U_10U_1_if_4_or_2_nl), inp_lookup_3_FpMantRNE_23U_11U_1_else_and_tmp);
  assign FpAdd_6U_10U_1_and_31_ssc = (~(FpAdd_6U_10U_1_and_2_tmp | FpAdd_6U_10U_1_is_inf_3_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_9_m1c;
  assign FpAdd_6U_10U_1_and_19_ssc = FpAdd_6U_10U_1_and_2_tmp & (~ FpAdd_6U_10U_1_is_inf_3_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_9_m1c;
  assign FpAdd_6U_10U_1_and_32_ssc = FpAdd_6U_10U_1_is_inf_3_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_9_m1c;
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_9_m1c = ~(IsNaN_6U_10U_9_land_3_lpi_1_dfm_8
      | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_19);
  assign FpAdd_6U_10U_1_and_2_tmp = (z_out_10[5]) & inp_lookup_3_FpMantRNE_23U_11U_1_else_and_tmp;
  assign nl_FpAdd_6U_10U_1_o_expo_sva_4 = ({FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_5 ,
      FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_4 , FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_3_0})
      + 6'b1;
  assign FpAdd_6U_10U_1_o_expo_sva_4 = nl_FpAdd_6U_10U_1_o_expo_sva_4[5:0];
  assign FpAdd_6U_10U_1_if_4_FpAdd_6U_10U_1_if_4_or_3_nl = FpAdd_6U_10U_1_and_22_ssc
      | (~ (z_out_11[5]));
  assign FpAdd_6U_10U_1_is_inf_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_1_and_22_ssc,
      (FpAdd_6U_10U_1_if_4_FpAdd_6U_10U_1_if_4_or_3_nl), inp_lookup_4_FpMantRNE_23U_11U_1_else_and_tmp);
  assign FpAdd_6U_10U_1_and_33_ssc = (~(FpAdd_6U_10U_1_and_3_tmp | FpAdd_6U_10U_1_is_inf_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_11_m1c;
  assign FpAdd_6U_10U_1_and_25_ssc = FpAdd_6U_10U_1_and_3_tmp & (~ FpAdd_6U_10U_1_is_inf_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_11_m1c;
  assign FpAdd_6U_10U_1_and_34_ssc = FpAdd_6U_10U_1_is_inf_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_11_m1c;
  assign FpAdd_6U_10U_1_FpAdd_6U_10U_1_nor_11_m1c = ~(IsNaN_6U_10U_9_land_lpi_1_dfm_8
      | IsNaN_6U_10U_2_land_lpi_1_dfm_st_18);
  assign FpAdd_6U_10U_1_and_3_tmp = (z_out_11[5]) & inp_lookup_4_FpMantRNE_23U_11U_1_else_and_tmp;
  assign nl_inp_lookup_1_FpMul_6U_10U_else_2_else_if_if_acc_nl = FpMul_6U_10U_else_2_else_ac_int_cctor_1_sva_2
      + 6'b1;
  assign inp_lookup_1_FpMul_6U_10U_else_2_else_if_if_acc_nl = nl_inp_lookup_1_FpMul_6U_10U_else_2_else_if_if_acc_nl[5:0];
  assign nand_643_nl = ~(inp_lookup_1_FpMul_6U_10U_else_2_else_if_if_acc_1_itm_5_1
      & (FpMul_6U_10U_p_mant_p1_1_sva_2[21]));
  assign FpMul_6U_10U_p_expo_1_lpi_1_dfm_1_mx0 = MUX_v_6_2_2((inp_lookup_1_FpMul_6U_10U_else_2_else_if_if_acc_nl),
      FpMul_6U_10U_else_2_else_ac_int_cctor_1_sva_2, nand_643_nl);
  assign FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp = ~((FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_1_sva_1==6'b111111));
  assign nl_FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_1_sva_1 = FpMul_6U_10U_p_expo_1_lpi_1_dfm_1_mx0
      + 6'b1;
  assign FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_1_sva_1 = nl_FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_1_sva_1[5:0];
  assign FpMul_6U_10U_is_inf_1_lpi_1_dfm_2 = ~(((inp_lookup_1_FpMul_6U_10U_else_2_else_if_if_acc_1_itm_5_1
      | (~ (FpMul_6U_10U_p_mant_p1_1_sva_2[21]))) & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_14_0_1)
      | FpMul_6U_10U_lor_6_lpi_1_dfm_4);
  assign FpMul_6U_10U_lor_9_lpi_1_dfm = (~((FpMul_6U_10U_o_expo_1_lpi_1_dfm!=6'b000000)))
      | FpMul_6U_10U_lor_6_lpi_1_dfm_4;
  assign FpMul_6U_10U_FpMul_6U_10U_nor_ssc = ~(IsNaN_6U_10U_1_land_1_lpi_1_dfm_6
      | IsNaN_6U_10U_land_1_lpi_1_dfm_6);
  assign FpMul_6U_10U_and_ssc = IsNaN_6U_10U_1_land_1_lpi_1_dfm_6 & (~ IsNaN_6U_10U_land_1_lpi_1_dfm_6);
  assign FpMul_6U_10U_FpMul_6U_10U_nor_8_nl = ~(inp_lookup_1_FpMantRNE_22U_11U_else_and_svs
      | FpMul_6U_10U_is_inf_1_lpi_1_dfm_2);
  assign FpMul_6U_10U_or_4_nl = ((~ FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp)
      & inp_lookup_1_FpMantRNE_22U_11U_else_and_svs) | FpMul_6U_10U_is_inf_1_lpi_1_dfm_2;
  assign FpMantWidthDec_6U_21U_10U_0U_0U_and_1_nl = FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp
      & inp_lookup_1_FpMantRNE_22U_11U_else_and_svs & (~ FpMul_6U_10U_is_inf_1_lpi_1_dfm_2);
  assign FpMul_6U_10U_o_expo_1_lpi_1_dfm = MUX1HOT_v_6_3_2(FpMul_6U_10U_p_expo_1_lpi_1_dfm_1_mx0,
      6'b111110, FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_1_sva_1, {(FpMul_6U_10U_FpMul_6U_10U_nor_8_nl)
      , (FpMul_6U_10U_or_4_nl) , (FpMantWidthDec_6U_21U_10U_0U_0U_and_1_nl)});
  assign nl_inp_lookup_2_FpMul_6U_10U_else_2_else_if_if_acc_nl = FpMul_6U_10U_else_2_else_ac_int_cctor_2_sva_2
      + 6'b1;
  assign inp_lookup_2_FpMul_6U_10U_else_2_else_if_if_acc_nl = nl_inp_lookup_2_FpMul_6U_10U_else_2_else_if_if_acc_nl[5:0];
  assign nand_642_nl = ~(inp_lookup_2_FpMul_6U_10U_else_2_else_if_if_acc_1_itm_5_1
      & (FpMul_6U_10U_p_mant_p1_2_sva_2[21]));
  assign FpMul_6U_10U_p_expo_2_lpi_1_dfm_1_mx0 = MUX_v_6_2_2((inp_lookup_2_FpMul_6U_10U_else_2_else_if_if_acc_nl),
      FpMul_6U_10U_else_2_else_ac_int_cctor_2_sva_2, nand_642_nl);
  assign FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp_1 = ~((FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_2_sva_1==6'b111111));
  assign nl_FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_2_sva_1 = FpMul_6U_10U_p_expo_2_lpi_1_dfm_1_mx0
      + 6'b1;
  assign FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_2_sva_1 = nl_FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_2_sva_1[5:0];
  assign FpMul_6U_10U_is_inf_2_lpi_1_dfm_2 = ~(((inp_lookup_2_FpMul_6U_10U_else_2_else_if_if_acc_1_itm_5_1
      | (~ (FpMul_6U_10U_p_mant_p1_2_sva_2[21]))) & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_14_0_1)
      | FpMul_6U_10U_lor_7_lpi_1_dfm_4);
  assign FpMul_6U_10U_lor_10_lpi_1_dfm = (~((FpMul_6U_10U_o_expo_2_lpi_1_dfm!=6'b000000)))
      | FpMul_6U_10U_lor_7_lpi_1_dfm_4;
  assign FpMul_6U_10U_FpMul_6U_10U_nor_1_ssc = ~(IsNaN_6U_10U_1_land_2_lpi_1_dfm_6
      | IsNaN_6U_10U_land_2_lpi_1_dfm_6);
  assign FpMul_6U_10U_and_2_ssc = IsNaN_6U_10U_1_land_2_lpi_1_dfm_6 & (~ IsNaN_6U_10U_land_2_lpi_1_dfm_6);
  assign FpMul_6U_10U_FpMul_6U_10U_nor_9_nl = ~(inp_lookup_2_FpMantRNE_22U_11U_else_and_svs
      | FpMul_6U_10U_is_inf_2_lpi_1_dfm_2);
  assign FpMul_6U_10U_or_5_nl = ((~ FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp_1)
      & inp_lookup_2_FpMantRNE_22U_11U_else_and_svs) | FpMul_6U_10U_is_inf_2_lpi_1_dfm_2;
  assign FpMantWidthDec_6U_21U_10U_0U_0U_and_3_nl = FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp_1
      & inp_lookup_2_FpMantRNE_22U_11U_else_and_svs & (~ FpMul_6U_10U_is_inf_2_lpi_1_dfm_2);
  assign FpMul_6U_10U_o_expo_2_lpi_1_dfm = MUX1HOT_v_6_3_2(FpMul_6U_10U_p_expo_2_lpi_1_dfm_1_mx0,
      6'b111110, FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_2_sva_1, {(FpMul_6U_10U_FpMul_6U_10U_nor_9_nl)
      , (FpMul_6U_10U_or_5_nl) , (FpMantWidthDec_6U_21U_10U_0U_0U_and_3_nl)});
  assign nl_inp_lookup_3_FpMul_6U_10U_else_2_else_if_if_acc_nl = FpMul_6U_10U_else_2_else_ac_int_cctor_3_sva_2
      + 6'b1;
  assign inp_lookup_3_FpMul_6U_10U_else_2_else_if_if_acc_nl = nl_inp_lookup_3_FpMul_6U_10U_else_2_else_if_if_acc_nl[5:0];
  assign nand_641_nl = ~(inp_lookup_3_FpMul_6U_10U_else_2_else_if_if_acc_1_itm_5_1
      & (FpMul_6U_10U_p_mant_p1_3_sva_2[21]));
  assign FpMul_6U_10U_p_expo_3_lpi_1_dfm_1_mx0 = MUX_v_6_2_2((inp_lookup_3_FpMul_6U_10U_else_2_else_if_if_acc_nl),
      FpMul_6U_10U_else_2_else_ac_int_cctor_3_sva_2, nand_641_nl);
  assign FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp_2 = ~((FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_3_sva_1==6'b111111));
  assign nl_FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_3_sva_1 = FpMul_6U_10U_p_expo_3_lpi_1_dfm_1_mx0
      + 6'b1;
  assign FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_3_sva_1 = nl_FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_3_sva_1[5:0];
  assign FpMul_6U_10U_is_inf_3_lpi_1_dfm_2 = ~(((inp_lookup_3_FpMul_6U_10U_else_2_else_if_if_acc_1_itm_5_1
      | (~ (FpMul_6U_10U_p_mant_p1_3_sva_2[21]))) & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_14_0_1)
      | FpMul_6U_10U_lor_8_lpi_1_dfm_4);
  assign FpMul_6U_10U_lor_11_lpi_1_dfm = (~((FpMul_6U_10U_o_expo_3_lpi_1_dfm!=6'b000000)))
      | FpMul_6U_10U_lor_8_lpi_1_dfm_4;
  assign FpMul_6U_10U_FpMul_6U_10U_nor_2_ssc = ~(IsNaN_6U_10U_1_land_3_lpi_1_dfm_6
      | IsNaN_6U_10U_land_3_lpi_1_dfm_6);
  assign FpMul_6U_10U_and_4_ssc = IsNaN_6U_10U_1_land_3_lpi_1_dfm_6 & (~ IsNaN_6U_10U_land_3_lpi_1_dfm_6);
  assign FpMul_6U_10U_FpMul_6U_10U_nor_10_nl = ~(inp_lookup_3_FpMantRNE_22U_11U_else_and_svs
      | FpMul_6U_10U_is_inf_3_lpi_1_dfm_2);
  assign FpMul_6U_10U_or_6_nl = ((~ FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp_2)
      & inp_lookup_3_FpMantRNE_22U_11U_else_and_svs) | FpMul_6U_10U_is_inf_3_lpi_1_dfm_2;
  assign FpMantWidthDec_6U_21U_10U_0U_0U_and_5_nl = FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp_2
      & inp_lookup_3_FpMantRNE_22U_11U_else_and_svs & (~ FpMul_6U_10U_is_inf_3_lpi_1_dfm_2);
  assign FpMul_6U_10U_o_expo_3_lpi_1_dfm = MUX1HOT_v_6_3_2(FpMul_6U_10U_p_expo_3_lpi_1_dfm_1_mx0,
      6'b111110, FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_3_sva_1, {(FpMul_6U_10U_FpMul_6U_10U_nor_10_nl)
      , (FpMul_6U_10U_or_6_nl) , (FpMantWidthDec_6U_21U_10U_0U_0U_and_5_nl)});
  assign nl_inp_lookup_4_FpMul_6U_10U_else_2_else_if_if_acc_nl = FpMul_6U_10U_else_2_else_ac_int_cctor_sva_2
      + 6'b1;
  assign inp_lookup_4_FpMul_6U_10U_else_2_else_if_if_acc_nl = nl_inp_lookup_4_FpMul_6U_10U_else_2_else_if_if_acc_nl[5:0];
  assign nand_640_nl = ~(inp_lookup_4_FpMul_6U_10U_else_2_else_if_if_acc_1_itm_5_1
      & (FpMul_6U_10U_p_mant_p1_sva_2[21]));
  assign FpMul_6U_10U_p_expo_lpi_1_dfm_1_mx0 = MUX_v_6_2_2((inp_lookup_4_FpMul_6U_10U_else_2_else_if_if_acc_nl),
      FpMul_6U_10U_else_2_else_ac_int_cctor_sva_2, nand_640_nl);
  assign FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp_3 = ~((FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_sva_1==6'b111111));
  assign nl_FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_sva_1 = FpMul_6U_10U_p_expo_lpi_1_dfm_1_mx0
      + 6'b1;
  assign FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_sva_1 = nl_FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_sva_1[5:0];
  assign FpMul_6U_10U_is_inf_lpi_1_dfm_2 = ~(((inp_lookup_4_FpMul_6U_10U_else_2_else_if_if_acc_1_itm_5_1
      | (~ (FpMul_6U_10U_p_mant_p1_sva_2[21]))) & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_14_0_1)
      | FpMul_6U_10U_lor_1_lpi_1_dfm_4);
  assign FpMul_6U_10U_lor_2_lpi_1_dfm = (~((FpMul_6U_10U_o_expo_lpi_1_dfm!=6'b000000)))
      | FpMul_6U_10U_lor_1_lpi_1_dfm_4;
  assign FpMul_6U_10U_FpMul_6U_10U_nor_3_ssc = ~(IsNaN_6U_10U_1_land_lpi_1_dfm_6
      | IsNaN_6U_10U_land_lpi_1_dfm_6);
  assign FpMul_6U_10U_and_6_ssc = IsNaN_6U_10U_1_land_lpi_1_dfm_6 & (~ IsNaN_6U_10U_land_lpi_1_dfm_6);
  assign FpMul_6U_10U_FpMul_6U_10U_nor_11_nl = ~(inp_lookup_4_FpMantRNE_22U_11U_else_and_svs
      | FpMul_6U_10U_is_inf_lpi_1_dfm_2);
  assign FpMul_6U_10U_or_7_nl = ((~ FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp_3)
      & inp_lookup_4_FpMantRNE_22U_11U_else_and_svs) | FpMul_6U_10U_is_inf_lpi_1_dfm_2;
  assign FpMantWidthDec_6U_21U_10U_0U_0U_and_7_nl = FpMantWidthDec_6U_21U_10U_0U_0U_if_1_unequal_tmp_3
      & inp_lookup_4_FpMantRNE_22U_11U_else_and_svs & (~ FpMul_6U_10U_is_inf_lpi_1_dfm_2);
  assign FpMul_6U_10U_o_expo_lpi_1_dfm = MUX1HOT_v_6_3_2(FpMul_6U_10U_p_expo_lpi_1_dfm_1_mx0,
      6'b111110, FpMantWidthDec_6U_21U_10U_0U_0U_o_expo_sva_1, {(FpMul_6U_10U_FpMul_6U_10U_nor_11_nl)
      , (FpMul_6U_10U_or_7_nl) , (FpMantWidthDec_6U_21U_10U_0U_0U_and_7_nl)});
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_1_sva = ({1'b1 , (~
      libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_20)}) + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_1_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_1_sva[4:0];
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_1_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((chn_inp_in_rsci_d_mxwt[277:268]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_or_mx0w1,
      or_dcpl_1005);
  assign IsZero_5U_10U_2_land_1_lpi_1_dfm = ~((chn_inp_in_rsci_d_mxwt[277:268]!=10'b0000000000)
      | (~ IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_1_sva));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_cse
      = ~(IsDenorm_5U_10U_2_land_1_lpi_1_dfm | IsInf_5U_10U_1_land_1_lpi_1_dfm);
  assign IsInf_5U_10U_1_land_1_lpi_1_dfm = ~((chn_inp_in_rsci_d_mxwt[277:268]!=10'b0000000000)
      | (~ IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_1_sva));
  assign IsNaN_5U_10U_1_land_1_lpi_1_dfm = IsDenorm_5U_10U_2_or_tmp & IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_1_sva;
  assign IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_1_sva = (chn_inp_in_rsci_d_mxwt[282:278]==5'b11111);
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_2_sva = ({1'b1 , (~
      libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_21)}) + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_2_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_2_sva[4:0];
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_2_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((chn_inp_in_rsci_d_mxwt[293:284]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_or_4_mx0w1,
      or_dcpl_1010);
  assign IsZero_5U_10U_2_land_2_lpi_1_dfm = ~((chn_inp_in_rsci_d_mxwt[293:284]!=10'b0000000000)
      | (~ IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_2_sva));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_1_cse
      = ~(IsDenorm_5U_10U_2_land_2_lpi_1_dfm | IsInf_5U_10U_1_land_2_lpi_1_dfm);
  assign IsInf_5U_10U_1_land_2_lpi_1_dfm = ~((chn_inp_in_rsci_d_mxwt[293:284]!=10'b0000000000)
      | (~ IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_2_sva));
  assign IsNaN_5U_10U_1_land_2_lpi_1_dfm = IsDenorm_5U_10U_2_or_1_tmp & IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_2_sva;
  assign IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_2_sva = (chn_inp_in_rsci_d_mxwt[298:294]==5'b11111);
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_3_sva = ({1'b1 , (~
      libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_22)}) + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_3_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_3_sva[4:0];
  assign IsZero_5U_10U_2_land_3_lpi_1_dfm = ~((chn_inp_in_rsci_d_mxwt[309:300]!=10'b0000000000)
      | (~ IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_3_sva));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_2_cse
      = ~(IsDenorm_5U_10U_2_land_3_lpi_1_dfm | IsInf_5U_10U_1_land_3_lpi_1_dfm);
  assign IsInf_5U_10U_1_land_3_lpi_1_dfm = ~((chn_inp_in_rsci_d_mxwt[309:300]!=10'b0000000000)
      | (~ IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_3_sva));
  assign IsNaN_5U_10U_1_land_3_lpi_1_dfm = IsDenorm_5U_10U_2_or_2_tmp & IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_3_sva;
  assign IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_3_sva = (chn_inp_in_rsci_d_mxwt[314:310]==5'b11111);
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_sva = ({1'b1 , (~ libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_23)})
      + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_2_if_1_if_acc_psp_sva[4:0];
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_lpi_1_dfm_3_mx0 = MUX_v_10_2_2((chn_inp_in_rsci_d_mxwt[325:316]),
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_or_12_mx0w1,
      or_dcpl_1015);
  assign IsZero_5U_10U_2_land_lpi_1_dfm = ~((chn_inp_in_rsci_d_mxwt[325:316]!=10'b0000000000)
      | (~ IsZero_5U_10U_2_IsZero_5U_10U_2_nor_cse_sva));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_FpExpoWidthInc_5U_6U_10U_1U_1U_1_nor_3_cse
      = ~(IsDenorm_5U_10U_2_land_lpi_1_dfm | IsInf_5U_10U_1_land_lpi_1_dfm);
  assign IsInf_5U_10U_1_land_lpi_1_dfm = ~((chn_inp_in_rsci_d_mxwt[325:316]!=10'b0000000000)
      | (~ IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_sva));
  assign IsNaN_5U_10U_1_land_lpi_1_dfm = IsDenorm_5U_10U_2_or_3_tmp & IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_sva;
  assign IsInf_5U_10U_1_IsInf_5U_10U_1_and_cse_sva = (chn_inp_in_rsci_d_mxwt[330:326]==5'b11111);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_9_0_1_lpi_1_dfm_2_mx0 = MUX_v_10_2_2(FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_9_0_1_lpi_1_dfm,
      10'b1111111111, IsInf_6U_23U_1_land_1_lpi_1_dfm_mx0w0);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_9_0_2_lpi_1_dfm_2_mx0 = MUX_v_10_2_2(FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_9_0_2_lpi_1_dfm,
      10'b1111111111, IsInf_6U_23U_1_land_2_lpi_1_dfm_mx0w0);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_9_0_3_lpi_1_dfm_2_mx0 = MUX_v_10_2_2(FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_9_0_3_lpi_1_dfm,
      10'b1111111111, IsInf_6U_23U_1_land_3_lpi_1_dfm_mx0w0);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_9_0_lpi_1_dfm_2_mx0 = MUX_v_10_2_2(FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_9_0_lpi_1_dfm,
      10'b1111111111, IsInf_6U_23U_1_land_lpi_1_dfm_mx0w0);
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_1_sva = ({1'b1 , (~ libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_24)})
      + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_1_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_1_sva[4:0];
  assign IsZero_5U_10U_land_1_lpi_1_dfm = ~((chn_inp_in_rsci_d_mxwt[405:396]!=10'b0000000000)
      | (~ IsZero_5U_10U_IsZero_5U_10U_nor_cse_1_sva));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_cse =
      ~(IsDenorm_5U_10U_land_1_lpi_1_dfm | IsInf_5U_10U_land_1_lpi_1_dfm);
  assign IsInf_5U_10U_land_1_lpi_1_dfm = ~((chn_inp_in_rsci_d_mxwt[405:396]!=10'b0000000000)
      | (~ IsInf_5U_10U_IsInf_5U_10U_and_cse_1_sva));
  assign IsNaN_5U_10U_land_1_lpi_1_dfm = IsDenorm_5U_10U_or_tmp & IsInf_5U_10U_IsInf_5U_10U_and_cse_1_sva;
  assign IsInf_5U_10U_IsInf_5U_10U_and_cse_1_sva = (chn_inp_in_rsci_d_mxwt[410:406]==5'b11111);
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_2_sva = ({1'b1 , (~ libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_25)})
      + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_2_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_2_sva[4:0];
  assign IsZero_5U_10U_land_2_lpi_1_dfm = ~((chn_inp_in_rsci_d_mxwt[421:412]!=10'b0000000000)
      | (~ IsZero_5U_10U_IsZero_5U_10U_nor_cse_2_sva));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_1_cse
      = ~(IsDenorm_5U_10U_land_2_lpi_1_dfm | IsInf_5U_10U_land_2_lpi_1_dfm);
  assign IsInf_5U_10U_land_2_lpi_1_dfm = ~((chn_inp_in_rsci_d_mxwt[421:412]!=10'b0000000000)
      | (~ IsInf_5U_10U_IsInf_5U_10U_and_cse_2_sva));
  assign IsNaN_5U_10U_land_2_lpi_1_dfm = IsDenorm_5U_10U_or_1_tmp & IsInf_5U_10U_IsInf_5U_10U_and_cse_2_sva;
  assign IsInf_5U_10U_IsInf_5U_10U_and_cse_2_sva = (chn_inp_in_rsci_d_mxwt[426:422]==5'b11111);
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_3_sva = ({1'b1 , (~ libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_26)})
      + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_3_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_3_sva[4:0];
  assign IsZero_5U_10U_land_3_lpi_1_dfm = ~((chn_inp_in_rsci_d_mxwt[437:428]!=10'b0000000000)
      | (~ IsZero_5U_10U_IsZero_5U_10U_nor_cse_3_sva));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_2_cse
      = ~(IsDenorm_5U_10U_land_3_lpi_1_dfm | IsInf_5U_10U_land_3_lpi_1_dfm);
  assign IsInf_5U_10U_land_3_lpi_1_dfm = ~((chn_inp_in_rsci_d_mxwt[437:428]!=10'b0000000000)
      | (~ IsInf_5U_10U_IsInf_5U_10U_and_cse_3_sva));
  assign IsNaN_5U_10U_land_3_lpi_1_dfm = IsDenorm_5U_10U_or_2_tmp & IsInf_5U_10U_IsInf_5U_10U_and_cse_3_sva;
  assign IsInf_5U_10U_IsInf_5U_10U_and_cse_3_sva = (chn_inp_in_rsci_d_mxwt[442:438]==5'b11111);
  assign nl_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_sva = ({1'b1 , (~ libraries_leading_sign_10_0_bc3b8703c8646a1ec2f1fe7a31faeefe3d5a_27)})
      + 5'b10001;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_sva = nl_FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_acc_psp_sva[4:0];
  assign IsZero_5U_10U_land_lpi_1_dfm = ~((chn_inp_in_rsci_d_mxwt[453:444]!=10'b0000000000)
      | (~ IsZero_5U_10U_IsZero_5U_10U_nor_cse_sva));
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_nor_3_cse
      = ~(IsDenorm_5U_10U_land_lpi_1_dfm | IsInf_5U_10U_land_lpi_1_dfm);
  assign IsInf_5U_10U_land_lpi_1_dfm = ~((chn_inp_in_rsci_d_mxwt[453:444]!=10'b0000000000)
      | (~ IsInf_5U_10U_IsInf_5U_10U_and_cse_sva));
  assign IsNaN_5U_10U_land_lpi_1_dfm = IsDenorm_5U_10U_or_3_tmp & IsInf_5U_10U_IsInf_5U_10U_and_cse_sva;
  assign IsInf_5U_10U_IsInf_5U_10U_and_cse_sva = (chn_inp_in_rsci_d_mxwt[458:454]==5'b11111);
  assign nl_inp_lookup_1_IntSaturation_51U_32U_else_if_acc_nl = conv_s2u_2_3(inp_lookup_if_else_o_acc_psp_1_sva[32:31])
      + 3'b1;
  assign inp_lookup_1_IntSaturation_51U_32U_else_if_acc_nl = nl_inp_lookup_1_IntSaturation_51U_32U_else_if_acc_nl[2:0];
  assign inp_lookup_1_IntSaturation_51U_32U_else_if_acc_itm_2_1 = readslicef_3_1_2((inp_lookup_1_IntSaturation_51U_32U_else_if_acc_nl));
  assign nl_inp_lookup_2_IntSaturation_51U_32U_else_if_acc_nl = conv_s2u_2_3(inp_lookup_if_else_o_acc_psp_2_sva[32:31])
      + 3'b1;
  assign inp_lookup_2_IntSaturation_51U_32U_else_if_acc_nl = nl_inp_lookup_2_IntSaturation_51U_32U_else_if_acc_nl[2:0];
  assign inp_lookup_2_IntSaturation_51U_32U_else_if_acc_itm_2_1 = readslicef_3_1_2((inp_lookup_2_IntSaturation_51U_32U_else_if_acc_nl));
  assign nl_inp_lookup_3_IntSaturation_51U_32U_else_if_acc_nl = conv_s2u_2_3(inp_lookup_if_else_o_acc_psp_3_sva[32:31])
      + 3'b1;
  assign inp_lookup_3_IntSaturation_51U_32U_else_if_acc_nl = nl_inp_lookup_3_IntSaturation_51U_32U_else_if_acc_nl[2:0];
  assign inp_lookup_3_IntSaturation_51U_32U_else_if_acc_itm_2_1 = readslicef_3_1_2((inp_lookup_3_IntSaturation_51U_32U_else_if_acc_nl));
  assign nl_inp_lookup_4_IntSaturation_51U_32U_else_if_acc_nl = conv_s2u_2_3(inp_lookup_if_else_o_acc_psp_sva[32:31])
      + 3'b1;
  assign inp_lookup_4_IntSaturation_51U_32U_else_if_acc_nl = nl_inp_lookup_4_IntSaturation_51U_32U_else_if_acc_nl[2:0];
  assign inp_lookup_4_IntSaturation_51U_32U_else_if_acc_itm_2_1 = readslicef_3_1_2((inp_lookup_4_IntSaturation_51U_32U_else_if_acc_nl));
  assign nl_inp_lookup_1_else_else_b0_mul_nl = $signed((chn_inp_in_crt_sva_1_331_268_1[15:0]))
      * $signed(conv_u2s_36_37({reg_inp_lookup_1_else_else_a0_acc_reg , reg_inp_lookup_1_else_else_a0_acc_1_reg
      , reg_inp_lookup_1_else_else_a0_acc_2_reg}));
  assign inp_lookup_1_else_else_b0_mul_nl = nl_inp_lookup_1_else_else_b0_mul_nl[51:0];
  assign nl_inp_lookup_else_else_o_acc_psp_1_sva = conv_s2s_52_53(inp_lookup_1_else_else_b0_mul_nl)
      + conv_s2s_51_53(inp_lookup_1_else_else_b1_mul_itm_2);
  assign inp_lookup_else_else_o_acc_psp_1_sva = nl_inp_lookup_else_else_o_acc_psp_1_sva[52:0];
  assign nl_inp_lookup_2_else_else_b0_mul_nl = $signed((chn_inp_in_crt_sva_1_331_268_1[31:16]))
      * $signed(conv_u2s_36_37({reg_inp_lookup_2_else_else_a0_acc_reg , reg_inp_lookup_2_else_else_a0_acc_1_reg
      , reg_inp_lookup_2_else_else_a0_acc_2_reg}));
  assign inp_lookup_2_else_else_b0_mul_nl = nl_inp_lookup_2_else_else_b0_mul_nl[51:0];
  assign nl_inp_lookup_else_else_o_acc_psp_2_sva = conv_s2s_52_53(inp_lookup_2_else_else_b0_mul_nl)
      + conv_s2s_51_53(inp_lookup_2_else_else_b1_mul_itm_2);
  assign inp_lookup_else_else_o_acc_psp_2_sva = nl_inp_lookup_else_else_o_acc_psp_2_sva[52:0];
  assign nl_inp_lookup_3_else_else_b0_mul_nl = $signed((chn_inp_in_crt_sva_1_331_268_1[47:32]))
      * $signed(conv_u2s_36_37({reg_inp_lookup_3_else_else_a0_acc_reg , reg_inp_lookup_3_else_else_a0_acc_1_reg
      , reg_inp_lookup_3_else_else_a0_acc_2_reg}));
  assign inp_lookup_3_else_else_b0_mul_nl = nl_inp_lookup_3_else_else_b0_mul_nl[51:0];
  assign nl_inp_lookup_else_else_o_acc_psp_3_sva = conv_s2s_52_53(inp_lookup_3_else_else_b0_mul_nl)
      + conv_s2s_51_53(inp_lookup_3_else_else_b1_mul_itm_2);
  assign inp_lookup_else_else_o_acc_psp_3_sva = nl_inp_lookup_else_else_o_acc_psp_3_sva[52:0];
  assign nl_inp_lookup_4_else_else_b0_mul_nl = $signed((chn_inp_in_crt_sva_1_331_268_1[63:48]))
      * $signed(conv_u2s_36_37({reg_inp_lookup_4_else_else_a0_acc_reg , reg_inp_lookup_4_else_else_a0_acc_1_reg
      , reg_inp_lookup_4_else_else_a0_acc_2_reg}));
  assign inp_lookup_4_else_else_b0_mul_nl = nl_inp_lookup_4_else_else_b0_mul_nl[51:0];
  assign nl_inp_lookup_else_else_o_acc_psp_sva = conv_s2s_52_53(inp_lookup_4_else_else_b0_mul_nl)
      + conv_s2s_51_53(inp_lookup_4_else_else_b1_mul_itm_2);
  assign inp_lookup_else_else_o_acc_psp_sva = nl_inp_lookup_else_else_o_acc_psp_sva[52:0];
  assign inp_lookup_1_IsZero_6U_10U_5_IsZero_6U_10U_5_nor_2 = ~((chn_inp_in_rsci_d_mxwt[282])
      | FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_3_0_mx0w0 | (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_3_mx0w0!=4'b0000));
  assign inp_lookup_3_IsZero_6U_10U_5_IsZero_6U_10U_5_nor_2 = ~((chn_inp_in_rsci_d_mxwt[314])
      | FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_3_0_mx0w0 | (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_3_mx0w0!=4'b0000));
  assign nl_inp_lookup_1_FpNormalize_8U_49U_1_acc_nl = ({1'b1 , (~ reg_FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_7_1_itm)})
      + conv_u2s_6_9(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_12)
      + 9'b1;
  assign inp_lookup_1_FpNormalize_8U_49U_1_acc_nl = nl_inp_lookup_1_FpNormalize_8U_49U_1_acc_nl[8:0];
  assign FpNormalize_8U_49U_1_oelse_not_9 = ((FpAdd_8U_23U_1_int_mant_p1_1_sva_3[48:0]!=49'b0000000000000000000000000000000000000000000000000))
      & (readslicef_9_1_8((inp_lookup_1_FpNormalize_8U_49U_1_acc_nl)));
  assign nl_inp_lookup_2_FpNormalize_8U_49U_1_acc_nl = ({1'b1 , (~ reg_FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_7_1_itm)})
      + conv_u2s_6_9(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_13)
      + 9'b1;
  assign inp_lookup_2_FpNormalize_8U_49U_1_acc_nl = nl_inp_lookup_2_FpNormalize_8U_49U_1_acc_nl[8:0];
  assign FpNormalize_8U_49U_1_oelse_not_11 = ((FpAdd_8U_23U_1_int_mant_p1_2_sva_3[48:0]!=49'b0000000000000000000000000000000000000000000000000))
      & (readslicef_9_1_8((inp_lookup_2_FpNormalize_8U_49U_1_acc_nl)));
  assign nl_inp_lookup_3_FpNormalize_8U_49U_1_acc_nl = ({1'b1 , (~ reg_FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_7_1_itm)})
      + conv_u2s_6_9(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_14)
      + 9'b1;
  assign inp_lookup_3_FpNormalize_8U_49U_1_acc_nl = nl_inp_lookup_3_FpNormalize_8U_49U_1_acc_nl[8:0];
  assign FpNormalize_8U_49U_1_oelse_not_13 = ((FpAdd_8U_23U_1_int_mant_p1_3_sva_3[48:0]!=49'b0000000000000000000000000000000000000000000000000))
      & (readslicef_9_1_8((inp_lookup_3_FpNormalize_8U_49U_1_acc_nl)));
  assign nl_inp_lookup_4_FpNormalize_8U_49U_1_acc_nl = ({1'b1 , (~ reg_FpMul_6U_10U_2_o_mant_lpi_1_dfm_7_1_reg)})
      + conv_u2s_6_9(libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_15)
      + 9'b1;
  assign inp_lookup_4_FpNormalize_8U_49U_1_acc_nl = nl_inp_lookup_4_FpNormalize_8U_49U_1_acc_nl[8:0];
  assign FpNormalize_8U_49U_1_oelse_not_15 = ((FpAdd_8U_23U_1_int_mant_p1_sva_3[48:0]!=49'b0000000000000000000000000000000000000000000000000))
      & (readslicef_9_1_8((inp_lookup_4_FpNormalize_8U_49U_1_acc_nl)));
  assign FpAdd_6U_10U_1_asn_124 = inp_lookup_1_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1
      & (FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_4[23]);
  assign nl_inp_lookup_1_FpNormalize_6U_23U_1_acc_nl = ({1'b1 , (~ FpAdd_6U_10U_1_qr_2_lpi_1_dfm_5)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_8)
      + 7'b1;
  assign inp_lookup_1_FpNormalize_6U_23U_1_acc_nl = nl_inp_lookup_1_FpNormalize_6U_23U_1_acc_nl[6:0];
  assign FpNormalize_6U_23U_1_oelse_not_9 = FpNormalize_6U_23U_1_if_or_itm_2 & (readslicef_7_1_6((inp_lookup_1_FpNormalize_6U_23U_1_acc_nl)));
  assign FpAdd_6U_10U_1_asn_126 = inp_lookup_2_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1
      & (FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_4[23]);
  assign nl_inp_lookup_2_FpNormalize_6U_23U_1_acc_nl = ({1'b1 , (~ FpAdd_6U_10U_1_qr_3_lpi_1_dfm_5)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_9)
      + 7'b1;
  assign inp_lookup_2_FpNormalize_6U_23U_1_acc_nl = nl_inp_lookup_2_FpNormalize_6U_23U_1_acc_nl[6:0];
  assign FpNormalize_6U_23U_1_oelse_not_11 = FpNormalize_6U_23U_1_if_or_1_itm_2 &
      (readslicef_7_1_6((inp_lookup_2_FpNormalize_6U_23U_1_acc_nl)));
  assign FpAdd_6U_10U_1_asn_128 = inp_lookup_3_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1
      & (FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_4[23]);
  assign nl_inp_lookup_3_FpNormalize_6U_23U_1_acc_nl = ({1'b1 , (~ FpAdd_6U_10U_1_qr_4_lpi_1_dfm_5)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_10)
      + 7'b1;
  assign inp_lookup_3_FpNormalize_6U_23U_1_acc_nl = nl_inp_lookup_3_FpNormalize_6U_23U_1_acc_nl[6:0];
  assign FpNormalize_6U_23U_1_oelse_not_13 = FpNormalize_6U_23U_1_if_or_2_itm_2 &
      (readslicef_7_1_6((inp_lookup_3_FpNormalize_6U_23U_1_acc_nl)));
  assign FpAdd_6U_10U_1_asn_130 = inp_lookup_4_FpAdd_6U_10U_1_if_3_if_acc_1_itm_5_1
      & (FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_4[23]);
  assign nl_inp_lookup_4_FpNormalize_6U_23U_1_acc_nl = ({1'b1 , (~ FpAdd_6U_10U_1_qr_lpi_1_dfm_5)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_11)
      + 7'b1;
  assign inp_lookup_4_FpNormalize_6U_23U_1_acc_nl = nl_inp_lookup_4_FpNormalize_6U_23U_1_acc_nl[6:0];
  assign FpNormalize_6U_23U_1_oelse_not_15 = FpNormalize_6U_23U_1_if_or_3_itm_2 &
      (readslicef_7_1_6((inp_lookup_4_FpNormalize_6U_23U_1_acc_nl)));
  assign FpAdd_6U_10U_asn_87 = FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_1_sva_2
      & (FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_4[23]);
  assign FpAdd_6U_10U_asn_89 = FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_2_sva_2
      & (FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_4[23]);
  assign FpAdd_6U_10U_asn_91 = FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_3_sva_2
      & (FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_4[23]);
  assign FpAdd_6U_10U_asn_93 = FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_sva_2
      & (FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_4[23]);
  assign inp_lookup_asn_98 = inp_lookup_else_unequal_tmp_38 & (~ (chn_inp_in_crt_sva_12_739_736_1[3]));
  assign inp_lookup_asn_102 = inp_lookup_if_unequal_tmp_19 & (chn_inp_in_crt_sva_12_739_736_1[3]);
  assign inp_lookup_asn_106 = inp_lookup_else_unequal_tmp_38 & (~ (chn_inp_in_crt_sva_12_739_736_1[0]));
  assign inp_lookup_asn_110 = inp_lookup_if_unequal_tmp_19 & (chn_inp_in_crt_sva_12_739_736_1[0]);
  assign inp_lookup_asn_114 = inp_lookup_else_unequal_tmp_38 & (~ (chn_inp_in_crt_sva_12_739_736_1[2]));
  assign inp_lookup_asn_118 = inp_lookup_if_unequal_tmp_19 & (chn_inp_in_crt_sva_12_739_736_1[2]);
  assign inp_lookup_asn_122 = inp_lookup_else_unequal_tmp_38 & (~ (chn_inp_in_crt_sva_12_739_736_1[1]));
  assign inp_lookup_asn_126 = inp_lookup_if_unequal_tmp_19 & (chn_inp_in_crt_sva_12_739_736_1[1]);
  assign inp_lookup_3_IsZero_6U_10U_2_aif_IsZero_6U_10U_2_aelse_nor_2 = ~((FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_3_mx1!=10'b0000000000));
  assign inp_lookup_1_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_2 = ~((FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_1_lpi_1_dfm_3_mx0!=10'b0000000000));
  assign FpAdd_6U_10U_mux_50_tmp_23 = MUX_s_1_2_2((FpAdd_6U_10U_asn_mx0w1[23]), (FpAdd_6U_10U_int_mant_p1_sva[23]),
      reg_inp_lookup_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse);
  assign FpAdd_6U_10U_mux_34_tmp_23 = MUX_s_1_2_2((FpAdd_6U_10U_asn_17_mx0w1[23]),
      (FpAdd_6U_10U_int_mant_p1_3_sva[23]), reg_inp_lookup_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse);
  assign FpAdd_6U_10U_mux_18_tmp_23 = MUX_s_1_2_2((FpAdd_6U_10U_asn_20_mx0w1[23]),
      (FpAdd_6U_10U_int_mant_p1_2_sva[23]), reg_inp_lookup_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse);
  assign FpAdd_6U_10U_mux_2_tmp_23 = MUX_s_1_2_2((FpAdd_6U_10U_asn_23_mx0w1[23]),
      (FpAdd_6U_10U_int_mant_p1_1_sva[23]), reg_inp_lookup_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse);
  assign and_dcpl_21 = main_stage_v_7 & (chn_inp_in_crt_sva_7_739_736_1[1]) & (cfg_precision_1_sva_st_84[1]);
  assign and_dcpl_38 = or_11_cse & (chn_inp_in_rsci_d_mxwt[736]);
  assign and_dcpl_40 = (cfg_precision_rsci_d==2'b10) & chn_inp_in_rsci_bawt;
  assign or_2_cse = (cfg_precision_rsci_d!=2'b10);
  assign and_dcpl_42 = or_2_cse & chn_inp_in_rsci_bawt;
  assign and_dcpl_49 = or_11_cse & (chn_inp_in_rsci_d_mxwt[737]);
  assign and_dcpl_57 = or_11_cse & (chn_inp_in_rsci_d_mxwt[738]);
  assign and_dcpl_65 = or_11_cse & (chn_inp_in_rsci_d_mxwt[739]);
  assign or_tmp_6 = (~ chn_inp_in_rsci_bawt) | (cfg_precision_rsci_d!=2'b10);
  assign or_tmp_8 = (~ main_stage_v_1) | (cfg_precision_1_sva_st_90!=2'b10);
  assign not_tmp_34 = ~((chn_inp_in_rsci_d_mxwt[162:128]!=35'b00000000000000000000000000000000000));
  assign or_tmp_21 = (~ main_stage_v_1) | (chn_inp_in_crt_sva_1_739_395_1[341]) |
      (cfg_precision_1_sva_st_90!=2'b10);
  assign mux_81_itm = MUX_s_1_2_2(or_tmp_21, or_471_cse, or_11_cse);
  assign mux_tmp_6 = MUX_s_1_2_2(main_stage_v_1, chn_inp_in_rsci_bawt, or_11_cse);
  assign not_tmp_45 = ~((chn_inp_in_rsci_d_mxwt[197:163]!=35'b00000000000000000000000000000000000));
  assign or_tmp_52 = (~ main_stage_v_1) | (chn_inp_in_crt_sva_1_739_395_1[342]) |
      (cfg_precision_1_sva_st_90!=2'b10);
  assign mux_87_itm = MUX_s_1_2_2(or_tmp_52, or_763_cse, or_11_cse);
  assign or_tmp_85 = (chn_inp_in_crt_sva_1_739_395_1[343]) | (~ main_stage_v_1) |
      (cfg_precision_1_sva_st_90!=2'b10);
  assign mux_95_itm = MUX_s_1_2_2(or_tmp_85, or_802_cse, or_11_cse);
  assign not_tmp_69 = ~((chn_inp_in_rsci_d_mxwt[267:233]!=35'b00000000000000000000000000000000000));
  assign or_tmp_114 = (chn_inp_in_crt_sva_1_739_395_1[344]) | (~ main_stage_v_1)
      | (cfg_precision_1_sva_st_90!=2'b10);
  assign or_114_cse = (chn_inp_in_rsci_d_mxwt[739]) | (~ chn_inp_in_rsci_bawt) |
      (cfg_precision_rsci_d!=2'b10);
  assign mux_100_itm = MUX_s_1_2_2(or_tmp_114, or_114_cse, or_11_cse);
  assign and_3402_nl = (chn_inp_in_crt_sva_1_739_395_1[341]) & (cfg_precision_1_sva_st_90==2'b10);
  assign nor_1710_nl = ~((~ (chn_inp_in_crt_sva_1_739_395_1[341])) | (cfg_precision_1_sva_st_90!=2'b10));
  assign mux_106_nl = MUX_s_1_2_2((nor_1710_nl), (and_3402_nl), inp_lookup_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3);
  assign nand_tmp_3 = ~(main_stage_v_1 & (mux_106_nl));
  assign mux_115_itm = MUX_s_1_2_2(or_2176_cse, or_tmp_8, or_11_cse);
  assign or_178_cse = (~((FpFractionToFloat_35U_6U_10U_1_mux_tmp[4:3]==2'b11) & (IntLeadZero_35U_1_leading_sign_35_0_rtn_1_sva_2[5])
      & inp_lookup_1_FpMantRNE_36U_11U_1_else_and_svs_2 & (~ IsNaN_6U_10U_6_nor_tmp)))
      | (~(FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_st_2 & (FpFractionToFloat_35U_6U_10U_1_mux_tmp[2:0]==3'b111)));
  assign nor_5_cse = ~(or_5873_cse | (~ inp_lookup_1_FpMul_6U_10U_2_else_2_if_acc_itm_6));
  assign not_tmp_101 = ~((cfg_precision_1_sva_st_90[1]) & IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_13);
  assign mux_tmp_50 = MUX_s_1_2_2(main_stage_v_2, main_stage_v_1, or_11_cse);
  assign nand_tmp_5 = ~(main_stage_v_1 & (chn_inp_in_crt_sva_1_739_395_1[342]) &
      (~ or_2010_cse));
  assign or_tmp_213 = ~(main_stage_v_1 & (chn_inp_in_crt_sva_1_739_395_1[342]) &
      (cfg_precision_1_sva_st_90==2'b10));
  assign or_tmp_234 = (~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[1]) |
      (cfg_precision_1_sva_st_91!=2'b10);
  assign or_tmp_238 = (~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[1]) |
      (cfg_precision_1_sva_st_91!=2'b10) | (~ inp_lookup_2_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs)
      | FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_3;
  assign or_tmp_241 = (~(FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_st_2 & inp_lookup_2_FpMantRNE_36U_11U_1_else_and_svs_2
      & (IntLeadZero_35U_1_leading_sign_35_0_rtn_2_sva_2[5]) & (~ IsNaN_6U_10U_6_nor_1_tmp)))
      | (FpFractionToFloat_35U_6U_10U_1_mux_40_tmp!=5'b11111);
  assign nor_13_cse = ~(or_5890_cse | (~ inp_lookup_2_FpMul_6U_10U_2_else_2_if_acc_itm_6));
  assign not_tmp_126 = ~((cfg_precision_1_sva_st_90[1]) & IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_13);
  assign nand_tmp_8 = ~((chn_inp_in_crt_sva_1_739_395_1[343]) & main_stage_v_1 &
      nor_1336_cse_1);
  assign or_tmp_277 = ~((chn_inp_in_crt_sva_2_739_736_1[2]) & main_stage_v_2 & (cfg_precision_1_sva_st_91==2'b10));
  assign or_tmp_306 = (chn_inp_in_crt_sva_2_739_736_1[2]) | (~ main_stage_v_2) |
      (cfg_precision_1_sva_st_91!=2'b10);
  assign nand_616_cse = ~((FpFractionToFloat_35U_6U_10U_1_mux_41_tmp==5'b11111) &
      (IntLeadZero_35U_1_leading_sign_35_0_rtn_3_sva_2[5]) & inp_lookup_3_FpMantRNE_36U_11U_1_else_and_svs_2
      & (~ IsNaN_6U_10U_6_nor_2_tmp) & FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_st_2);
  assign not_tmp_152 = ~((cfg_precision_1_sva_st_90[1]) & IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_13);
  assign nand_tmp_12 = ~((chn_inp_in_crt_sva_1_739_395_1[344]) & main_stage_v_1 &
      nor_1336_cse_1);
  assign or_tmp_347 = ~((chn_inp_in_crt_sva_1_739_395_1[344]) & main_stage_v_1 &
      (cfg_precision_1_sva_st_90==2'b10));
  assign or_tmp_374 = (~ inp_lookup_4_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs)
      | FpMul_6U_10U_2_lor_1_lpi_1_dfm_st_3 | (~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[3])
      | (cfg_precision_1_sva_st_91!=2'b10);
  assign mux_197_itm = MUX_s_1_2_2(or_2282_cse, or_2176_cse, or_11_cse);
  assign or_tmp_439 = (cfg_precision_1_sva_st_91!=2'b10);
  assign and_tmp_29 = main_stage_v_2 & (chn_inp_in_crt_sva_2_739_736_1[0]) & or_tmp_439;
  assign or_tmp_440 = (cfg_precision_1_sva_st_80!=2'b10);
  assign not_tmp_182 = ~((cfg_precision_1_sva_st_80[1]) & (nor_1210_cse | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_15));
  assign nor_1640_nl = ~((cfg_precision_1_sva_st_80[0]) | not_tmp_182);
  assign mux_204_nl = MUX_s_1_2_2((nor_1640_nl), or_tmp_440, chn_inp_in_crt_sva_3_739_736_1[0]);
  assign and_tmp_33 = main_stage_v_3 & (mux_204_nl);
  assign mux_203_nl = MUX_s_1_2_2((~ or_tmp_439), or_tmp_439, chn_inp_in_crt_sva_2_739_736_1[0]);
  assign and_132_nl = main_stage_v_2 & (mux_203_nl);
  assign mux_tmp_127 = MUX_s_1_2_2(and_tmp_33, (and_132_nl), or_11_cse);
  assign or_454_nl = (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[0]) | (cfg_precision_1_sva_st_80[0])
      | not_tmp_182;
  assign mux_tmp_133 = MUX_s_1_2_2((or_454_nl), or_5800_cse, or_11_cse);
  assign or_tmp_461 = (~(FpMul_6U_10U_2_lor_6_lpi_1_dfm_st_4 | (~ inp_lookup_1_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4)
      | (~ inp_lookup_1_FpMul_6U_10U_2_else_2_else_slc_FpMul_6U_10U_2_p_mant_p1_21_itm_2)))
      | (chn_inp_in_crt_sva_3_739_736_1[0]) | (cfg_precision_1_sva_st_80!=2'b10);
  assign nand_tmp_14 = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ main_stage_v_3) | or_tmp_461;
  assign and_tmp_34 = main_stage_v_3 & or_tmp_461;
  assign or_tmp_463 = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ and_tmp_34);
  assign and_tmp_35 = main_stage_v_2 & (chn_inp_in_crt_sva_2_739_736_1[1]) & or_tmp_439;
  assign or_504_cse = (~ inp_lookup_2_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs)
      | FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_3;
  assign or_506_nl = (cfg_precision_1_sva_st_80!=2'b10) | (~ IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_15);
  assign mux_tmp_163 = MUX_s_1_2_2(or_tmp_440, (or_506_nl), or_504_cse);
  assign mux_242_nl = MUX_s_1_2_2((~ mux_tmp_163), or_tmp_440, chn_inp_in_crt_sva_3_739_736_1[1]);
  assign and_tmp_38 = main_stage_v_3 & (mux_242_nl);
  assign mux_240_nl = MUX_s_1_2_2((~ or_tmp_439), or_tmp_439, chn_inp_in_crt_sva_2_739_736_1[1]);
  assign and_138_nl = main_stage_v_2 & (mux_240_nl);
  assign mux_tmp_165 = MUX_s_1_2_2(and_tmp_38, (and_138_nl), or_11_cse);
  assign or_515_nl = (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[1]) | mux_tmp_163;
  assign mux_tmp_171 = MUX_s_1_2_2((or_515_nl), or_tmp_234, or_11_cse);
  assign or_tmp_523 = (~(FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_4 | (~ inp_lookup_2_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4)
      | (~ inp_lookup_2_FpMul_6U_10U_2_else_2_else_slc_FpMul_6U_10U_2_p_mant_p1_21_itm_2)))
      | (chn_inp_in_crt_sva_3_739_736_1[1]) | (cfg_precision_1_sva_st_80!=2'b10);
  assign nand_tmp_16 = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ main_stage_v_3) | or_tmp_523;
  assign and_tmp_39 = main_stage_v_3 & or_tmp_523;
  assign or_tmp_525 = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ and_tmp_39);
  assign and_tmp_42 = (chn_inp_in_crt_sva_2_739_736_1[2]) & main_stage_v_2 & or_tmp_439;
  assign or_570_nl = (cfg_precision_1_sva_st_80!=2'b10) | (~ IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_15);
  assign mux_tmp_201 = MUX_s_1_2_2(or_tmp_440, (or_570_nl), or_5372_cse);
  assign mux_280_nl = MUX_s_1_2_2((~ mux_tmp_201), or_tmp_440, chn_inp_in_crt_sva_3_739_736_1[2]);
  assign and_tmp_45 = main_stage_v_3 & (mux_280_nl);
  assign and_145_nl = main_stage_v_2 & or_tmp_439;
  assign mux_278_nl = MUX_s_1_2_2((~ or_2176_cse), (and_145_nl), chn_inp_in_crt_sva_2_739_736_1[2]);
  assign mux_tmp_203 = MUX_s_1_2_2(and_tmp_45, (mux_278_nl), or_11_cse);
  assign or_577_nl = (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[2]) | mux_tmp_201;
  assign mux_tmp_209 = MUX_s_1_2_2((or_577_nl), or_tmp_306, or_11_cse);
  assign or_tmp_584 = (~((~ IsNaN_6U_10U_5_land_3_lpi_1_dfm_5) | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_15))
      | (chn_inp_in_crt_sva_3_739_736_1[2]) | (cfg_precision_1_sva_st_80[0]) | (~((cfg_precision_1_sva_st_80[1])
      & or_5372_cse));
  assign and_tmp_48 = main_stage_v_3 & or_tmp_584;
  assign nand_tmp_18 = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ main_stage_v_3) | or_tmp_584;
  assign or_tmp_597 = (~(FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_4 | (~ inp_lookup_3_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4)
      | (~ inp_lookup_3_FpMul_6U_10U_2_else_2_else_slc_FpMul_6U_10U_2_p_mant_p1_21_itm_2)))
      | (chn_inp_in_crt_sva_3_739_736_1[2]) | (cfg_precision_1_sva_st_80!=2'b10);
  assign nand_tmp_20 = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ main_stage_v_3) | or_tmp_597;
  assign and_tmp_49 = main_stage_v_3 & or_tmp_597;
  assign or_tmp_599 = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ and_tmp_49);
  assign or_tmp_621 = ~((chn_inp_in_rsci_d_mxwt[739]) & chn_inp_in_rsci_bawt & (cfg_precision_rsci_d==2'b10));
  assign and_tmp_50 = main_stage_v_2 & (chn_inp_in_crt_sva_2_739_736_1[3]) & or_tmp_439;
  assign or_tmp_630 = (cfg_precision_1_sva_st_80!=2'b10) | (~ reg_chn_inp_out_rsci_ld_core_psct_cse)
      | chn_inp_out_rsci_bawt;
  assign or_tmp_631 = (~((cfg_precision_1_sva_st_80!=2'b10))) | (~ reg_chn_inp_out_rsci_ld_core_psct_cse)
      | chn_inp_out_rsci_bawt;
  assign mux_321_nl = MUX_s_1_2_2(or_tmp_631, or_tmp_630, chn_inp_in_crt_sva_3_739_736_1[3]);
  assign mux_322_nl = MUX_s_1_2_2(or_11_cse, (mux_321_nl), main_stage_v_3);
  assign or_635_nl = (~(FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_3 | (~ inp_lookup_4_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs)
      | (cfg_precision_1_sva_st_80!=2'b10))) | (~ reg_chn_inp_out_rsci_ld_core_psct_cse)
      | chn_inp_out_rsci_bawt;
  assign mux_323_nl = MUX_s_1_2_2((or_635_nl), or_tmp_630, chn_inp_in_crt_sva_3_739_736_1[3]);
  assign mux_324_nl = MUX_s_1_2_2(or_11_cse, (mux_323_nl), main_stage_v_3);
  assign mux_tmp_247 = MUX_s_1_2_2((mux_324_nl), (mux_322_nl), IsNaN_6U_10U_2_land_lpi_1_dfm_st_15);
  assign mux_326_nl = MUX_s_1_2_2(or_tmp_630, or_tmp_631, chn_inp_in_crt_sva_3_739_736_1[3]);
  assign nand_22_nl = ~(main_stage_v_3 & (~ (mux_326_nl)));
  assign or_636_nl = FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_3 | (~ inp_lookup_4_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs)
      | (cfg_precision_1_sva_st_80!=2'b10) | (~ reg_chn_inp_out_rsci_ld_core_psct_cse)
      | chn_inp_out_rsci_bawt;
  assign mux_327_nl = MUX_s_1_2_2((or_636_nl), or_tmp_631, chn_inp_in_crt_sva_3_739_736_1[3]);
  assign nand_23_nl = ~(main_stage_v_3 & (~ (mux_327_nl)));
  assign mux_tmp_250 = MUX_s_1_2_2((nand_23_nl), (nand_22_nl), IsNaN_6U_10U_2_land_lpi_1_dfm_st_15);
  assign and_3346_cse = (chn_inp_in_crt_sva_2_739_736_1[3]) & main_stage_v_2;
  assign mux_tmp_251 = MUX_s_1_2_2((~ mux_tmp_250), mux_tmp_247, and_3346_cse);
  assign or_645_nl = FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_3 | (~ inp_lookup_4_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs)
      | (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt;
  assign mux_337_nl = MUX_s_1_2_2((or_645_nl), or_11_cse, IsNaN_6U_10U_2_land_lpi_1_dfm_st_15);
  assign nand_tmp_24 = (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[3]) |
      (cfg_precision_1_sva_st_80!=2'b10) | (mux_337_nl);
  assign or_647_nl = IsNaN_6U_10U_2_land_lpi_1_dfm_st_15 | nor_572_cse | (~ reg_chn_inp_out_rsci_ld_core_psct_cse)
      | chn_inp_out_rsci_bawt;
  assign mux_tmp_260 = MUX_s_1_2_2(or_11_cse, (or_647_nl), nor_1800_cse);
  assign mux_339_nl = MUX_s_1_2_2(nand_tmp_24, (~ mux_tmp_260), inp_lookup_4_FpMul_6U_10U_1_else_2_if_acc_itm_6_1);
  assign mux_tmp_262 = MUX_s_1_2_2((mux_339_nl), nand_tmp_24, or_648_cse);
  assign nor_74_cse = ~((~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[3])
      | (cfg_precision_1_sva_st_91!=2'b10));
  assign mux_tmp_278 = MUX_s_1_2_2(main_stage_v_4, main_stage_v_3, or_11_cse);
  assign or_tmp_679 = (chn_inp_in_crt_sva_2_739_736_1[0]) | (cfg_precision_1_sva_st_91!=2'b10);
  assign not_tmp_282 = ~((cfg_precision_1_sva_st_80[1]) & IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_15);
  assign or_tmp_701 = (~((~ IsNaN_6U_10U_5_land_1_lpi_1_dfm_6) | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_16))
      | (chn_inp_in_crt_sva_4_739_736_1[0]) | (cfg_precision_1_sva_st_81!=2'b10);
  assign nand_tmp_29 = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ main_stage_v_4) | or_tmp_701;
  assign and_tmp_54 = main_stage_v_4 & or_tmp_701;
  assign or_tmp_704 = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ and_tmp_54);
  assign or_tmp_736 = (chn_inp_in_crt_sva_2_739_736_1[1]) | (cfg_precision_1_sva_st_91!=2'b10);
  assign or_tmp_753 = (~((~ IsNaN_6U_10U_5_land_2_lpi_1_dfm_6) | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_16))
      | (chn_inp_in_crt_sva_4_739_736_1[1]) | (cfg_precision_1_sva_st_81!=2'b10);
  assign nand_tmp_37 = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ main_stage_v_4) | or_tmp_753;
  assign and_tmp_56 = main_stage_v_4 & or_tmp_753;
  assign or_tmp_756 = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ and_tmp_56);
  assign not_tmp_345 = ~((cfg_precision_1_sva_st_81[1]) & IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_16);
  assign or_tmp_792 = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[2]) | (cfg_precision_1_sva_st_81[0])
      | not_tmp_345;
  assign not_tmp_346 = ~(main_stage_v_4 & ((chn_inp_in_crt_sva_4_739_736_1[2]) |
      (cfg_precision_1_sva_st_81[0]) | not_tmp_345));
  assign or_tmp_798 = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | not_tmp_346;
  assign or_tmp_808 = (~((~ IsNaN_6U_10U_5_land_3_lpi_1_dfm_6) | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_16))
      | (chn_inp_in_crt_sva_4_739_736_1[2]) | (cfg_precision_1_sva_st_81!=2'b10);
  assign nand_tmp_45 = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ main_stage_v_4) | or_tmp_808;
  assign and_tmp_59 = main_stage_v_4 & or_tmp_808;
  assign or_tmp_811 = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ and_tmp_59);
  assign nand_tmp_47 = ~(main_stage_v_4 & (~((~((chn_inp_in_crt_sva_4_739_736_1[3])
      | (~ FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_4))) | (cfg_precision_1_sva_st_81!=2'b10))));
  assign nand_tmp_50 = ~(main_stage_v_4 & (~(((chn_inp_in_crt_sva_4_739_736_1[3])
      & IsNaN_8U_23U_2_land_lpi_1_dfm_st_7) | (cfg_precision_1_sva_st_81!=2'b10))));
  assign not_tmp_374 = ~((cfg_precision_1_sva_st_82[1]) & main_stage_v_5);
  assign or_tmp_850 = (~ (chn_inp_in_crt_sva_5_739_736_1[0])) | (cfg_precision_1_sva_st_82[0])
      | not_tmp_374;
  assign or_tmp_880 = ~((chn_inp_in_crt_sva_5_739_736_1[1]) & (cfg_precision_1_sva_st_82==2'b10)
      & main_stage_v_5);
  assign nand_tmp_53 = ~(main_stage_v_4 & (~((~((chn_inp_in_crt_sva_4_739_736_1[2])
      | (~ FpAdd_6U_10U_1_is_a_greater_acc_2_itm_6))) | (cfg_precision_1_sva_st_81!=2'b10))));
  assign or_tmp_899 = ~((chn_inp_in_crt_sva_5_739_736_1[2]) & (cfg_precision_1_sva_st_82==2'b10)
      & main_stage_v_5);
  assign or_tmp_945 = (~ (chn_inp_in_crt_sva_5_739_736_1[3])) | (cfg_precision_1_sva_st_82[0])
      | not_tmp_374;
  assign or_tmp_957 = (cfg_precision_1_sva_st_82[0]) | not_tmp_374;
  assign or_tmp_959 = (cfg_precision_1_sva_st_83!=2'b10) | (~ main_stage_v_6);
  assign mux_516_itm = MUX_s_1_2_2(or_tmp_959, or_tmp_957, or_11_cse);
  assign not_tmp_424 = ~((chn_inp_in_crt_sva_6_739_736_1[0]) & main_stage_v_6);
  assign or_tmp_962 = (cfg_precision_1_sva_st_83!=2'b10) | not_tmp_424;
  assign or_968_nl = (~ inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5)
      | (cfg_precision_1_sva_st_82[0]) | not_tmp_374;
  assign or_970_nl = inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
      | (cfg_precision_1_sva_st_82[0]) | not_tmp_374;
  assign mux_tmp_441 = MUX_s_1_2_2((or_970_nl), (or_968_nl), inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6);
  assign mux_tmp_444 = MUX_s_1_2_2(mux_tmp_441, or_tmp_957, chn_inp_in_crt_sva_5_739_736_1[0]);
  assign not_tmp_428 = ~((cfg_precision_1_sva_st_83[1]) & (chn_inp_in_crt_sva_6_739_736_1[1])
      & main_stage_v_6);
  assign nand_570_cse = ~((cfg_precision_1_sva_st_83[1]) & main_stage_v_6);
  assign or_tmp_990 = (cfg_precision_1_sva_st_83[0]) | nand_570_cse;
  assign mux_530_itm = MUX_s_1_2_2(or_tmp_990, or_3167_cse, or_11_cse);
  assign or_tmp_992 = (cfg_precision_1_sva_st_83[0]) | not_tmp_428;
  assign nand_568_nl = ~(inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6
      & (cfg_precision_1_sva_st_82==2'b10) & main_stage_v_5);
  assign or_999_nl = inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6
      | (cfg_precision_1_sva_st_82!=2'b10) | (~ main_stage_v_5);
  assign mux_tmp_454 = MUX_s_1_2_2((or_999_nl), (nand_568_nl), inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5);
  assign mux_tmp_457 = MUX_s_1_2_2(mux_tmp_454, or_3167_cse, chn_inp_in_crt_sva_5_739_736_1[1]);
  assign mux_540_itm = MUX_s_1_2_2(or_tmp_959, or_3167_cse, or_11_cse);
  assign or_tmp_1009 = ~((chn_inp_in_crt_sva_6_739_736_1[2]) & (cfg_precision_1_sva_st_83==2'b10)
      & main_stage_v_6);
  assign mux_502_nl = MUX_s_1_2_2((~ inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5),
      inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5,
      inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6);
  assign not_tmp_442 = ~(main_stage_v_5 & (mux_502_nl));
  assign nand_566_nl = ~(IsNaN_8U_23U_3_land_3_lpi_1_dfm_7 & (cfg_precision_1_sva_st_83==2'b10)
      & main_stage_v_6);
  assign or_1018_nl = IsNaN_8U_23U_3_land_3_lpi_1_dfm_7 | (cfg_precision_1_sva_st_83!=2'b10)
      | (~ main_stage_v_6);
  assign mux_tmp_465 = MUX_s_1_2_2((or_1018_nl), (nand_566_nl), IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_itm_11);
  assign or_1022_nl = (cfg_precision_1_sva_st_82!=2'b10) | not_tmp_442;
  assign mux_tmp_467 = MUX_s_1_2_2((or_1022_nl), or_3167_cse, chn_inp_in_crt_sva_5_739_736_1[2]);
  assign or_tmp_1038 = ~((chn_inp_in_crt_sva_6_739_736_1[3]) & (cfg_precision_1_sva_st_83==2'b10)
      & main_stage_v_6);
  assign or_1043_nl = (~ inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5)
      | (cfg_precision_1_sva_st_82[0]) | not_tmp_374;
  assign or_1045_nl = inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
      | (cfg_precision_1_sva_st_82[0]) | not_tmp_374;
  assign mux_tmp_475 = MUX_s_1_2_2((or_1045_nl), (or_1043_nl), inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5);
  assign mux_tmp_478 = MUX_s_1_2_2(mux_tmp_475, or_tmp_957, chn_inp_in_crt_sva_5_739_736_1[3]);
  assign or_tmp_1058 = ~((chn_inp_in_crt_sva_7_739_736_1[0]) & (cfg_precision_1_sva_st_84==2'b10)
      & main_stage_v_7);
  assign mux_559_itm = MUX_s_1_2_2(or_tmp_1058, or_tmp_962, or_11_cse);
  assign or_tmp_1060 = IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_tmp | IsNaN_8U_23U_4_nor_tmp;
  assign nor_tmp_139 = (chn_inp_in_crt_sva_6_739_736_1[0]) & inp_lookup_1_FpMantRNE_24U_11U_else_and_svs;
  assign or_tmp_1098 = (cfg_precision_1_sva_st_83!=2'b10) | (chn_inp_in_crt_sva_6_739_736_1[0])
      | (~ main_stage_v_6);
  assign or_tmp_1106 = (cfg_precision_1_sva_st_84[0]) | (~ and_dcpl_21);
  assign mux_573_itm = MUX_s_1_2_2(or_tmp_1106, or_tmp_992, or_11_cse);
  assign nor_tmp_146 = (chn_inp_in_crt_sva_6_739_736_1[1]) & inp_lookup_2_FpMantRNE_24U_11U_else_and_svs;
  assign or_tmp_1143 = (cfg_precision_1_sva_st_83!=2'b10) | (chn_inp_in_crt_sva_6_739_736_1[1])
      | (~ main_stage_v_6);
  assign nand_557_cse = ~((cfg_precision_1_sva_st_84[1]) & main_stage_v_7);
  assign or_tmp_1147 = (cfg_precision_1_sva_st_84[0]) | nand_557_cse;
  assign mux_586_itm = MUX_s_1_2_2(or_tmp_1147, or_tmp_990, or_11_cse);
  assign or_tmp_1151 = ~((chn_inp_in_crt_sva_7_739_736_1[2]) & (cfg_precision_1_sva_st_84==2'b10)
      & main_stage_v_7);
  assign mux_587_itm = MUX_s_1_2_2(or_tmp_1151, or_tmp_1009, or_11_cse);
  assign or_tmp_1182 = (cfg_precision_1_sva_st_84!=2'b10) | (~ main_stage_v_7);
  assign or_tmp_1185 = (chn_inp_in_crt_sva_6_739_736_1[2]) | (cfg_precision_1_sva_st_83!=2'b10)
      | (~ main_stage_v_6);
  assign or_tmp_1198 = ~((chn_inp_in_crt_sva_7_739_736_1[3]) & (cfg_precision_1_sva_st_84==2'b10)
      & main_stage_v_7);
  assign mux_599_itm = MUX_s_1_2_2(or_tmp_1198, or_tmp_1038, or_11_cse);
  assign or_tmp_1232 = (chn_inp_in_crt_sva_7_739_736_1[3]) | (cfg_precision_1_sva_st_84!=2'b10)
      | (~ main_stage_v_7);
  assign or_tmp_1239 = (chn_inp_in_crt_sva_6_739_736_1[3]) | (cfg_precision_1_sva_st_83!=2'b10)
      | (~ main_stage_v_6);
  assign or_tmp_1253 = (~ (chn_inp_in_crt_sva_8_739_736_1[0])) | (cfg_precision_1_sva_st_85!=2'b10)
      | (~(IsNaN_6U_10U_land_1_lpi_1_dfm_5 & main_stage_v_8));
  assign or_tmp_1255 = ~((chn_inp_in_crt_sva_8_739_736_1[0]) & (cfg_precision_1_sva_st_85==2'b10)
      & main_stage_v_8);
  assign nor_tmp_161 = (chn_inp_in_crt_sva_7_739_736_1[0]) & FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_tmp;
  assign or_1280_nl = (cfg_precision_1_sva_st_85!=2'b10) | (~ main_stage_v_8);
  assign mux_623_itm = MUX_s_1_2_2((or_1280_nl), or_tmp_1182, or_11_cse);
  assign nor_tmp_166 = FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_2_tmp & (chn_inp_in_crt_sva_7_739_736_1[1]);
  assign not_tmp_537 = ~((cfg_precision_1_sva_st_85[1]) & (chn_inp_in_crt_sva_8_739_736_1[1])
      & main_stage_v_8);
  assign or_tmp_1302 = (cfg_precision_1_sva_st_85[0]) | not_tmp_537;
  assign nand_544_cse = ~((cfg_precision_1_sva_st_85[1]) & main_stage_v_8);
  assign or_1306_nl = (cfg_precision_1_sva_st_85[0]) | nand_544_cse;
  assign mux_632_itm = MUX_s_1_2_2((or_1306_nl), or_tmp_1147, or_11_cse);
  assign or_tmp_1310 = ~((chn_inp_in_crt_sva_8_739_736_1[2]) & IsNaN_6U_10U_land_3_lpi_1_dfm_5
      & (cfg_precision_1_sva_st_85==2'b10) & main_stage_v_8);
  assign or_tmp_1312 = ~((chn_inp_in_crt_sva_8_739_736_1[2]) & (cfg_precision_1_sva_st_85==2'b10)
      & main_stage_v_8);
  assign nor_tmp_172 = (chn_inp_in_crt_sva_7_739_736_1[2]) & FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_4_tmp;
  assign and_3289_nl = (~(inp_lookup_3_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp
      & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_12_1_1 & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_12_0_1
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_21==4'b1111))) & nor_tmp_172;
  assign mux_636_nl = MUX_s_1_2_2((and_3289_nl), nor_tmp_172, IsNaN_6U_10U_IsNaN_6U_10U_nor_2_tmp);
  assign nor_1476_nl = ~((~ (cfg_precision_1_sva_st_84[1])) | (~ main_stage_v_7)
      | (cfg_precision_1_sva_st_84[0]) | (mux_636_nl));
  assign nor_1477_nl = ~((chn_inp_in_crt_sva_8_739_736_1[2]) | (~ main_stage_v_8)
      | (cfg_precision_1_sva_st_85!=2'b10));
  assign mux_637_nl = MUX_s_1_2_2(nor_1493_cse, (nor_1477_nl), reg_FpMul_6U_10U_lor_5_lpi_1_dfm_3_cse);
  assign or_1319_nl = (~ IsNaN_6U_10U_1_land_3_lpi_1_dfm_5) | IsNaN_6U_10U_land_3_lpi_1_dfm_5;
  assign mux_638_nl = MUX_s_1_2_2(nor_1493_cse, (mux_637_nl), or_1319_nl);
  assign not_tmp_546 = MUX_s_1_2_2((mux_638_nl), (nor_1476_nl), or_11_cse);
  assign or_tmp_1338 = ~((chn_inp_in_crt_sva_8_739_736_1[3]) & IsNaN_6U_10U_land_lpi_1_dfm_5
      & (cfg_precision_1_sva_st_85==2'b10) & main_stage_v_8);
  assign or_tmp_1340 = ~((chn_inp_in_crt_sva_8_739_736_1[3]) & (cfg_precision_1_sva_st_85==2'b10)
      & main_stage_v_8);
  assign nor_tmp_176 = (chn_inp_in_crt_sva_7_739_736_1[3]) & FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_6_tmp;
  assign or_tmp_1363 = IsNaN_6U_10U_1_land_1_lpi_1_dfm_5 | IsNaN_6U_10U_land_1_lpi_1_dfm_5;
  assign or_tmp_1369 = IsNaN_6U_10U_land_1_lpi_1_dfm_6 | IsNaN_6U_10U_1_land_1_lpi_1_dfm_6;
  assign or_tmp_1389 = ~((chn_inp_in_crt_sva_9_739_736_1[0]) & main_stage_v_9 & (cfg_precision_1_sva_st_86==2'b10));
  assign mux_659_itm = MUX_s_1_2_2(or_tmp_1389, or_tmp_1255, or_11_cse);
  assign or_tmp_1393 = IsNaN_6U_10U_1_land_2_lpi_1_dfm_5 | IsNaN_6U_10U_land_2_lpi_1_dfm_5;
  assign or_tmp_1399 = IsNaN_6U_10U_land_2_lpi_1_dfm_6 | IsNaN_6U_10U_1_land_2_lpi_1_dfm_6;
  assign or_tmp_1418 = ~((chn_inp_in_crt_sva_9_739_736_1[1]) & main_stage_v_9 & (cfg_precision_1_sva_st_100==2'b10));
  assign mux_666_itm = MUX_s_1_2_2(or_tmp_1418, or_tmp_1302, or_11_cse);
  assign or_tmp_1422 = IsNaN_6U_10U_1_land_3_lpi_1_dfm_5 | IsNaN_6U_10U_land_3_lpi_1_dfm_5;
  assign or_tmp_1428 = IsNaN_6U_10U_land_3_lpi_1_dfm_6 | IsNaN_6U_10U_1_land_3_lpi_1_dfm_6;
  assign or_tmp_1444 = ~((chn_inp_in_crt_sva_9_739_736_1[2]) & main_stage_v_9 & (cfg_precision_1_sva_st_112==2'b10));
  assign mux_673_itm = MUX_s_1_2_2(or_tmp_1444, or_tmp_1312, or_11_cse);
  assign or_tmp_1448 = IsNaN_6U_10U_1_land_lpi_1_dfm_5 | IsNaN_6U_10U_land_lpi_1_dfm_5;
  assign or_tmp_1454 = IsNaN_6U_10U_land_lpi_1_dfm_6 | IsNaN_6U_10U_1_land_lpi_1_dfm_6;
  assign or_tmp_1467 = ~((chn_inp_in_crt_sva_9_739_736_1[3]) & main_stage_v_9 & (cfg_precision_1_sva_st_124==2'b10));
  assign mux_680_itm = MUX_s_1_2_2(or_tmp_1467, or_tmp_1340, or_11_cse);
  assign or_tmp_1502 = (~ (chn_inp_in_crt_sva_10_739_736_1[0])) | (cfg_precision_1_sva_st_87[0])
      | nand_653_cse;
  assign nor_tmp_199 = (chn_inp_in_crt_sva_10_739_736_1[0]) & main_stage_v_10;
  assign or_tmp_1537 = (~ (chn_inp_in_crt_sva_10_739_736_1[1])) | (cfg_precision_1_sva_st_101[0])
      | nand_652_cse;
  assign nor_tmp_208 = (chn_inp_in_crt_sva_10_739_736_1[1]) & main_stage_v_10;
  assign nor_tmp_216 = (chn_inp_in_crt_sva_10_739_736_1[2]) & main_stage_v_10;
  assign nor_tmp_224 = (chn_inp_in_crt_sva_10_739_736_1[3]) & main_stage_v_10;
  assign not_tmp_698 = ~((cfg_precision_1_sva_st_88[1]) & main_stage_v_11);
  assign nor_tmp_227 = (chn_inp_in_crt_sva_11_739_736_1[0]) & main_stage_v_11;
  assign not_tmp_703 = ~((cfg_precision_1_sva_st_102[1]) & main_stage_v_11);
  assign nor_tmp_230 = (chn_inp_in_crt_sva_11_739_736_1[1]) & main_stage_v_11;
  assign not_tmp_708 = ~((cfg_precision_1_sva_st_114[1]) & main_stage_v_11);
  assign nor_tmp_232 = (chn_inp_in_crt_sva_11_739_736_1[2]) & main_stage_v_11;
  assign not_tmp_711 = ~((cfg_precision_1_sva_st_126[1]) & main_stage_v_11);
  assign nor_tmp_234 = (chn_inp_in_crt_sva_11_739_736_1[3]) & main_stage_v_11;
  assign mux_tmp_698 = MUX_s_1_2_2(main_stage_v_11, main_stage_v_10, or_11_cse);
  assign or_tmp_1661 = (~(FpAdd_6U_10U_mux_2_tmp_23 | (~ FpNormalize_6U_23U_if_FpNormalize_6U_23U_if_nand_tmp)))
      | (~ (chn_inp_in_crt_sva_11_739_736_1[0])) | (cfg_precision_1_sva_st_88[0])
      | not_tmp_698;
  assign or_tmp_1665 = inp_lookup_1_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2
      | reg_FpNormalize_6U_23U_lor_1_lpi_1_dfm_4_cse | (~ main_stage_v_12) | (~ (chn_inp_in_crt_sva_12_739_736_1[0]))
      | (cfg_precision_1_sva_st_89!=2'b10);
  assign or_tmp_1671 = ~(main_stage_v_12 & (chn_inp_in_crt_sva_12_739_736_1[0]) &
      (cfg_precision_1_sva_st_89==2'b10));
  assign mux_782_itm = MUX_s_1_2_2(or_tmp_1671, or_1621_cse, or_11_cse);
  assign or_tmp_1687 = (~(IsNaN_6U_10U_2_land_1_lpi_1_dfm_25 | IsNaN_6U_10U_3_land_1_lpi_1_dfm_7))
      | (~ (chn_inp_in_crt_sva_11_739_736_1[0])) | (cfg_precision_1_sva_st_88[0])
      | not_tmp_698;
  assign or_1686_nl = (~ IsNaN_6U_10U_2_land_1_lpi_1_dfm_25) | (~ (chn_inp_in_crt_sva_11_739_736_1[0]))
      | (cfg_precision_1_sva_st_88[0]) | not_tmp_698;
  assign mux_tmp_708 = MUX_s_1_2_2(or_tmp_1687, (or_1686_nl), IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_23);
  assign or_tmp_1690 = ~(main_stage_v_12 & IsNaN_6U_10U_2_land_1_lpi_1_dfm_26 & (chn_inp_in_crt_sva_12_739_736_1[0])
      & (cfg_precision_1_sva_st_89==2'b10));
  assign or_tmp_1697 = ~(inp_lookup_2_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2
      & main_stage_v_12 & (chn_inp_in_crt_sva_12_739_736_1[1]) & (cfg_precision_1_sva_st_103==2'b10));
  assign or_tmp_1699 = inp_lookup_2_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2
      | (~ main_stage_v_12) | reg_FpNormalize_6U_23U_lor_2_lpi_1_dfm_4_cse | (~ (chn_inp_in_crt_sva_12_739_736_1[1]))
      | (cfg_precision_1_sva_st_103!=2'b10);
  assign or_tmp_1701 = ~(main_stage_v_12 & (chn_inp_in_crt_sva_12_739_736_1[1]) &
      (cfg_precision_1_sva_st_103==2'b10));
  assign mux_tmp_715 = MUX_s_1_2_2(or_tmp_1699, or_tmp_1701, FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_4[23]);
  assign mux_799_itm = MUX_s_1_2_2(or_tmp_1701, or_1632_cse, or_11_cse);
  assign or_tmp_1724 = IsNaN_6U_10U_2_land_2_lpi_1_dfm_25 | IsNaN_6U_10U_3_land_2_lpi_1_dfm_7;
  assign or_tmp_1728 = ~(FpAdd_6U_10U_or_17_cse & main_stage_v_12 & (chn_inp_in_crt_sva_12_739_736_1[1])
      & (cfg_precision_1_sva_st_103==2'b10));
  assign or_tmp_1734 = (~(FpAdd_6U_10U_mux_34_tmp_23 | (~ FpNormalize_6U_23U_if_FpNormalize_6U_23U_if_nand_2_tmp)))
      | (~ (chn_inp_in_crt_sva_11_739_736_1[2])) | (cfg_precision_1_sva_st_114[0])
      | not_tmp_708;
  assign not_tmp_733 = ~((cfg_precision_1_sva_st_115[1]) & (chn_inp_in_crt_sva_12_739_736_1[2])
      & main_stage_v_12);
  assign or_tmp_1736 = (~(inp_lookup_3_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2
      | (~ FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_3_sva_2))) |
      (cfg_precision_1_sva_st_115[0]) | not_tmp_733;
  assign or_tmp_1741 = inp_lookup_3_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2
      | (cfg_precision_1_sva_st_115[0]) | not_tmp_733;
  assign or_1752_nl = (cfg_precision_1_sva_st_115[0]) | not_tmp_733;
  assign mux_816_itm = MUX_s_1_2_2((or_1752_nl), or_1645_cse, or_11_cse);
  assign or_tmp_1770 = IsNaN_6U_10U_2_land_3_lpi_1_dfm_25 | IsNaN_6U_10U_3_land_3_lpi_1_dfm_7;
  assign or_tmp_1774 = FpAdd_6U_10U_FpAdd_6U_10U_nor_9_m1c | (cfg_precision_1_sva_st_115[0])
      | not_tmp_733;
  assign or_tmp_1784 = inp_lookup_4_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2
      | reg_FpNormalize_6U_23U_lor_lpi_1_dfm_4_cse | (~ main_stage_v_12) | (~ (chn_inp_in_crt_sva_12_739_736_1[3]))
      | (cfg_precision_1_sva_st_127!=2'b10);
  assign or_tmp_1786 = ~(main_stage_v_12 & (chn_inp_in_crt_sva_12_739_736_1[3]) &
      (cfg_precision_1_sva_st_127==2'b10));
  assign mux_829_itm = MUX_s_1_2_2(or_tmp_1786, or_1658_cse, or_11_cse);
  assign or_tmp_1806 = (~(IsNaN_6U_10U_2_land_lpi_1_dfm_25 | IsNaN_6U_10U_3_land_lpi_1_dfm_7))
      | (~ (chn_inp_in_crt_sva_11_739_736_1[3])) | (cfg_precision_1_sva_st_126[0])
      | not_tmp_711;
  assign or_1805_nl = (~ IsNaN_6U_10U_2_land_lpi_1_dfm_25) | (~ (chn_inp_in_crt_sva_11_739_736_1[3]))
      | (cfg_precision_1_sva_st_126[0]) | not_tmp_711;
  assign mux_tmp_754 = MUX_s_1_2_2(or_tmp_1806, (or_1805_nl), IsNaN_6U_10U_2_land_lpi_1_dfm_st_22);
  assign or_tmp_1818 = (chn_inp_in_crt_sva_11_739_736_1[0]) | (~ main_stage_v_11);
  assign nor_tmp_250 = inp_lookup_if_unequal_tmp_19 & (chn_inp_in_crt_sva_12_739_736_1[0])
      & main_stage_v_12;
  assign or_tmp_1826 = (chn_inp_in_crt_sva_11_739_736_1[3]) | (~ main_stage_v_11);
  assign nor_tmp_252 = inp_lookup_if_unequal_tmp_19 & (chn_inp_in_crt_sva_12_739_736_1[3])
      & main_stage_v_12;
  assign or_tmp_1840 = (chn_inp_in_crt_sva_11_739_736_1[1]) | (~ main_stage_v_11);
  assign nor_tmp_253 = (chn_inp_in_crt_sva_11_739_736_1[1]) & inp_lookup_if_unequal_tmp_12
      & main_stage_v_11;
  assign or_tmp_1845 = (chn_inp_in_crt_sva_11_739_736_1[2]) | inp_lookup_else_unequal_tmp_37
      | (~ main_stage_v_11);
  assign or_tmp_1849 = (chn_inp_in_crt_sva_11_739_736_1[2]) | (~ main_stage_v_11);
  assign nor_tmp_256 = inp_lookup_if_unequal_tmp_19 & (chn_inp_in_crt_sva_12_739_736_1[2])
      & main_stage_v_12;
  assign or_tmp_1856 = (chn_inp_in_crt_sva_11_739_736_1[1]) | inp_lookup_else_unequal_tmp_37
      | (~ main_stage_v_11);
  assign not_tmp_772 = ~(IsNaN_6U_10U_7_land_1_lpi_1_dfm_6 | (~(FpMul_6U_10U_2_lor_6_lpi_1_dfm_6
      | (~(FpMul_6U_10U_2_FpMul_6U_10U_2_and_itm_2 & ((~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_2)
      | inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4))))));
  assign not_tmp_773 = ~((cfg_precision_1_sva_st_80[1]) & (IsNaN_6U_10U_6_land_1_lpi_1_dfm_5
      | not_tmp_772));
  assign nor_1382_nl = ~((chn_inp_in_crt_sva_3_739_736_1[0]) | (cfg_precision_1_sva_st_80!=2'b10)
      | IsNaN_6U_10U_6_land_1_lpi_1_dfm_5 | not_tmp_772);
  assign or_5698_nl = (chn_inp_in_crt_sva_3_739_736_1[0]) | (cfg_precision_1_sva_st_80[0])
      | not_tmp_773;
  assign or_1866_nl = FpMul_6U_10U_1_lor_6_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_15;
  assign mux_857_nl = MUX_s_1_2_2((or_5698_nl), (nor_1382_nl), or_1866_nl);
  assign nand_tmp_90 = ~(main_stage_v_3 & (mux_857_nl));
  assign not_tmp_776 = ~((~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[0])
      | (cfg_precision_1_sva_st_80[0]) | not_tmp_773);
  assign or_tmp_1891 = nor_884_cse | (chn_inp_in_crt_sva_3_739_736_1[0]) | (cfg_precision_1_sva_st_80[0])
      | (~((cfg_precision_1_sva_st_80[1]) & or_5369_cse));
  assign and_tmp_111 = main_stage_v_3 & or_tmp_1891;
  assign nand_tmp_91 = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ main_stage_v_3) | or_tmp_1891;
  assign nor_1371_cse = ~(FpMul_6U_10U_2_lor_7_lpi_1_dfm_6 | (~(FpMul_6U_10U_2_FpMul_6U_10U_2_and_16_itm_2
      & ((~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_2) |
      inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4))));
  assign not_tmp_789 = ~(IsNaN_6U_10U_7_land_2_lpi_1_dfm_6 | nor_1371_cse);
  assign not_tmp_790 = ~((cfg_precision_1_sva_st_80[1]) & (IsNaN_6U_10U_6_land_2_lpi_1_dfm_5
      | not_tmp_789));
  assign nor_1369_nl = ~((chn_inp_in_crt_sva_3_739_736_1[1]) | (cfg_precision_1_sva_st_80!=2'b10)
      | IsNaN_6U_10U_6_land_2_lpi_1_dfm_5 | not_tmp_789);
  assign or_5697_nl = (chn_inp_in_crt_sva_3_739_736_1[1]) | (cfg_precision_1_sva_st_80[0])
      | not_tmp_790;
  assign or_1904_nl = FpMul_6U_10U_1_lor_7_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_15;
  assign mux_874_nl = MUX_s_1_2_2((or_5697_nl), (nor_1369_nl), or_1904_nl);
  assign nand_tmp_94 = ~(main_stage_v_3 & (mux_874_nl));
  assign not_tmp_793 = ~((~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[1])
      | (cfg_precision_1_sva_st_80[0]) | not_tmp_790);
  assign or_tmp_1929 = nor_880_cse | (chn_inp_in_crt_sva_3_739_736_1[1]) | (cfg_precision_1_sva_st_80[0])
      | (~((cfg_precision_1_sva_st_80[1]) & or_504_cse));
  assign and_tmp_116 = main_stage_v_3 & or_tmp_1929;
  assign nand_tmp_95 = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ main_stage_v_3) | or_tmp_1929;
  assign not_tmp_806 = ~(IsNaN_6U_10U_7_land_3_lpi_1_dfm_6 | (~(FpMul_6U_10U_2_lor_8_lpi_1_dfm_6
      | (~(FpMul_6U_10U_2_FpMul_6U_10U_2_and_17_itm_2 & ((~ FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_2)
      | inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4))))));
  assign not_tmp_807 = ~((cfg_precision_1_sva_st_80[1]) & (IsNaN_6U_10U_6_land_3_lpi_1_dfm_5
      | not_tmp_806));
  assign nor_1356_nl = ~((chn_inp_in_crt_sva_3_739_736_1[2]) | (cfg_precision_1_sva_st_80!=2'b10)
      | IsNaN_6U_10U_6_land_3_lpi_1_dfm_5 | not_tmp_806);
  assign or_5696_nl = (chn_inp_in_crt_sva_3_739_736_1[2]) | (cfg_precision_1_sva_st_80[0])
      | not_tmp_807;
  assign or_1942_nl = FpMul_6U_10U_1_lor_8_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_15;
  assign mux_891_nl = MUX_s_1_2_2((or_5696_nl), (nor_1356_nl), or_1942_nl);
  assign nand_tmp_98 = ~(main_stage_v_3 & (mux_891_nl));
  assign not_tmp_810 = ~((~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[2])
      | (cfg_precision_1_sva_st_80[0]) | not_tmp_807);
  assign or_tmp_1967 = nor_875_cse | (chn_inp_in_crt_sva_3_739_736_1[3]) | (cfg_precision_1_sva_st_80[0])
      | (~((cfg_precision_1_sva_st_80[1]) & or_3779_cse));
  assign and_tmp_121 = main_stage_v_3 & or_tmp_1967;
  assign nand_tmp_99 = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ main_stage_v_3) | or_tmp_1967;
  assign or_1970_cse = (cfg_precision_1_sva_st_90!=2'b10) | (chn_inp_in_crt_sva_1_739_395_1[344]);
  assign or_tmp_2199 = inp_lookup_2_FpMantRNE_22U_11U_2_else_and_tmp | FpMul_6U_10U_2_lor_7_lpi_1_dfm_5;
  assign or_tmp_2234 = inp_lookup_3_FpMantRNE_22U_11U_2_else_and_tmp | FpMul_6U_10U_2_lor_8_lpi_1_dfm_5;
  assign not_tmp_940 = ~((cfg_precision_1_sva_st_80[1]) & mux_1015_cse);
  assign or_2361_nl = (~ inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4)
      | (cfg_precision_1_sva_st_80!=2'b10);
  assign or_2362_nl = inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4
      | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_tmp_950 = MUX_s_1_2_2((or_2362_nl), (or_2361_nl), inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4);
  assign or_2398_nl = (~ inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4)
      | (cfg_precision_1_sva_st_80!=2'b10);
  assign or_2399_nl = inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4
      | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_tmp_966 = MUX_s_1_2_2((or_2399_nl), (or_2398_nl), inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4);
  assign or_2400_nl = (~ inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5)
      | (cfg_precision_1_sva_st_81!=2'b10);
  assign or_2401_nl = inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5
      | (cfg_precision_1_sva_st_81!=2'b10);
  assign mux_tmp_967 = MUX_s_1_2_2((or_2401_nl), (or_2400_nl), inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5);
  assign nor_1175_nl = ~((~ inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4)
      | (cfg_precision_1_sva_st_81!=2'b10));
  assign nor_1176_nl = ~(inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4
      | (cfg_precision_1_sva_st_81!=2'b10));
  assign mux_1057_nl = MUX_s_1_2_2((nor_1176_nl), (nor_1175_nl), inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5);
  assign nand_tmp_126 = ~(main_stage_v_4 & (chn_inp_in_crt_sva_4_739_736_1[3]) &
      (mux_1057_nl));
  assign or_tmp_2441 = IsNaN_6U_10U_4_land_lpi_1_dfm_5 | IsNaN_6U_10U_5_land_lpi_1_dfm_6;
  assign mux_1066_itm = MUX_s_1_2_2(or_tmp_957, or_3850_cse, or_11_cse);
  assign mux_1067_itm = MUX_s_1_2_2(or_3167_cse, or_3850_cse, or_11_cse);
  assign or_tmp_2486 = (chn_inp_in_crt_sva_5_739_736_1[0]) | (cfg_precision_1_sva_st_82[0])
      | not_tmp_374;
  assign or_tmp_2490 = (chn_inp_in_crt_sva_5_739_736_1[1]) | (cfg_precision_1_sva_st_82!=2'b10)
      | (~ main_stage_v_5);
  assign or_tmp_2494 = (chn_inp_in_crt_sva_5_739_736_1[2]) | (cfg_precision_1_sva_st_82!=2'b10)
      | (~ main_stage_v_5);
  assign or_tmp_2498 = (chn_inp_in_crt_sva_5_739_736_1[3]) | (cfg_precision_1_sva_st_82[0])
      | not_tmp_374;
  assign or_2507_nl = nor_1593_cse | (chn_inp_in_crt_sva_5_739_736_1[0]) | IsNaN_8U_23U_3_land_1_lpi_1_dfm_6
      | IsNaN_6U_10U_8_land_1_lpi_1_dfm_6;
  assign or_2508_nl = (chn_inp_in_crt_sva_5_739_736_1[0]) | IsNaN_8U_23U_3_land_1_lpi_1_dfm_6
      | IsNaN_6U_10U_8_land_1_lpi_1_dfm_6;
  assign mux_tmp_1008 = MUX_s_1_2_2((or_2508_nl), (or_2507_nl), IsNaN_8U_23U_2_land_1_lpi_1_dfm_9);
  assign nor_1155_nl = ~((~ main_stage_v_4) | (cfg_precision_1_sva_st_81!=2'b10)
      | (~((chn_inp_in_crt_sva_4_739_736_1[0]) | IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_tmp
      | FpAdd_6U_10U_1_is_a_greater_acc_itm_6 | inp_lookup_1_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp
      | mux_476_cse)));
  assign or_2509_nl = inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
      | mux_tmp_1008;
  assign nand_135_nl = ~(inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
      & (~ mux_tmp_1008));
  assign mux_1087_nl = MUX_s_1_2_2((nand_135_nl), (or_2509_nl), inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6);
  assign nor_1157_nl = ~((cfg_precision_1_sva_st_82[0]) | (~((cfg_precision_1_sva_st_82[1])
      & main_stage_v_5 & (mux_1087_nl))));
  assign not_tmp_1029 = MUX_s_1_2_2((nor_1157_nl), (nor_1155_nl), or_11_cse);
  assign and_tmp_158 = IsNaN_8U_23U_2_land_1_lpi_1_dfm_9 & nor_1593_cse;
  assign or_2528_nl = (~ inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5)
      | (~ main_stage_v_5) | (chn_inp_in_crt_sva_5_739_736_1[0]) | (cfg_precision_1_sva_st_82!=2'b10);
  assign or_2530_nl = inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
      | (~ main_stage_v_5) | (chn_inp_in_crt_sva_5_739_736_1[0]) | (cfg_precision_1_sva_st_82!=2'b10);
  assign mux_tmp_1015 = MUX_s_1_2_2((or_2530_nl), (or_2528_nl), inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6);
  assign or_tmp_2531 = (~ main_stage_v_5) | (chn_inp_in_crt_sva_5_739_736_1[0]) |
      (cfg_precision_1_sva_st_82!=2'b10);
  assign or_2535_nl = (~ chn_inp_in_crt_sva_4_411_1) | (cfg_precision_1_sva_st_81!=2'b10);
  assign or_2536_nl = chn_inp_in_crt_sva_4_411_1 | (cfg_precision_1_sva_st_81!=2'b10);
  assign mux_1099_nl = MUX_s_1_2_2((or_2536_nl), (or_2535_nl), inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5);
  assign mux_1100_nl = MUX_s_1_2_2((mux_1099_nl), or_3379_cse, chn_inp_in_crt_sva_4_739_736_1[0]);
  assign nand_tmp_138 = ~(main_stage_v_4 & (~ (mux_1100_nl)));
  assign or_2544_nl = nor_1587_cse | (chn_inp_in_crt_sva_5_739_736_1[1]) | IsNaN_8U_23U_3_land_2_lpi_1_dfm_6
      | IsNaN_6U_10U_8_land_2_lpi_1_dfm_4;
  assign or_2545_nl = (chn_inp_in_crt_sva_5_739_736_1[1]) | IsNaN_8U_23U_3_land_2_lpi_1_dfm_6
      | IsNaN_6U_10U_8_land_2_lpi_1_dfm_4;
  assign mux_tmp_1025 = MUX_s_1_2_2((or_2545_nl), (or_2544_nl), IsNaN_8U_23U_2_land_2_lpi_1_dfm_9);
  assign nor_1147_nl = ~((~ main_stage_v_4) | (cfg_precision_1_sva_st_81!=2'b10)
      | (~((chn_inp_in_crt_sva_4_739_736_1[1]) | IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_1_tmp
      | FpAdd_6U_10U_1_is_a_greater_acc_1_itm_6 | inp_lookup_2_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp
      | mux_485_cse)));
  assign or_2546_nl = inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
      | mux_tmp_1025;
  assign nand_139_nl = ~(inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
      & (~ mux_tmp_1025));
  assign mux_1104_nl = MUX_s_1_2_2((nand_139_nl), (or_2546_nl), inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6);
  assign nor_1149_nl = ~((~ main_stage_v_5) | (cfg_precision_1_sva_st_82[0]) | (~((cfg_precision_1_sva_st_82[1])
      & (mux_1104_nl))));
  assign not_tmp_1046 = MUX_s_1_2_2((nor_1149_nl), (nor_1147_nl), or_11_cse);
  assign and_tmp_162 = IsNaN_8U_23U_2_land_2_lpi_1_dfm_9 & nor_1587_cse;
  assign or_2565_nl = (~ inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5)
      | (~ main_stage_v_5) | (chn_inp_in_crt_sva_5_739_736_1[1]) | (cfg_precision_1_sva_st_82!=2'b10);
  assign or_2567_nl = inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
      | (~ main_stage_v_5) | (chn_inp_in_crt_sva_5_739_736_1[1]) | (cfg_precision_1_sva_st_82!=2'b10);
  assign mux_tmp_1032 = MUX_s_1_2_2((or_2567_nl), (or_2565_nl), inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6);
  assign or_2572_nl = (~ chn_inp_in_crt_sva_4_427_1) | (cfg_precision_1_sva_st_81!=2'b10);
  assign or_2573_nl = chn_inp_in_crt_sva_4_427_1 | (cfg_precision_1_sva_st_81!=2'b10);
  assign mux_1116_nl = MUX_s_1_2_2((or_2573_nl), (or_2572_nl), inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5);
  assign mux_1117_nl = MUX_s_1_2_2((mux_1116_nl), or_3379_cse, chn_inp_in_crt_sva_4_739_736_1[1]);
  assign nand_tmp_142 = ~(main_stage_v_4 & (~ (mux_1117_nl)));
  assign or_2581_nl = nor_1584_cse | (chn_inp_in_crt_sva_5_739_736_1[2]) | IsNaN_8U_23U_3_land_3_lpi_1_dfm_6
      | IsNaN_6U_10U_8_land_3_lpi_1_dfm_4;
  assign or_2582_nl = (chn_inp_in_crt_sva_5_739_736_1[2]) | IsNaN_8U_23U_3_land_3_lpi_1_dfm_6
      | IsNaN_6U_10U_8_land_3_lpi_1_dfm_4;
  assign mux_tmp_1042 = MUX_s_1_2_2((or_2582_nl), (or_2581_nl), IsNaN_8U_23U_2_land_3_lpi_1_dfm_9);
  assign nor_1139_nl = ~((~ main_stage_v_4) | (cfg_precision_1_sva_st_81!=2'b10)
      | (~((chn_inp_in_crt_sva_4_739_736_1[2]) | IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_2_tmp
      | FpAdd_6U_10U_1_is_a_greater_acc_2_itm_6 | inp_lookup_3_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp
      | mux_500_cse)));
  assign or_2583_nl = inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
      | mux_tmp_1042;
  assign nand_143_nl = ~(inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
      & (~ mux_tmp_1042));
  assign mux_1121_nl = MUX_s_1_2_2((nand_143_nl), (or_2583_nl), inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6);
  assign nor_1141_nl = ~((~ main_stage_v_5) | (cfg_precision_1_sva_st_82[0]) | (~((cfg_precision_1_sva_st_82[1])
      & (mux_1121_nl))));
  assign not_tmp_1063 = MUX_s_1_2_2((nor_1141_nl), (nor_1139_nl), or_11_cse);
  assign and_tmp_166 = IsNaN_8U_23U_2_land_3_lpi_1_dfm_9 & nor_1584_cse;
  assign or_2602_nl = (~ inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5)
      | (~ main_stage_v_5) | (chn_inp_in_crt_sva_5_739_736_1[2]) | (cfg_precision_1_sva_st_82!=2'b10);
  assign or_2604_nl = inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
      | (~ main_stage_v_5) | (chn_inp_in_crt_sva_5_739_736_1[2]) | (cfg_precision_1_sva_st_82!=2'b10);
  assign mux_tmp_1049 = MUX_s_1_2_2((or_2604_nl), (or_2602_nl), inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6);
  assign or_2609_nl = (~ chn_inp_in_crt_sva_4_443_1) | (cfg_precision_1_sva_st_81!=2'b10);
  assign or_2610_nl = chn_inp_in_crt_sva_4_443_1 | (cfg_precision_1_sva_st_81!=2'b10);
  assign mux_1133_nl = MUX_s_1_2_2((or_2610_nl), (or_2609_nl), inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5);
  assign mux_1134_nl = MUX_s_1_2_2((mux_1133_nl), or_3379_cse, chn_inp_in_crt_sva_4_739_736_1[2]);
  assign nand_tmp_146 = ~(main_stage_v_4 & (~ (mux_1134_nl)));
  assign mux_tmp_1059 = MUX_s_1_2_2((~ inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5),
      inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5,
      inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5);
  assign nor_1131_nl = ~((~ main_stage_v_4) | (cfg_precision_1_sva_st_81!=2'b10)
      | (~((chn_inp_in_crt_sva_4_739_736_1[3]) | IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_3_tmp
      | FpAdd_6U_10U_1_is_a_greater_acc_3_itm_6_1 | inp_lookup_4_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp
      | mux_1140_cse)));
  assign or_2619_nl = nor_1130_cse | (chn_inp_in_crt_sva_5_739_736_1[3]) | IsNaN_8U_23U_3_land_lpi_1_dfm_5
      | IsNaN_6U_10U_8_land_lpi_1_dfm_4 | mux_tmp_1059;
  assign or_2621_nl = (chn_inp_in_crt_sva_5_739_736_1[3]) | IsNaN_8U_23U_3_land_lpi_1_dfm_5
      | IsNaN_6U_10U_8_land_lpi_1_dfm_4 | mux_tmp_1059;
  assign mux_1138_nl = MUX_s_1_2_2((or_2621_nl), (or_2619_nl), IsNaN_8U_23U_2_land_lpi_1_dfm_9);
  assign nor_1133_nl = ~((~ main_stage_v_5) | (cfg_precision_1_sva_st_82[0]) | (~((cfg_precision_1_sva_st_82[1])
      & (mux_1138_nl))));
  assign not_tmp_1080 = MUX_s_1_2_2((nor_1133_nl), (nor_1131_nl), or_11_cse);
  assign or_2640_nl = (~ inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5)
      | (~ main_stage_v_5) | (chn_inp_in_crt_sva_5_739_736_1[3]) | (cfg_precision_1_sva_st_82!=2'b10);
  assign or_2642_nl = inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
      | (~ main_stage_v_5) | (chn_inp_in_crt_sva_5_739_736_1[3]) | (cfg_precision_1_sva_st_82!=2'b10);
  assign mux_tmp_1067 = MUX_s_1_2_2((or_2642_nl), (or_2640_nl), inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5);
  assign or_tmp_2643 = (~ main_stage_v_5) | (chn_inp_in_crt_sva_5_739_736_1[3]) |
      (cfg_precision_1_sva_st_82!=2'b10);
  assign mux_1151_nl = MUX_s_1_2_2(or_2445_cse, or_2444_cse, chn_inp_in_crt_sva_4_459_1);
  assign mux_1152_nl = MUX_s_1_2_2((mux_1151_nl), or_3379_cse, chn_inp_in_crt_sva_4_739_736_1[3]);
  assign nand_tmp_148 = ~(main_stage_v_4 & (~ (mux_1152_nl)));
  assign or_tmp_2695 = IsNaN_6U_10U_9_land_lpi_1_dfm_7 | IsNaN_6U_10U_2_land_lpi_1_dfm_st_17;
  assign not_tmp_1108 = ~(or_tmp_2695 & main_stage_v_6);
  assign or_2698_nl = (cfg_precision_1_sva_st_83!=2'b10) | not_tmp_1108;
  assign mux_tmp_1092 = MUX_s_1_2_2((or_2698_nl), or_tmp_959, chn_inp_in_crt_sva_6_739_736_1[3]);
  assign or_2701_nl = (cfg_precision_1_sva_st_84!=2'b10) | (~(IsNaN_6U_10U_2_land_lpi_1_dfm_st_18
      & main_stage_v_7));
  assign or_2699_nl = (chn_inp_in_crt_sva_7_739_736_1[3]) | IsNaN_6U_10U_9_land_lpi_1_dfm_8;
  assign mux_1171_nl = MUX_s_1_2_2((or_2701_nl), or_tmp_1182, or_2699_nl);
  assign mux_1172_itm = MUX_s_1_2_2((mux_1171_nl), mux_tmp_1092, or_11_cse);
  assign or_tmp_2703 = IsNaN_6U_10U_9_land_3_lpi_1_dfm_7 | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_18;
  assign or_5684_itm = IsNaN_6U_10U_9_land_2_lpi_1_dfm_7 | (chn_inp_in_crt_sva_6_739_736_1[1])
      | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_18;
  assign or_tmp_2710 = (cfg_precision_1_sva_st_83[0]) | (~((cfg_precision_1_sva_st_83[1])
      & or_5684_itm & main_stage_v_6));
  assign mux_1176_nl = MUX_s_1_2_2(or_tmp_1147, or_tmp_2710, or_11_cse);
  assign and_3195_nl = main_stage_v_7 & IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_19;
  assign mux_1177_nl = MUX_s_1_2_2((and_3195_nl), main_stage_v_7, chn_inp_in_crt_sva_7_739_736_1[1]);
  assign or_2714_nl = (cfg_precision_1_sva_st_84[0]) | (~((cfg_precision_1_sva_st_84[1])
      & (mux_1177_nl)));
  assign mux_1178_nl = MUX_s_1_2_2((or_2714_nl), or_tmp_2710, or_11_cse);
  assign mux_1179_itm = MUX_s_1_2_2((mux_1178_nl), (mux_1176_nl), IsNaN_6U_10U_9_land_2_lpi_1_dfm_8);
  assign or_5683_itm = (chn_inp_in_crt_sva_6_739_736_1[0]) | IsNaN_6U_10U_9_land_1_lpi_1_dfm_7
      | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_18;
  assign or_tmp_2717 = (cfg_precision_1_sva_st_83!=2'b10) | (~(or_5683_itm & main_stage_v_6));
  assign mux_1180_nl = MUX_s_1_2_2(or_tmp_1182, or_tmp_2717, or_11_cse);
  assign mux_1181_nl = MUX_s_1_2_2(or_tmp_1058, or_tmp_2717, or_11_cse);
  assign mux_1182_itm = MUX_s_1_2_2((mux_1181_nl), (mux_1180_nl), FpAdd_6U_10U_1_or_12_cse);
  assign or_tmp_2723 = IsNaN_6U_10U_9_land_1_lpi_1_dfm_7 | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_18;
  assign or_tmp_2738 = IsNaN_6U_10U_9_land_2_lpi_1_dfm_7 | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_18;
  assign or_tmp_2768 = nor_1913_cse | (cfg_precision_1_sva_st_83!=2'b10) | (~ main_stage_v_6);
  assign or_tmp_2804 = (cfg_precision_1_sva_st_85[0]) | (~((cfg_precision_1_sva_st_85[1])
      & (chn_inp_in_crt_sva_8_739_736_1[1]) & IsNaN_6U_10U_land_2_lpi_1_dfm_5 & main_stage_v_8));
  assign and_3400_nl = main_stage_v_9 & (cfg_precision_1_sva_st_86==2'b10);
  assign nor_1058_nl = ~((~ main_stage_v_9) | (cfg_precision_1_sva_st_86!=2'b10));
  assign mux_1236_nl = MUX_s_1_2_2((nor_1058_nl), (and_3400_nl), inp_lookup_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_4);
  assign nand_tmp_162 = ~((chn_inp_in_crt_sva_9_739_736_1[0]) & (mux_1236_nl));
  assign and_3399_nl = main_stage_v_9 & (cfg_precision_1_sva_st_100==2'b10);
  assign nor_1056_nl = ~((~ main_stage_v_9) | (cfg_precision_1_sva_st_100!=2'b10));
  assign mux_1238_nl = MUX_s_1_2_2((nor_1056_nl), (and_3399_nl), inp_lookup_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_4);
  assign nand_tmp_163 = ~((chn_inp_in_crt_sva_9_739_736_1[1]) & (mux_1238_nl));
  assign and_3398_nl = main_stage_v_9 & (cfg_precision_1_sva_st_112==2'b10);
  assign nor_1054_nl = ~((~ main_stage_v_9) | (cfg_precision_1_sva_st_112!=2'b10));
  assign mux_1240_nl = MUX_s_1_2_2((nor_1054_nl), (and_3398_nl), inp_lookup_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_4);
  assign nand_tmp_164 = ~((chn_inp_in_crt_sva_9_739_736_1[2]) & (mux_1240_nl));
  assign and_3175_nl = main_stage_v_9 & (cfg_precision_1_sva_st_124==2'b10);
  assign nor_1052_nl = ~((~ main_stage_v_9) | (cfg_precision_1_sva_st_124!=2'b10));
  assign mux_1242_nl = MUX_s_1_2_2((nor_1052_nl), (and_3175_nl), inp_lookup_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_4);
  assign nand_tmp_165 = ~((chn_inp_in_crt_sva_9_739_736_1[3]) & (mux_1242_nl));
  assign or_tmp_2924 = (chn_inp_in_crt_sva_10_739_736_1[3]) | inp_lookup_else_unequal_tmp_36
      | (~ main_stage_v_10);
  assign or_tmp_2935 = (chn_inp_in_crt_sva_10_739_736_1[2]) | inp_lookup_else_unequal_tmp_36
      | (~ main_stage_v_10);
  assign not_tmp_1202 = ~((IsNaN_6U_10U_3_land_3_lpi_1_dfm_6 | IsNaN_6U_10U_2_land_3_lpi_1_dfm_24)
      & main_stage_v_10);
  assign or_tmp_2953 = (chn_inp_in_crt_sva_10_739_736_1[1]) | inp_lookup_else_unequal_tmp_36
      | (~ main_stage_v_10);
  assign not_tmp_1208 = ~((cfg_precision_1_sva_st_101[1]) & (IsNaN_6U_10U_3_land_2_lpi_1_dfm_6
      | IsNaN_6U_10U_2_land_2_lpi_1_dfm_24) & main_stage_v_10);
  assign or_tmp_2974 = (chn_inp_in_crt_sva_10_739_736_1[0]) | inp_lookup_else_unequal_tmp_36
      | (~ main_stage_v_10);
  assign not_tmp_1212 = ~((cfg_precision_1_sva_st_87[1]) & (IsNaN_6U_10U_3_land_1_lpi_1_dfm_6
      | IsNaN_6U_10U_2_land_1_lpi_1_dfm_24) & main_stage_v_10);
  assign and_tmp_181 = main_stage_v_10 & or_3291_cse;
  assign mux_tmp_1183 = MUX_s_1_2_2(main_stage_v_10, and_tmp_181, chn_inp_in_crt_sva_10_739_736_1[3]);
  assign and_tmp_182 = (chn_inp_in_crt_sva_10_739_736_1[3]) & mux_tmp_1183;
  assign or_tmp_2986 = (chn_inp_in_crt_sva_10_739_736_1[3]) | (~ main_stage_v_10);
  assign mux_tmp_1187 = MUX_s_1_2_2(main_stage_v_10, and_tmp_181, chn_inp_in_crt_sva_10_739_736_1[2]);
  assign and_tmp_184 = (chn_inp_in_crt_sva_10_739_736_1[2]) & mux_tmp_1187;
  assign or_tmp_2990 = (chn_inp_in_crt_sva_10_739_736_1[2]) | (~ main_stage_v_10);
  assign and_tmp_187 = (chn_inp_in_crt_sva_10_739_736_1[1]) & main_stage_v_10 & or_3291_cse;
  assign or_tmp_2993 = (chn_inp_in_crt_sva_10_739_736_1[1]) | (~ main_stage_v_10);
  assign mux_tmp_1195 = MUX_s_1_2_2(main_stage_v_10, and_tmp_181, chn_inp_in_crt_sva_10_739_736_1[0]);
  assign and_tmp_188 = (chn_inp_in_crt_sva_10_739_736_1[0]) & mux_tmp_1195;
  assign or_tmp_2997 = (chn_inp_in_crt_sva_10_739_736_1[0]) | (~ main_stage_v_10);
  assign or_tmp_2999 = (cfg_precision_1_sva_19!=2'b10) | (~ (chn_inp_in_crt_sva_9_739_736_1[0]))
      | IsNaN_6U_10U_2_land_1_lpi_1_dfm_23;
  assign or_tmp_3002 = (cfg_precision_1_sva_20!=2'b10) | (~ (chn_inp_in_crt_sva_10_739_736_1[0]))
      | IsNaN_6U_10U_2_land_1_lpi_1_dfm_24;
  assign or_tmp_3007 = (cfg_precision_1_sva_19!=2'b10) | (~ (chn_inp_in_crt_sva_9_739_736_1[0]));
  assign or_tmp_3011 = (cfg_precision_1_sva_20!=2'b10) | (~ (chn_inp_in_crt_sva_10_739_736_1[0]));
  assign and_3169_cse = or_3489_cse & main_stage_v_9;
  assign mux_tmp_1209 = MUX_s_1_2_2(and_3113_cse, and_3169_cse, chn_inp_in_crt_sva_9_739_736_1[0]);
  assign or_tmp_3017 = (cfg_precision_1_sva_19!=2'b10) | (~ (chn_inp_in_crt_sva_9_739_736_1[1]))
      | IsNaN_6U_10U_2_land_2_lpi_1_dfm_23;
  assign or_tmp_3020 = (cfg_precision_1_sva_20!=2'b10) | (~ (chn_inp_in_crt_sva_10_739_736_1[1]))
      | IsNaN_6U_10U_2_land_2_lpi_1_dfm_24;
  assign or_tmp_3025 = (cfg_precision_1_sva_19!=2'b10) | (~ (chn_inp_in_crt_sva_9_739_736_1[1]));
  assign or_tmp_3029 = (cfg_precision_1_sva_20!=2'b10) | (~ (chn_inp_in_crt_sva_10_739_736_1[1]));
  assign mux_tmp_1221 = MUX_s_1_2_2(and_3111_cse, and_3169_cse, chn_inp_in_crt_sva_9_739_736_1[1]);
  assign or_tmp_3035 = (cfg_precision_1_sva_19!=2'b10) | (~ (chn_inp_in_crt_sva_9_739_736_1[2]))
      | IsNaN_6U_10U_2_land_3_lpi_1_dfm_23;
  assign or_tmp_3038 = (cfg_precision_1_sva_20!=2'b10) | (~ (chn_inp_in_crt_sva_10_739_736_1[2]))
      | IsNaN_6U_10U_2_land_3_lpi_1_dfm_24;
  assign or_tmp_3043 = (cfg_precision_1_sva_19!=2'b10) | (~ (chn_inp_in_crt_sva_9_739_736_1[2]));
  assign or_tmp_3047 = (cfg_precision_1_sva_20!=2'b10) | (~ (chn_inp_in_crt_sva_10_739_736_1[2]));
  assign mux_tmp_1233 = MUX_s_1_2_2(and_3110_cse, and_3169_cse, chn_inp_in_crt_sva_9_739_736_1[2]);
  assign or_tmp_3053 = (cfg_precision_1_sva_19!=2'b10) | (~ (chn_inp_in_crt_sva_9_739_736_1[3]))
      | IsNaN_6U_10U_2_land_lpi_1_dfm_23;
  assign or_tmp_3056 = (cfg_precision_1_sva_20!=2'b10) | (~ (chn_inp_in_crt_sva_10_739_736_1[3]))
      | IsNaN_6U_10U_2_land_lpi_1_dfm_24;
  assign or_tmp_3061 = (cfg_precision_1_sva_19!=2'b10) | (~ (chn_inp_in_crt_sva_9_739_736_1[3]));
  assign or_tmp_3065 = (cfg_precision_1_sva_20!=2'b10) | (~ (chn_inp_in_crt_sva_10_739_736_1[3]));
  assign mux_tmp_1245 = MUX_s_1_2_2(and_3112_cse, and_3169_cse, chn_inp_in_crt_sva_9_739_736_1[3]);
  assign or_tmp_3087 = IsNaN_6U_10U_7_land_2_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_14;
  assign or_tmp_3123 = (chn_inp_in_crt_sva_3_739_736_1[1]) | (cfg_precision_1_sva_st_80!=2'b10)
      | IsNaN_6U_10U_6_land_2_lpi_1_dfm_5 | IsNaN_6U_10U_7_land_2_lpi_1_dfm_6 | nor_1371_cse;
  assign or_tmp_3132 = IsNaN_6U_10U_9_land_lpi_1_dfm_6 | IsNaN_6U_10U_8_land_lpi_1_dfm_4;
  assign or_3150_nl = (~((chn_inp_in_crt_sva_5_739_736_1[3]) | IsNaN_6U_10U_9_land_lpi_1_dfm_6
      | IsNaN_6U_10U_8_land_lpi_1_dfm_4)) | (cfg_precision_1_sva_st_82[0]) | not_tmp_374;
  assign mux_1347_itm = MUX_s_1_2_2(mux_tmp_1092, (or_3150_nl), or_11_cse);
  assign or_tmp_3152 = (~((chn_inp_in_crt_sva_5_739_736_1[2]) | IsNaN_6U_10U_9_land_3_lpi_1_dfm_6
      | IsNaN_6U_10U_8_land_3_lpi_1_dfm_4)) | (cfg_precision_1_sva_st_82!=2'b10)
      | (~ main_stage_v_5);
  assign or_tmp_3153 = IsNaN_6U_10U_9_land_3_lpi_1_dfm_6 | IsNaN_6U_10U_8_land_3_lpi_1_dfm_4;
  assign or_tmp_3156 = (chn_inp_in_crt_sva_5_739_736_1[2]) | (~(or_tmp_3153 & (cfg_precision_1_sva_st_82==2'b10)
      & main_stage_v_5));
  assign or_tmp_3160 = (chn_inp_in_crt_sva_6_739_736_1[2]) | (~(or_tmp_2703 & (cfg_precision_1_sva_st_83==2'b10)
      & main_stage_v_6));
  assign or_tmp_3180 = IsNaN_6U_10U_9_land_2_lpi_1_dfm_6 | IsNaN_6U_10U_8_land_2_lpi_1_dfm_4;
  assign or_3198_nl = (~((chn_inp_in_crt_sva_5_739_736_1[1]) | IsNaN_6U_10U_9_land_2_lpi_1_dfm_6
      | IsNaN_6U_10U_8_land_2_lpi_1_dfm_4)) | (cfg_precision_1_sva_st_82!=2'b10)
      | (~ main_stage_v_5);
  assign mux_1362_itm = MUX_s_1_2_2(or_tmp_2710, (or_3198_nl), or_11_cse);
  assign or_tmp_3200 = IsNaN_6U_10U_9_land_1_lpi_1_dfm_6 | IsNaN_6U_10U_8_land_1_lpi_1_dfm_6;
  assign or_3219_nl = (~((chn_inp_in_crt_sva_5_739_736_1[0]) | IsNaN_6U_10U_9_land_1_lpi_1_dfm_6
      | IsNaN_6U_10U_8_land_1_lpi_1_dfm_6)) | (cfg_precision_1_sva_st_82[0]) | not_tmp_374;
  assign mux_1367_itm = MUX_s_1_2_2(or_tmp_2717, (or_3219_nl), or_11_cse);
  assign or_tmp_3224 = (chn_inp_in_crt_sva_9_739_736_1[3]) | inp_lookup_else_unequal_tmp_35
      | (~ main_stage_v_9);
  assign or_tmp_3227 = (chn_inp_in_crt_sva_9_739_736_1[2]) | inp_lookup_else_unequal_tmp_35
      | (~ main_stage_v_9);
  assign or_tmp_3230 = (chn_inp_in_crt_sva_9_739_736_1[1]) | inp_lookup_else_unequal_tmp_35
      | (~ main_stage_v_9);
  assign or_tmp_3233 = (chn_inp_in_crt_sva_9_739_736_1[0]) | inp_lookup_else_unequal_tmp_35
      | (~ main_stage_v_9);
  assign or_tmp_3235 = (chn_inp_in_crt_sva_9_739_736_1[3]) | (~ main_stage_v_9);
  assign or_tmp_3246 = (chn_inp_in_crt_sva_9_739_736_1[2]) | (~ main_stage_v_9);
  assign or_tmp_3257 = (chn_inp_in_crt_sva_9_739_736_1[1]) | (~ main_stage_v_9);
  assign or_tmp_3268 = (chn_inp_in_crt_sva_9_739_736_1[0]) | (~ main_stage_v_9);
  assign not_tmp_1369 = ~(main_stage_v_9 & (chn_inp_in_crt_sva_9_739_736_1[0]));
  assign nor_tmp_464 = ((chn_inp_in_crt_sva_9_739_736_1!=4'b0000)) & main_stage_v_9;
  assign not_tmp_1373 = ~(main_stage_v_9 & (chn_inp_in_crt_sva_9_739_736_1[1]));
  assign not_tmp_1377 = ~(main_stage_v_9 & (chn_inp_in_crt_sva_9_739_736_1[2]));
  assign not_tmp_1381 = ~(main_stage_v_9 & (chn_inp_in_crt_sva_9_739_736_1[3]));
  assign or_3337_nl = (~ FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_7_0_1)
      | (cfg_precision_1_sva_st_91!=2'b10);
  assign or_3339_nl = FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_7_0_1
      | (cfg_precision_1_sva_st_91!=2'b10);
  assign mux_tmp_1367 = MUX_s_1_2_2((or_3339_nl), (or_3337_nl), FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_7_1_1);
  assign not_tmp_1388 = MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_7_0_1,
      (~ FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_7_0_1), FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_7_1_1);
  assign mux_1449_nl = MUX_s_1_2_2((~ FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_7_0_1),
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_7_0_1, FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_7_1_1);
  assign not_tmp_1391 = ~((cfg_precision_1_sva_st_91[1]) & (mux_1449_nl));
  assign not_tmp_1425 = ~((cfg_precision_1_sva_st_81[1]) & main_stage_v_4);
  assign and_3124_cse = main_stage_v_7 & (chn_inp_in_crt_sva_7_739_736_1[0]);
  assign or_3472_nl = (~ (chn_inp_in_crt_sva_7_739_736_1[0])) | (cfg_precision_1_sva_st_84!=2'b10);
  assign mux_tmp_1450 = MUX_s_1_2_2(main_stage_v_7, and_3124_cse, or_3472_nl);
  assign and_3122_nl = main_stage_v_7 & (chn_inp_in_crt_sva_7_739_736_1[1]);
  assign nor_500_nl = ~((cfg_precision_1_sva_st_84!=2'b10) | (~ (chn_inp_in_crt_sva_7_739_736_1[1])));
  assign mux_tmp_1452 = MUX_s_1_2_2((and_3122_nl), main_stage_v_7, nor_500_nl);
  assign and_3120_cse = main_stage_v_7 & (chn_inp_in_crt_sva_7_739_736_1[2]);
  assign or_3478_nl = (~ (chn_inp_in_crt_sva_7_739_736_1[2])) | (cfg_precision_1_sva_st_84!=2'b10);
  assign mux_tmp_1454 = MUX_s_1_2_2(main_stage_v_7, and_3120_cse, or_3478_nl);
  assign and_3118_cse = main_stage_v_7 & (chn_inp_in_crt_sva_7_739_736_1[3]);
  assign or_3480_nl = (~ (chn_inp_in_crt_sva_7_739_736_1[3])) | (cfg_precision_1_sva_st_84!=2'b10);
  assign mux_tmp_1458 = MUX_s_1_2_2(main_stage_v_7, and_3118_cse, or_3480_nl);
  assign or_tmp_3510 = (chn_inp_in_crt_sva_8_739_736_1[3]) | (~ main_stage_v_8);
  assign mux_1558_itm = MUX_s_1_2_2(or_tmp_3235, or_tmp_3510, or_11_cse);
  assign or_tmp_3512 = (chn_inp_in_crt_sva_8_739_736_1[2]) | (~ main_stage_v_8);
  assign mux_1559_itm = MUX_s_1_2_2(or_tmp_3246, or_tmp_3512, or_11_cse);
  assign or_tmp_3514 = (chn_inp_in_crt_sva_8_739_736_1[1]) | (~ main_stage_v_8);
  assign mux_1560_itm = MUX_s_1_2_2(or_tmp_3257, or_tmp_3514, or_11_cse);
  assign or_tmp_3516 = (chn_inp_in_crt_sva_8_739_736_1[0]) | (~ main_stage_v_8);
  assign mux_1561_itm = MUX_s_1_2_2(or_tmp_3268, or_tmp_3516, or_11_cse);
  assign mux_tmp_1485 = (chn_inp_in_crt_sva_8_739_736_1[3]) & main_stage_v_8 & or_3484_cse;
  assign mux_tmp_1488 = (chn_inp_in_crt_sva_8_739_736_1[2]) & main_stage_v_8 & or_3484_cse;
  assign mux_tmp_1494 = (chn_inp_in_crt_sva_8_739_736_1[0]) & main_stage_v_8 & or_3484_cse;
  assign nor_tmp_522 = ((chn_inp_in_crt_sva_8_739_736_1!=4'b0000)) & main_stage_v_8;
  assign or_tmp_3530 = (~ main_stage_v_7) | (chn_inp_in_crt_sva_7_739_736_1[0]) |
      (~ inp_lookup_else_unequal_tmp_33);
  assign or_tmp_3534 = (~ main_stage_v_7) | (chn_inp_in_crt_sva_7_739_736_1[1]) |
      (~ inp_lookup_else_unequal_tmp_33);
  assign or_tmp_3538 = (~ main_stage_v_7) | (chn_inp_in_crt_sva_7_739_736_1[2]) |
      (~ inp_lookup_else_unequal_tmp_33);
  assign or_tmp_3542 = (~ main_stage_v_7) | (chn_inp_in_crt_sva_7_739_736_1[3]) |
      (~ inp_lookup_else_unequal_tmp_33);
  assign nor_tmp_532 = (chn_inp_in_crt_sva_6_739_736_1[0]) & main_stage_v_6;
  assign nor_tmp_533 = (chn_inp_in_crt_sva_6_739_736_1[3]) & main_stage_v_6;
  assign nor_tmp_535 = (chn_inp_in_crt_sva_6_739_736_1[1]) & main_stage_v_6;
  assign and_3106_cse = (chn_inp_in_crt_sva_6_739_736_1[2]) & main_stage_v_6;
  assign mux_tmp_1509 = MUX_s_1_2_2(and_3106_cse, main_stage_v_6, chn_inp_in_crt_sva_6_739_736_1[2]);
  assign and_310_cse = main_stage_v_7 & or_3558_cse;
  assign mux_tmp_1511 = MUX_s_1_2_2(and_3118_cse, and_310_cse, chn_inp_in_crt_sva_7_739_736_1[3]);
  assign mux_tmp_1513 = MUX_s_1_2_2(and_3120_cse, and_310_cse, chn_inp_in_crt_sva_7_739_736_1[2]);
  assign mux_tmp_1518 = MUX_s_1_2_2(and_3124_cse, and_310_cse, chn_inp_in_crt_sva_7_739_736_1[0]);
  assign nor_tmp_545 = ((chn_inp_in_crt_sva_7_739_736_1!=4'b0000)) & main_stage_v_7;
  assign or_tmp_3562 = (~ main_stage_v_7) | (chn_inp_in_crt_sva_7_739_736_1[3]);
  assign or_tmp_3564 = (~ main_stage_v_7) | (chn_inp_in_crt_sva_7_739_736_1[2]);
  assign or_tmp_3566 = (~ main_stage_v_7) | (chn_inp_in_crt_sva_7_739_736_1[1]);
  assign or_tmp_3568 = (~ main_stage_v_7) | (chn_inp_in_crt_sva_7_739_736_1[0]);
  assign nor_tmp_551 = (chn_inp_in_crt_sva_5_739_736_1[0]) & main_stage_v_5;
  assign nor_tmp_552 = (chn_inp_in_crt_sva_5_739_736_1[1]) & main_stage_v_5;
  assign nor_tmp_553 = (chn_inp_in_crt_sva_5_739_736_1[2]) & main_stage_v_5;
  assign nor_tmp_555 = (chn_inp_in_crt_sva_5_739_736_1[3]) & main_stage_v_5;
  assign nand_326_cse = ~(inp_lookup_else_unequal_tmp_32 & main_stage_v_6);
  assign or_tmp_3612 = (chn_inp_in_crt_sva_6_739_736_1[3]) | nand_326_cse;
  assign or_tmp_3614 = (chn_inp_in_crt_sva_6_739_736_1[2]) | nand_326_cse;
  assign or_tmp_3616 = (chn_inp_in_crt_sva_6_739_736_1[1]) | nand_326_cse;
  assign or_tmp_3618 = (chn_inp_in_crt_sva_6_739_736_1[0]) | nand_326_cse;
  assign nor_tmp_560 = ((cfg_precision_1_sva_16!=2'b10)) & main_stage_v_6;
  assign mux_tmp_1543 = nor_tmp_560 & (chn_inp_in_crt_sva_6_739_736_1[3]);
  assign mux_tmp_1545 = MUX_s_1_2_2(and_3106_cse, nor_tmp_560, chn_inp_in_crt_sva_6_739_736_1[2]);
  assign mux_tmp_1548 = (chn_inp_in_crt_sva_6_739_736_1[1]) & nor_tmp_560;
  assign mux_tmp_1553 = (chn_inp_in_crt_sva_6_739_736_1[0]) & nor_tmp_560;
  assign nor_tmp_569 = ((chn_inp_in_crt_sva_6_739_736_1!=4'b0000)) & main_stage_v_6;
  assign or_tmp_3627 = (chn_inp_in_crt_sva_6_739_736_1[3]) | (~ main_stage_v_6);
  assign or_tmp_3629 = (chn_inp_in_crt_sva_6_739_736_1[2]) | (~ main_stage_v_6);
  assign or_tmp_3631 = (chn_inp_in_crt_sva_6_739_736_1[1]) | (~ main_stage_v_6);
  assign or_tmp_3633 = (chn_inp_in_crt_sva_6_739_736_1[0]) | (~ main_stage_v_6);
  assign and_tmp_225 = main_stage_v_4 & (chn_inp_in_crt_sva_4_739_736_1[0]);
  assign and_tmp_226 = main_stage_v_4 & (chn_inp_in_crt_sva_4_739_736_1[3]);
  assign and_tmp_227 = main_stage_v_4 & (chn_inp_in_crt_sva_4_739_736_1[1]);
  assign and_tmp_228 = main_stage_v_4 & (chn_inp_in_crt_sva_4_739_736_1[2]);
  assign not_tmp_1550 = ~(main_stage_v_5 & or_3384_cse);
  assign mux_tmp_1573 = MUX_s_1_2_2(not_tmp_1550, or_3716_cse, chn_inp_in_crt_sva_5_739_736_1[3]);
  assign mux_tmp_1575 = MUX_s_1_2_2(not_tmp_1550, or_3718_cse, chn_inp_in_crt_sva_5_739_736_1[2]);
  assign mux_tmp_1577 = MUX_s_1_2_2(not_tmp_1550, or_3720_cse, chn_inp_in_crt_sva_5_739_736_1[1]);
  assign mux_tmp_1579 = MUX_s_1_2_2(not_tmp_1550, or_3722_cse, chn_inp_in_crt_sva_5_739_736_1[0]);
  assign mux_tmp_1581 = main_stage_v_5 & or_3384_cse & (chn_inp_in_crt_sva_5_739_736_1[3]);
  assign mux_tmp_1583 = main_stage_v_5 & or_3384_cse & (chn_inp_in_crt_sva_5_739_736_1[2]);
  assign mux_tmp_1585 = main_stage_v_5 & or_3384_cse & (chn_inp_in_crt_sva_5_739_736_1[1]);
  assign mux_tmp_1587 = main_stage_v_5 & or_3384_cse & (chn_inp_in_crt_sva_5_739_736_1[0]);
  assign nand_tmp_218 = ~(main_stage_v_4 & (~((~ or_3379_cse) | (chn_inp_in_crt_sva_4_739_736_1[0]))));
  assign nand_tmp_219 = ~(main_stage_v_4 & (~((~ or_3379_cse) | (chn_inp_in_crt_sva_4_739_736_1[1]))));
  assign nand_tmp_220 = ~(main_stage_v_4 & (~((~ or_3379_cse) | (chn_inp_in_crt_sva_4_739_736_1[2]))));
  assign nand_tmp_221 = ~(main_stage_v_4 & (~((~ or_3379_cse) | (chn_inp_in_crt_sva_4_739_736_1[3]))));
  assign or_3781_nl = FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_4 | (~ inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5)
      | (cfg_precision_1_sva_st_81!=2'b10);
  assign mux_1694_nl = MUX_s_1_2_2((or_3781_nl), or_3379_cse, chn_inp_in_crt_sva_4_739_736_1[3]);
  assign nand_tmp_222 = ~(main_stage_v_4 & (~ (mux_1694_nl)));
  assign or_tmp_3798 = (~((~ inp_lookup_2_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp)
      | FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_1_itm_23_1)) | FpAdd_8U_23U_1_is_a_greater_acc_1_itm_8_1
      | IsNaN_6U_10U_5_land_2_lpi_1_dfm_5 | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10);
  assign or_tmp_3802 = (~((~((FpMul_6U_10U_1_p_mant_p1_2_sva[21]) | (~ inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4)
      | FpMul_6U_10U_1_lor_7_lpi_1_dfm_5)) | IsNaN_6U_10U_5_land_2_lpi_1_dfm_5))
      | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_15 | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10);
  assign or_tmp_3819 = (~((~ inp_lookup_3_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp)
      | FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_2_itm_23_1)) | FpAdd_8U_23U_1_is_a_greater_acc_2_itm_8_1
      | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10);
  assign or_tmp_3836 = (~((~((FpMul_6U_10U_1_p_mant_p1_sva[21]) | FpMul_6U_10U_1_lor_1_lpi_1_dfm_5
      | (~ inp_lookup_4_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs_2)))
      | IsNaN_6U_10U_5_land_lpi_1_dfm_5)) | IsNaN_6U_10U_2_land_lpi_1_dfm_st_15;
  assign and_tmp_240 = main_stage_v_4 & or_3379_cse & (chn_inp_in_crt_sva_4_739_736_1[3]);
  assign and_tmp_242 = main_stage_v_4 & or_3379_cse & (chn_inp_in_crt_sva_4_739_736_1[2]);
  assign and_tmp_244 = main_stage_v_4 & or_3379_cse & (chn_inp_in_crt_sva_4_739_736_1[1]);
  assign and_tmp_246 = main_stage_v_4 & or_3379_cse & (chn_inp_in_crt_sva_4_739_736_1[0]);
  assign or_tmp_3973 = FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_3 | (~ inp_lookup_3_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs)
      | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10);
  assign nand_tmp_230 = ~(main_stage_v_3 & (~((chn_inp_in_crt_sva_3_739_736_1[3])
      | (~ or_tmp_440))));
  assign nand_tmp_231 = ~(main_stage_v_3 & (~((~ or_tmp_440) | (chn_inp_in_crt_sva_3_739_736_1[2]))));
  assign nand_tmp_232 = ~(main_stage_v_3 & (~((~ or_tmp_440) | (chn_inp_in_crt_sva_3_739_736_1[1]))));
  assign nand_tmp_233 = ~(main_stage_v_3 & (~((~ or_tmp_440) | (chn_inp_in_crt_sva_3_739_736_1[0]))));
  assign or_3998_nl = (cfg_precision_1_sva_st_90!=2'b10) | IsNaN_8U_23U_2_land_1_lpi_1_dfm_st_6;
  assign mux_1821_nl = MUX_s_1_2_2(or_2010_cse, (or_3998_nl), chn_inp_in_crt_sva_1_739_395_1[341]);
  assign nand_tmp_234 = ~(main_stage_v_1 & (~ (mux_1821_nl)));
  assign or_4001_nl = (cfg_precision_1_sva_st_90!=2'b10) | IsNaN_8U_23U_2_land_2_lpi_1_dfm_st_6;
  assign mux_1825_nl = MUX_s_1_2_2(or_2010_cse, (or_4001_nl), chn_inp_in_crt_sva_1_739_395_1[342]);
  assign nand_tmp_235 = ~(main_stage_v_1 & (~ (mux_1825_nl)));
  assign nor_tmp_653 = ((~ nor_1336_cse_1) | (chn_inp_in_crt_sva_1_739_395_1[341]))
      & main_stage_v_1;
  assign nor_tmp_656 = ((~ nor_1340_cse) | (chn_inp_in_crt_sva_2_739_736_1[0])) &
      main_stage_v_2;
  assign nor_tmp_657 = ((~ nor_1336_cse_1) | (chn_inp_in_crt_sva_1_739_395_1[342]))
      & main_stage_v_1;
  assign nor_tmp_660 = ((~ nor_1340_cse) | (chn_inp_in_crt_sva_2_739_736_1[1])) &
      main_stage_v_2;
  assign nor_tmp_661 = (nor_758_cse | (chn_inp_in_crt_sva_1_739_395_1[343])) & main_stage_v_1;
  assign nor_tmp_664 = ((~ nor_1340_cse) | (chn_inp_in_crt_sva_2_739_736_1[2])) &
      main_stage_v_2;
  assign nor_tmp_665 = (nor_756_cse | (chn_inp_in_crt_sva_1_739_395_1[344])) & main_stage_v_1;
  assign nor_tmp_668 = ((~ nor_1340_cse) | (chn_inp_in_crt_sva_2_739_736_1[3])) &
      main_stage_v_2;
  assign and_dcpl_78 = (~ chn_inp_out_rsci_bawt) & reg_chn_inp_out_rsci_ld_core_psct_cse;
  assign or_dcpl_4 = and_dcpl_78 | (~ main_stage_v_12);
  assign and_dcpl_96 = or_11_cse & main_stage_v_12;
  assign and_dcpl_98 = (~ main_stage_v_12) & chn_inp_out_rsci_bawt & reg_chn_inp_out_rsci_ld_core_psct_cse;
  assign or_dcpl_8 = and_dcpl_78 | (~ main_stage_v_1);
  assign and_dcpl_105 = or_11_cse & (~ (chn_inp_in_rsci_d_mxwt[736]));
  assign and_dcpl_106 = inp_lookup_else_if_unequal_tmp_mx0w1 & or_11_cse;
  assign and_dcpl_107 = ~((chn_inp_in_rsci_d_mxwt[160]) | (chn_inp_in_rsci_d_mxwt[162]));
  assign and_dcpl_109 = ~((chn_inp_in_rsci_d_mxwt[159:158]!=2'b00));
  assign and_dcpl_132 = ~((chn_inp_in_rsci_d_mxwt[132:131]!=2'b00));
  assign and_dcpl_138 = (~((chn_inp_in_rsci_d_mxwt[148]) | (chn_inp_in_rsci_d_mxwt[161])
      | (chn_inp_in_rsci_d_mxwt[128]))) & (~((chn_inp_in_rsci_d_mxwt[130:129]!=2'b00)));
  assign and_dcpl_141 = ~((~ and_dcpl_138) | (~ and_dcpl_132) | (chn_inp_in_rsci_d_mxwt[133])
      | (chn_inp_in_rsci_d_mxwt[134]) | (chn_inp_in_rsci_d_mxwt[135]) | (chn_inp_in_rsci_d_mxwt[136])
      | (chn_inp_in_rsci_d_mxwt[137]) | (chn_inp_in_rsci_d_mxwt[138]) | (chn_inp_in_rsci_d_mxwt[139])
      | (chn_inp_in_rsci_d_mxwt[140]) | (chn_inp_in_rsci_d_mxwt[141]) | (chn_inp_in_rsci_d_mxwt[142])
      | (chn_inp_in_rsci_d_mxwt[143]) | (chn_inp_in_rsci_d_mxwt[144]) | (chn_inp_in_rsci_d_mxwt[145])
      | (chn_inp_in_rsci_d_mxwt[146]) | (chn_inp_in_rsci_d_mxwt[147]) | (chn_inp_in_rsci_d_mxwt[149])
      | (chn_inp_in_rsci_d_mxwt[150]) | (chn_inp_in_rsci_d_mxwt[151]) | (chn_inp_in_rsci_d_mxwt[152])
      | (chn_inp_in_rsci_d_mxwt[153]) | (chn_inp_in_rsci_d_mxwt[154]) | (chn_inp_in_rsci_d_mxwt[155])
      | (chn_inp_in_rsci_d_mxwt[156]) | (chn_inp_in_rsci_d_mxwt[157]) | (~ and_dcpl_109)
      | (~ and_dcpl_107) | (~ or_11_cse));
  assign and_dcpl_142 = (cfg_precision_rsci_d==2'b10);
  assign and_dcpl_144 = and_dcpl_142 & (~ (chn_inp_in_rsci_d_mxwt[736])) & or_11_cse;
  assign or_dcpl_44 = or_2_cse | (chn_inp_in_rsci_d_mxwt[736]);
  assign and_dcpl_145 = or_dcpl_44 & or_11_cse;
  assign and_dcpl_173 = ~((~ and_dcpl_138) | (~ and_dcpl_132) | (chn_inp_in_rsci_d_mxwt[133])
      | (chn_inp_in_rsci_d_mxwt[134]) | (chn_inp_in_rsci_d_mxwt[135]) | (chn_inp_in_rsci_d_mxwt[136])
      | (chn_inp_in_rsci_d_mxwt[137]) | (chn_inp_in_rsci_d_mxwt[138]) | (chn_inp_in_rsci_d_mxwt[139])
      | (chn_inp_in_rsci_d_mxwt[140]) | (chn_inp_in_rsci_d_mxwt[141]) | (chn_inp_in_rsci_d_mxwt[142])
      | (chn_inp_in_rsci_d_mxwt[143]) | (chn_inp_in_rsci_d_mxwt[144]) | (chn_inp_in_rsci_d_mxwt[145])
      | (chn_inp_in_rsci_d_mxwt[146]) | (chn_inp_in_rsci_d_mxwt[147]) | (chn_inp_in_rsci_d_mxwt[149])
      | (chn_inp_in_rsci_d_mxwt[150]) | (chn_inp_in_rsci_d_mxwt[151]) | (chn_inp_in_rsci_d_mxwt[152])
      | (chn_inp_in_rsci_d_mxwt[153]) | (chn_inp_in_rsci_d_mxwt[154]) | (chn_inp_in_rsci_d_mxwt[155])
      | (chn_inp_in_rsci_d_mxwt[156]) | (chn_inp_in_rsci_d_mxwt[157]) | (~ and_dcpl_109)
      | (~ and_dcpl_107));
  assign and_dcpl_176 = or_11_cse & (~ (chn_inp_in_rsci_d_mxwt[737]));
  assign and_dcpl_177 = inp_lookup_else_if_unequal_tmp_1_mx0w1 & or_11_cse;
  assign and_dcpl_178 = ~((chn_inp_in_rsci_d_mxwt[170]) | (chn_inp_in_rsci_d_mxwt[193]));
  assign and_dcpl_180 = ~((chn_inp_in_rsci_d_mxwt[192]) | (chn_inp_in_rsci_d_mxwt[194]));
  assign and_dcpl_203 = ~((chn_inp_in_rsci_d_mxwt[166:165]!=2'b00));
  assign and_dcpl_209 = (~((chn_inp_in_rsci_d_mxwt[197:195]!=3'b000))) & (~((chn_inp_in_rsci_d_mxwt[164:163]!=2'b00)));
  assign and_dcpl_212 = ~((~ and_dcpl_209) | (~ and_dcpl_203) | (chn_inp_in_rsci_d_mxwt[167])
      | (chn_inp_in_rsci_d_mxwt[168]) | (chn_inp_in_rsci_d_mxwt[169]) | (chn_inp_in_rsci_d_mxwt[171])
      | (chn_inp_in_rsci_d_mxwt[172]) | (chn_inp_in_rsci_d_mxwt[173]) | (chn_inp_in_rsci_d_mxwt[174])
      | (chn_inp_in_rsci_d_mxwt[175]) | (chn_inp_in_rsci_d_mxwt[176]) | (chn_inp_in_rsci_d_mxwt[177])
      | (chn_inp_in_rsci_d_mxwt[178]) | (chn_inp_in_rsci_d_mxwt[179]) | (chn_inp_in_rsci_d_mxwt[180])
      | (chn_inp_in_rsci_d_mxwt[181]) | (chn_inp_in_rsci_d_mxwt[182]) | (chn_inp_in_rsci_d_mxwt[183])
      | (chn_inp_in_rsci_d_mxwt[184]) | (chn_inp_in_rsci_d_mxwt[185]) | (chn_inp_in_rsci_d_mxwt[186])
      | (chn_inp_in_rsci_d_mxwt[187]) | (chn_inp_in_rsci_d_mxwt[188]) | (chn_inp_in_rsci_d_mxwt[189])
      | (chn_inp_in_rsci_d_mxwt[190]) | (chn_inp_in_rsci_d_mxwt[191]) | (~ and_dcpl_180)
      | (~ and_dcpl_178) | (~ or_11_cse));
  assign and_dcpl_214 = and_dcpl_142 & (~ (chn_inp_in_rsci_d_mxwt[737])) & or_11_cse;
  assign or_dcpl_80 = or_2_cse | (chn_inp_in_rsci_d_mxwt[737]);
  assign and_dcpl_215 = or_dcpl_80 & or_11_cse;
  assign and_dcpl_243 = ~((~ and_dcpl_209) | (~ and_dcpl_203) | (chn_inp_in_rsci_d_mxwt[167])
      | (chn_inp_in_rsci_d_mxwt[168]) | (chn_inp_in_rsci_d_mxwt[169]) | (chn_inp_in_rsci_d_mxwt[171])
      | (chn_inp_in_rsci_d_mxwt[172]) | (chn_inp_in_rsci_d_mxwt[173]) | (chn_inp_in_rsci_d_mxwt[174])
      | (chn_inp_in_rsci_d_mxwt[175]) | (chn_inp_in_rsci_d_mxwt[176]) | (chn_inp_in_rsci_d_mxwt[177])
      | (chn_inp_in_rsci_d_mxwt[178]) | (chn_inp_in_rsci_d_mxwt[179]) | (chn_inp_in_rsci_d_mxwt[180])
      | (chn_inp_in_rsci_d_mxwt[181]) | (chn_inp_in_rsci_d_mxwt[182]) | (chn_inp_in_rsci_d_mxwt[183])
      | (chn_inp_in_rsci_d_mxwt[184]) | (chn_inp_in_rsci_d_mxwt[185]) | (chn_inp_in_rsci_d_mxwt[186])
      | (chn_inp_in_rsci_d_mxwt[187]) | (chn_inp_in_rsci_d_mxwt[188]) | (chn_inp_in_rsci_d_mxwt[189])
      | (chn_inp_in_rsci_d_mxwt[190]) | (chn_inp_in_rsci_d_mxwt[191]) | (~ and_dcpl_180)
      | (~ and_dcpl_178));
  assign and_dcpl_246 = or_11_cse & (~ (chn_inp_in_rsci_d_mxwt[738]));
  assign and_dcpl_247 = or_79_cse & or_11_cse;
  assign and_dcpl_248 = ~((chn_inp_in_rsci_d_mxwt[199:198]!=2'b00));
  assign and_dcpl_250 = ~((chn_inp_in_rsci_d_mxwt[232]) | (chn_inp_in_rsci_d_mxwt[202]));
  assign and_dcpl_273 = ~((chn_inp_in_rsci_d_mxwt[207:206]!=2'b00));
  assign and_dcpl_279 = (~((chn_inp_in_rsci_d_mxwt[200]) | (chn_inp_in_rsci_d_mxwt[201])
      | (chn_inp_in_rsci_d_mxwt[203]))) & (~((chn_inp_in_rsci_d_mxwt[205:204]!=2'b00)));
  assign and_dcpl_282 = ~((~ and_dcpl_279) | (~ and_dcpl_273) | (chn_inp_in_rsci_d_mxwt[231:208]!=24'b000000000000000000000000)
      | (~ and_dcpl_250) | (~ and_dcpl_248) | (~ or_11_cse));
  assign and_dcpl_284 = and_dcpl_142 & (~ (chn_inp_in_rsci_d_mxwt[738])) & or_11_cse;
  assign or_dcpl_116 = or_2_cse | (chn_inp_in_rsci_d_mxwt[738]);
  assign and_dcpl_285 = or_dcpl_116 & or_11_cse;
  assign and_dcpl_313 = ~((~ and_dcpl_279) | (~ and_dcpl_273) | (chn_inp_in_rsci_d_mxwt[231:208]!=24'b000000000000000000000000)
      | (~ and_dcpl_250) | (~ and_dcpl_248));
  assign and_dcpl_316 = or_11_cse & (~ (chn_inp_in_rsci_d_mxwt[739]));
  assign and_dcpl_317 = inp_lookup_else_if_unequal_tmp_3_mx0w1 & or_11_cse;
  assign and_dcpl_318 = ~((chn_inp_in_rsci_d_mxwt[267:266]!=2'b00));
  assign and_dcpl_320 = ~((chn_inp_in_rsci_d_mxwt[265:264]!=2'b00));
  assign and_dcpl_343 = ~((chn_inp_in_rsci_d_mxwt[235:234]!=2'b00));
  assign and_dcpl_349 = (~((chn_inp_in_rsci_d_mxwt[244]) | (chn_inp_in_rsci_d_mxwt[238])
      | (chn_inp_in_rsci_d_mxwt[237]))) & (~((chn_inp_in_rsci_d_mxwt[239]) | (chn_inp_in_rsci_d_mxwt[233])));
  assign and_dcpl_352 = ~((~ and_dcpl_349) | (~ and_dcpl_343) | (chn_inp_in_rsci_d_mxwt[236])
      | (chn_inp_in_rsci_d_mxwt[240]) | (chn_inp_in_rsci_d_mxwt[241]) | (chn_inp_in_rsci_d_mxwt[242])
      | (chn_inp_in_rsci_d_mxwt[243]) | (chn_inp_in_rsci_d_mxwt[245]) | (chn_inp_in_rsci_d_mxwt[246])
      | (chn_inp_in_rsci_d_mxwt[247]) | (chn_inp_in_rsci_d_mxwt[248]) | (chn_inp_in_rsci_d_mxwt[249])
      | (chn_inp_in_rsci_d_mxwt[250]) | (chn_inp_in_rsci_d_mxwt[251]) | (chn_inp_in_rsci_d_mxwt[252])
      | (chn_inp_in_rsci_d_mxwt[253]) | (chn_inp_in_rsci_d_mxwt[254]) | (chn_inp_in_rsci_d_mxwt[255])
      | (chn_inp_in_rsci_d_mxwt[256]) | (chn_inp_in_rsci_d_mxwt[257]) | (chn_inp_in_rsci_d_mxwt[258])
      | (chn_inp_in_rsci_d_mxwt[259]) | (chn_inp_in_rsci_d_mxwt[260]) | (chn_inp_in_rsci_d_mxwt[261])
      | (chn_inp_in_rsci_d_mxwt[262]) | (chn_inp_in_rsci_d_mxwt[263]) | (~ and_dcpl_320)
      | (~ and_dcpl_318) | (~ or_11_cse));
  assign and_dcpl_354 = and_dcpl_142 & (~ (chn_inp_in_rsci_d_mxwt[739])) & or_11_cse;
  assign or_dcpl_152 = or_2_cse | (chn_inp_in_rsci_d_mxwt[739]);
  assign and_dcpl_355 = or_dcpl_152 & or_11_cse;
  assign and_dcpl_383 = ~((~ and_dcpl_349) | (~ and_dcpl_343) | (chn_inp_in_rsci_d_mxwt[236])
      | (chn_inp_in_rsci_d_mxwt[240]) | (chn_inp_in_rsci_d_mxwt[241]) | (chn_inp_in_rsci_d_mxwt[242])
      | (chn_inp_in_rsci_d_mxwt[243]) | (chn_inp_in_rsci_d_mxwt[245]) | (chn_inp_in_rsci_d_mxwt[246])
      | (chn_inp_in_rsci_d_mxwt[247]) | (chn_inp_in_rsci_d_mxwt[248]) | (chn_inp_in_rsci_d_mxwt[249])
      | (chn_inp_in_rsci_d_mxwt[250]) | (chn_inp_in_rsci_d_mxwt[251]) | (chn_inp_in_rsci_d_mxwt[252])
      | (chn_inp_in_rsci_d_mxwt[253]) | (chn_inp_in_rsci_d_mxwt[254]) | (chn_inp_in_rsci_d_mxwt[255])
      | (chn_inp_in_rsci_d_mxwt[256]) | (chn_inp_in_rsci_d_mxwt[257]) | (chn_inp_in_rsci_d_mxwt[258])
      | (chn_inp_in_rsci_d_mxwt[259]) | (chn_inp_in_rsci_d_mxwt[260]) | (chn_inp_in_rsci_d_mxwt[261])
      | (chn_inp_in_rsci_d_mxwt[262]) | (chn_inp_in_rsci_d_mxwt[263]) | (~ and_dcpl_320)
      | (~ and_dcpl_318));
  assign and_dcpl_390 = or_11_cse & (~ FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_5);
  assign and_dcpl_393 = or_11_cse & (~ (chn_inp_in_crt_sva_1_739_395_1[341]));
  assign and_dcpl_394 = or_11_cse & (chn_inp_in_crt_sva_1_739_395_1[341]);
  assign and_dcpl_398 = or_11_cse & (~ FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_5);
  assign and_dcpl_401 = or_11_cse & (~ (chn_inp_in_crt_sva_1_739_395_1[342]));
  assign and_dcpl_402 = or_11_cse & (chn_inp_in_crt_sva_1_739_395_1[342]);
  assign and_dcpl_406 = or_11_cse & (~ FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_5);
  assign and_dcpl_409 = or_11_cse & (~ (chn_inp_in_crt_sva_1_739_395_1[343]));
  assign and_dcpl_410 = or_11_cse & (chn_inp_in_crt_sva_1_739_395_1[343]);
  assign and_dcpl_412 = or_11_cse & (~ FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2);
  assign and_dcpl_415 = or_11_cse & (~ (chn_inp_in_crt_sva_1_739_395_1[344]));
  assign and_dcpl_416 = or_11_cse & (chn_inp_in_crt_sva_1_739_395_1[344]);
  assign and_dcpl_419 = or_11_cse & main_stage_v_2;
  assign and_dcpl_423 = (cfg_precision_1_sva_st_91==2'b10);
  assign and_dcpl_427 = or_11_cse & (chn_inp_in_crt_sva_2_739_736_1[0]);
  assign and_dcpl_428 = ~((chn_inp_in_crt_sva_2_739_736_1[0]) | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_14);
  assign and_dcpl_433 = (~ (chn_inp_in_crt_sva_2_739_736_1[0])) & IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_14;
  assign and_dcpl_437 = and_dcpl_423 & (chn_inp_in_crt_sva_2_739_736_1[0]) & main_stage_v_2;
  assign and_dcpl_453 = and_dcpl_423 & (~ (chn_inp_in_crt_sva_2_739_736_1[0])) &
      and_dcpl_419;
  assign and_dcpl_454 = ~((cfg_precision_1_sva_st_80[0]) | (chn_inp_in_crt_sva_3_739_736_1[0]));
  assign or_dcpl_159 = or_tmp_439 | (chn_inp_in_crt_sva_2_739_736_1[0]) | (~ main_stage_v_2);
  assign and_dcpl_458 = or_dcpl_159 & (cfg_precision_1_sva_st_80[1]) & and_dcpl_454
      & main_stage_v_3 & or_11_cse;
  assign and_dcpl_459 = or_11_cse & (~ (chn_inp_in_crt_sva_2_739_736_1[0]));
  assign and_dcpl_464 = or_11_cse & (chn_inp_in_crt_sva_2_739_736_1[1]);
  assign and_dcpl_465 = ~(IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_14 | IsNaN_6U_10U_7_land_2_lpi_1_dfm_5);
  assign and_dcpl_468 = (~ IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_14) & IsNaN_6U_10U_7_land_2_lpi_1_dfm_5;
  assign and_dcpl_471 = IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_14 & (~ (chn_inp_in_crt_sva_2_739_736_1[1]));
  assign and_dcpl_488 = or_11_cse & (~ (chn_inp_in_crt_sva_2_739_736_1[1]));
  assign or_dcpl_163 = or_tmp_439 | (chn_inp_in_crt_sva_2_739_736_1[1]) | (~ main_stage_v_2);
  assign and_dcpl_495 = or_dcpl_163 & (cfg_precision_1_sva_st_80==2'b10) & (~ (chn_inp_in_crt_sva_3_739_736_1[1]))
      & main_stage_v_3 & or_11_cse;
  assign and_dcpl_496 = or_11_cse & (chn_inp_in_crt_sva_2_739_736_1[2]);
  assign and_dcpl_498 = and_dcpl_423 & main_stage_v_2;
  assign and_dcpl_504 = (~ IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_14) & IsNaN_6U_10U_7_land_3_lpi_1_dfm_5;
  assign and_dcpl_524 = or_11_cse & (~ (chn_inp_in_crt_sva_2_739_736_1[2]));
  assign and_dcpl_526 = (cfg_precision_1_sva_st_80[1]) & (~ (chn_inp_in_crt_sva_3_739_736_1[2]));
  assign or_dcpl_167 = or_tmp_439 | (~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[2]);
  assign and_dcpl_530 = or_dcpl_167 & (~ (cfg_precision_1_sva_st_80[0])) & and_dcpl_526
      & main_stage_v_3 & or_11_cse;
  assign and_dcpl_535 = or_11_cse & (chn_inp_in_crt_sva_2_739_736_1[3]);
  assign and_dcpl_539 = (~ IsNaN_6U_10U_2_land_lpi_1_dfm_st_14) & IsNaN_6U_10U_7_land_lpi_1_dfm_5;
  assign and_dcpl_559 = or_11_cse & (~ (chn_inp_in_crt_sva_2_739_736_1[3]));
  assign and_dcpl_560 = or_11_cse & main_stage_v_3;
  assign and_dcpl_564 = or_11_cse & (chn_inp_in_crt_sva_3_739_736_1[0]);
  assign and_dcpl_565 = or_11_cse & (~ (chn_inp_in_crt_sva_3_739_736_1[0]));
  assign and_dcpl_567 = (cfg_precision_1_sva_st_80==2'b10) & (~ (chn_inp_in_crt_sva_3_739_736_1[0]));
  assign and_dcpl_573 = (or_tmp_440 | (chn_inp_in_crt_sva_3_739_736_1[0]) | (~ main_stage_v_3))
      & (cfg_precision_1_sva_st_81==2'b10) & (~ (chn_inp_in_crt_sva_4_739_736_1[0]))
      & main_stage_v_4 & or_11_cse;
  assign and_dcpl_575 = (or_tmp_440 | (chn_inp_in_crt_sva_3_739_736_1[0])) & or_11_cse;
  assign and_dcpl_582 = or_11_cse & (chn_inp_in_crt_sva_3_739_736_1[1]);
  assign and_dcpl_583 = or_11_cse & (~ (chn_inp_in_crt_sva_3_739_736_1[1]));
  assign and_dcpl_584 = (cfg_precision_1_sva_st_80==2'b10);
  assign and_dcpl_585 = and_dcpl_584 & (~ (chn_inp_in_crt_sva_3_739_736_1[1]));
  assign and_dcpl_591 = (or_tmp_440 | (chn_inp_in_crt_sva_3_739_736_1[1]) | (~ main_stage_v_3))
      & (cfg_precision_1_sva_st_81==2'b10) & (~ (chn_inp_in_crt_sva_4_739_736_1[1]))
      & main_stage_v_4 & or_11_cse;
  assign and_dcpl_593 = (or_tmp_440 | (chn_inp_in_crt_sva_3_739_736_1[1])) & or_11_cse;
  assign and_dcpl_597 = ~(IsNaN_6U_10U_5_land_2_lpi_1_dfm_5 | (chn_inp_in_crt_sva_3_739_736_1[1]));
  assign and_dcpl_600 = or_11_cse & (chn_inp_in_crt_sva_3_739_736_1[2]);
  assign and_dcpl_601 = or_11_cse & (~ (chn_inp_in_crt_sva_3_739_736_1[2]));
  assign and_dcpl_603 = and_dcpl_584 & (~ (chn_inp_in_crt_sva_3_739_736_1[2]));
  assign and_dcpl_609 = (or_tmp_440 | (chn_inp_in_crt_sva_3_739_736_1[2]) | (~ main_stage_v_3))
      & (cfg_precision_1_sva_st_81==2'b10) & (~ (chn_inp_in_crt_sva_4_739_736_1[2]))
      & main_stage_v_4 & or_11_cse;
  assign and_dcpl_611 = (or_tmp_440 | (chn_inp_in_crt_sva_3_739_736_1[2])) & or_11_cse;
  assign and_dcpl_613 = (~ (chn_inp_in_crt_sva_3_739_736_1[2])) & main_stage_v_3
      & or_11_cse;
  assign and_dcpl_615 = ~(IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_15 | (cfg_precision_1_sva_st_80[0]));
  assign and_dcpl_627 = ~(IsNaN_6U_10U_5_land_3_lpi_1_dfm_5 | (chn_inp_in_crt_sva_3_739_736_1[2]));
  assign and_dcpl_630 = or_11_cse & (chn_inp_in_crt_sva_3_739_736_1[3]);
  assign and_dcpl_631 = or_11_cse & (~ (chn_inp_in_crt_sva_3_739_736_1[3]));
  assign and_dcpl_633 = and_dcpl_584 & (~ (chn_inp_in_crt_sva_3_739_736_1[3]));
  assign or_dcpl_186 = or_tmp_440 | (chn_inp_in_crt_sva_3_739_736_1[3]) | (~ main_stage_v_3);
  assign and_dcpl_639 = or_dcpl_186 & (cfg_precision_1_sva_st_81==2'b10) & (~ (chn_inp_in_crt_sva_4_739_736_1[3]))
      & main_stage_v_4 & or_11_cse;
  assign or_tmp_4220 = (chn_inp_in_crt_sva_3_739_736_1[3]) | (cfg_precision_1_sva_st_80!=2'b10);
  assign and_dcpl_641 = or_tmp_4220 & or_11_cse;
  assign and_dcpl_642 = (~ (chn_inp_in_crt_sva_3_739_736_1[3])) & IsNaN_6U_10U_5_land_lpi_1_dfm_5;
  assign and_dcpl_645 = ~((chn_inp_in_crt_sva_3_739_736_1[3]) | IsNaN_6U_10U_5_land_lpi_1_dfm_5);
  assign and_dcpl_654 = or_11_cse & (chn_inp_in_crt_sva_4_739_736_1[0]);
  assign and_dcpl_655 = or_11_cse & (~ (chn_inp_in_crt_sva_4_739_736_1[0]));
  assign and_dcpl_662 = or_11_cse & (chn_inp_in_crt_sva_4_739_736_1[1]);
  assign and_dcpl_663 = or_11_cse & (~ (chn_inp_in_crt_sva_4_739_736_1[1]));
  assign and_dcpl_670 = or_11_cse & (chn_inp_in_crt_sva_4_739_736_1[2]);
  assign and_dcpl_671 = or_11_cse & (~ (chn_inp_in_crt_sva_4_739_736_1[2]));
  assign mux_tmp_1821 = MUX_s_1_2_2((chn_inp_in_crt_sva_5_739_736_1[2]), (chn_inp_in_crt_sva_4_739_736_1[2]),
      or_11_cse);
  assign and_dcpl_678 = or_11_cse & (chn_inp_in_crt_sva_4_739_736_1[3]);
  assign and_dcpl_679 = or_11_cse & (~ (chn_inp_in_crt_sva_4_739_736_1[3]));
  assign and_dcpl_688 = or_11_cse & (~ IsNaN_8U_23U_3_land_1_lpi_1_dfm_6);
  assign and_dcpl_690 = or_11_cse & (chn_inp_in_crt_sva_5_739_736_1[0]);
  assign and_dcpl_691 = or_11_cse & (~ (chn_inp_in_crt_sva_5_739_736_1[0]));
  assign and_dcpl_699 = or_11_cse & (~ IsNaN_8U_23U_3_land_2_lpi_1_dfm_6);
  assign and_dcpl_701 = or_11_cse & (chn_inp_in_crt_sva_5_739_736_1[1]);
  assign and_dcpl_702 = or_11_cse & (~ (chn_inp_in_crt_sva_5_739_736_1[1]));
  assign and_dcpl_712 = or_11_cse & (chn_inp_in_crt_sva_5_739_736_1[2]);
  assign and_dcpl_713 = or_11_cse & (~ (chn_inp_in_crt_sva_5_739_736_1[2]));
  assign nor_tmp_686 = IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_4 & (chn_inp_in_crt_sva_6_739_736_1[2]);
  assign and_dcpl_717 = or_11_cse & (~ IsNaN_8U_23U_3_land_lpi_1_dfm_5);
  assign and_dcpl_719 = or_11_cse & (chn_inp_in_crt_sva_5_739_736_1[3]);
  assign and_dcpl_720 = or_11_cse & (~ (chn_inp_in_crt_sva_5_739_736_1[3]));
  assign and_dcpl_740 = or_11_cse & (~ (chn_inp_in_crt_sva_6_739_736_1[0]));
  assign and_dcpl_741 = or_11_cse & (chn_inp_in_crt_sva_6_739_736_1[0]);
  assign and_dcpl_752 = or_11_cse & (~ (chn_inp_in_crt_sva_6_739_736_1[1]));
  assign and_dcpl_753 = or_11_cse & (chn_inp_in_crt_sva_6_739_736_1[1]);
  assign and_dcpl_764 = or_11_cse & (~ (chn_inp_in_crt_sva_6_739_736_1[2]));
  assign and_dcpl_765 = or_11_cse & (chn_inp_in_crt_sva_6_739_736_1[2]);
  assign and_dcpl_776 = or_11_cse & (~ (chn_inp_in_crt_sva_6_739_736_1[3]));
  assign and_dcpl_777 = or_11_cse & (chn_inp_in_crt_sva_6_739_736_1[3]);
  assign and_dcpl_784 = or_11_cse & (chn_inp_in_crt_sva_7_739_736_1[0]);
  assign and_dcpl_785 = or_11_cse & (~ (chn_inp_in_crt_sva_7_739_736_1[0]));
  assign and_dcpl_787 = IsNaN_6U_10U_IsNaN_6U_10U_nor_tmp & (chn_inp_in_crt_sva_7_739_736_1[0])
      & or_11_cse;
  assign and_dcpl_798 = (~ IsNaN_6U_10U_IsNaN_6U_10U_nor_tmp) & (chn_inp_in_crt_sva_7_739_736_1[0])
      & or_11_cse;
  assign and_dcpl_801 = ~((chn_inp_in_crt_sva_7_739_736_1[0]) | IsNaN_6U_10U_8_land_1_lpi_1_dfm_7
      | IsNaN_6U_10U_9_land_1_lpi_1_dfm_8);
  assign and_dcpl_807 = or_11_cse & (chn_inp_in_crt_sva_7_739_736_1[1]);
  assign and_dcpl_808 = or_11_cse & (~ (chn_inp_in_crt_sva_7_739_736_1[1]));
  assign and_dcpl_810 = (chn_inp_in_crt_sva_7_739_736_1[1]) & IsNaN_6U_10U_IsNaN_6U_10U_nor_1_tmp
      & or_11_cse;
  assign and_dcpl_821 = (chn_inp_in_crt_sva_7_739_736_1[1]) & (~ IsNaN_6U_10U_IsNaN_6U_10U_nor_1_tmp)
      & or_11_cse;
  assign and_dcpl_825 = or_11_cse & (~ IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_19);
  assign and_dcpl_831 = or_11_cse & (chn_inp_in_crt_sva_7_739_736_1[2]);
  assign and_dcpl_832 = or_11_cse & (~ (chn_inp_in_crt_sva_7_739_736_1[2]));
  assign and_dcpl_834 = (chn_inp_in_crt_sva_7_739_736_1[2]) & IsNaN_6U_10U_IsNaN_6U_10U_nor_2_tmp
      & or_11_cse;
  assign and_dcpl_845 = (chn_inp_in_crt_sva_7_739_736_1[2]) & (~ IsNaN_6U_10U_IsNaN_6U_10U_nor_2_tmp)
      & or_11_cse;
  assign and_dcpl_847 = or_11_cse & (~ IsNaN_6U_10U_9_land_3_lpi_1_dfm_8);
  assign and_dcpl_856 = or_11_cse & (chn_inp_in_crt_sva_7_739_736_1[3]);
  assign and_dcpl_857 = or_11_cse & (~ (chn_inp_in_crt_sva_7_739_736_1[3]));
  assign and_dcpl_859 = (chn_inp_in_crt_sva_7_739_736_1[3]) & IsNaN_6U_10U_IsNaN_6U_10U_nor_3_tmp
      & or_11_cse;
  assign and_dcpl_870 = (chn_inp_in_crt_sva_7_739_736_1[3]) & (~ IsNaN_6U_10U_IsNaN_6U_10U_nor_3_tmp)
      & or_11_cse;
  assign and_dcpl_872 = ~(IsNaN_6U_10U_9_land_lpi_1_dfm_8 | (chn_inp_in_crt_sva_7_739_736_1[3]));
  assign and_dcpl_874 = or_11_cse & (~ IsNaN_6U_10U_2_land_lpi_1_dfm_st_18);
  assign or_dcpl_257 = (cfg_precision_1_sva_st_125!=2'b10);
  assign or_dcpl_264 = (cfg_precision_1_sva_st_89!=2'b10);
  assign or_dcpl_267 = or_dcpl_264 | (~ (chn_inp_in_crt_sva_12_739_736_1[0]));
  assign or_dcpl_269 = (cfg_precision_1_sva_st_103!=2'b10) | (~ (chn_inp_in_crt_sva_12_739_736_1[1]));
  assign or_dcpl_276 = (~ (chn_inp_in_crt_sva_12_739_736_1[2])) | (cfg_precision_1_sva_st_115!=2'b10);
  assign or_dcpl_278 = (cfg_precision_1_sva_st_127!=2'b10) | (~ (chn_inp_in_crt_sva_12_739_736_1[3]));
  assign and_dcpl_927 = (cfg_precision_1_sva_st_87==2'b10);
  assign nor_689_nl = ~(FpAdd_6U_10U_is_a_greater_oif_aelse_acc_itm_10_1 | (~ inp_lookup_1_FpAdd_6U_10U_is_a_greater_oif_equal_tmp));
  assign mux_tmp_1835 = MUX_s_1_2_2((nor_689_nl), inp_lookup_1_FpAdd_6U_10U_is_a_greater_oif_equal_svs,
      reg_inp_lookup_1_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse);
  assign or_dcpl_280 = mux_tmp_1835 | reg_inp_lookup_1_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse;
  assign and_dcpl_930 = or_dcpl_280 & and_dcpl_927 & (chn_inp_in_crt_sva_10_739_736_1[0])
      & or_11_cse;
  assign and_dcpl_935 = (~ mux_tmp_1835) & (cfg_precision_1_sva_st_87==2'b10) & (~
      reg_inp_lookup_1_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse) & (chn_inp_in_crt_sva_10_739_736_1[0])
      & or_11_cse;
  assign and_dcpl_936 = ((cfg_precision_1_sva_st_87!=2'b10) | (~ (chn_inp_in_crt_sva_10_739_736_1[0])))
      & or_11_cse;
  assign and_dcpl_937 = (cfg_precision_1_sva_st_101==2'b10);
  assign nor_691_nl = ~((~ inp_lookup_2_FpAdd_6U_10U_is_a_greater_oif_equal_tmp)
      | FpAdd_6U_10U_is_a_greater_oif_aelse_acc_1_itm_10_1);
  assign mux_tmp_1836 = MUX_s_1_2_2((nor_691_nl), inp_lookup_2_FpAdd_6U_10U_is_a_greater_oif_equal_svs,
      reg_inp_lookup_2_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse);
  assign or_dcpl_283 = mux_tmp_1836 | reg_inp_lookup_2_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse;
  assign and_dcpl_940 = or_dcpl_283 & and_dcpl_937 & (chn_inp_in_crt_sva_10_739_736_1[1])
      & or_11_cse;
  assign and_dcpl_941 = (chn_inp_in_crt_sva_10_739_736_1[1]) & (~ reg_inp_lookup_2_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse);
  assign and_dcpl_943 = (~ mux_tmp_1836) & or_11_cse;
  assign and_dcpl_944 = and_dcpl_943 & and_dcpl_937 & and_dcpl_941;
  assign and_dcpl_945 = ((cfg_precision_1_sva_st_101!=2'b10) | (~ (chn_inp_in_crt_sva_10_739_736_1[1])))
      & or_11_cse;
  assign and_dcpl_947 = (cfg_precision_1_sva_st_113==2'b10) & (chn_inp_in_crt_sva_10_739_736_1[2]);
  assign nand_241_nl = ~(reg_inp_lookup_3_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse
      & (~ inp_lookup_3_FpAdd_6U_10U_is_a_greater_oif_equal_svs));
  assign and_3053_nl = reg_inp_lookup_3_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse
      & inp_lookup_3_FpAdd_6U_10U_is_a_greater_oif_equal_svs;
  assign nor_692_nl = ~(FpAdd_6U_10U_is_a_greater_oif_aelse_acc_2_itm_10_1 | (~ inp_lookup_3_FpAdd_6U_10U_is_a_greater_oif_equal_tmp));
  assign mux_tmp_1837 = MUX_s_1_2_2((and_3053_nl), (nand_241_nl), nor_692_nl);
  assign or_dcpl_286 = mux_tmp_1837 | reg_inp_lookup_3_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse;
  assign and_dcpl_949 = or_dcpl_286 & and_dcpl_947 & or_11_cse;
  assign and_dcpl_954 = (~ mux_tmp_1837) & (cfg_precision_1_sva_st_113==2'b10) &
      (chn_inp_in_crt_sva_10_739_736_1[2]) & (~ reg_inp_lookup_3_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse)
      & or_11_cse;
  assign and_dcpl_955 = ((cfg_precision_1_sva_st_113!=2'b10) | (~ (chn_inp_in_crt_sva_10_739_736_1[2])))
      & or_11_cse;
  assign and_dcpl_958 = (cfg_precision_1_sva_st_125==2'b10) & (chn_inp_in_crt_sva_10_739_736_1[3])
      & or_11_cse;
  assign nor_696_nl = ~(FpAdd_6U_10U_is_a_greater_oif_aelse_acc_3_itm_10_1 | (~ inp_lookup_4_FpAdd_6U_10U_is_a_greater_oif_equal_tmp));
  assign mux_tmp_1838 = MUX_s_1_2_2((nor_696_nl), inp_lookup_4_FpAdd_6U_10U_is_a_greater_oif_equal_svs,
      reg_inp_lookup_4_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse);
  assign or_dcpl_289 = mux_tmp_1838 | reg_inp_lookup_4_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse;
  assign and_dcpl_959 = or_dcpl_289 & and_dcpl_958;
  assign and_dcpl_961 = (~ mux_tmp_1838) & (~ reg_inp_lookup_4_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse)
      & and_dcpl_958;
  assign and_dcpl_962 = (or_dcpl_257 | (~ (chn_inp_in_crt_sva_10_739_736_1[3])))
      & or_11_cse;
  assign or_dcpl_294 = (~ main_stage_v_8) | (cfg_precision_1_sva_st_85[0]);
  assign or_dcpl_295 = or_dcpl_294 | (~ (cfg_precision_1_sva_st_85[1]));
  assign or_dcpl_336 = (~ main_stage_v_7) | (cfg_precision_1_sva_st_84[0]);
  assign or_dcpl_342 = (~ main_stage_v_6) | (cfg_precision_1_sva_st_83[0]);
  assign or_dcpl_357 = ~(main_stage_v_6 & (chn_inp_in_crt_sva_6_739_736_1[1]));
  assign or_dcpl_409 = and_dcpl_78 | (~ main_stage_v_4);
  assign and_dcpl_1007 = or_5809_cse & (cfg_precision_1_sva_st_80==2'b10) & (~ (chn_inp_in_crt_sva_3_739_736_1[3]))
      & main_stage_v_3 & or_11_cse;
  assign and_dcpl_1009 = and_dcpl_423 & (~ (chn_inp_in_crt_sva_2_739_736_1[3])) &
      and_dcpl_419;
  assign mux_tmp_1845 = MUX_s_1_2_2((chn_inp_in_crt_sva_2_739_736_1[2]), (chn_inp_in_crt_sva_1_739_395_1[343]),
      or_11_cse);
  assign and_dcpl_1060 = or_11_cse & (~ (cfg_precision_rsci_d[0]));
  assign or_dcpl_499 = (chn_inp_in_rsci_d_mxwt[344:342]!=3'b111) | (~((chn_inp_in_rsci_d_mxwt[346:345]==2'b11)
      & IsDenorm_5U_10U_3_or_tmp));
  assign or_dcpl_542 = (chn_inp_in_rsci_d_mxwt[360:358]!=3'b111) | (~((chn_inp_in_rsci_d_mxwt[362:361]==2'b11)
      & IsDenorm_5U_10U_3_or_1_tmp));
  assign or_dcpl_585 = (chn_inp_in_rsci_d_mxwt[376:374]!=3'b111) | (~((chn_inp_in_rsci_d_mxwt[378:377]==2'b11)
      & IsDenorm_5U_10U_3_or_2_tmp));
  assign or_dcpl_628 = (chn_inp_in_rsci_d_mxwt[392:390]!=3'b111) | (~((chn_inp_in_rsci_d_mxwt[394:393]==2'b11)
      & IsDenorm_5U_10U_3_or_3_tmp));
  assign or_dcpl_630 = or_2_cse | (~ chn_inp_in_rsci_bawt);
  assign or_dcpl_631 = or_dcpl_630 | and_dcpl_78 | (chn_inp_in_rsci_d_mxwt[736]);
  assign or_dcpl_634 = or_dcpl_630 | and_dcpl_78 | (chn_inp_in_rsci_d_mxwt[737]);
  assign or_dcpl_637 = or_dcpl_630 | and_dcpl_78 | (chn_inp_in_rsci_d_mxwt[738]);
  assign or_dcpl_640 = or_dcpl_630 | and_dcpl_78 | (chn_inp_in_rsci_d_mxwt[739]);
  assign and_dcpl_1217 = and_4210_cse & IsNaN_8U_23U_land_lpi_1_dfm_4;
  assign and_dcpl_1219 = and_4210_cse & (~ IsNaN_8U_23U_land_lpi_1_dfm_4);
  assign and_dcpl_1224 = IsNaN_8U_23U_land_3_lpi_1_dfm_4 & (chn_inp_in_crt_sva_1_739_395_1[343])
      & or_11_cse;
  assign and_dcpl_1226 = (~ IsNaN_8U_23U_land_3_lpi_1_dfm_4) & (chn_inp_in_crt_sva_1_739_395_1[343])
      & or_11_cse;
  assign and_dcpl_1230 = IsNaN_8U_23U_land_1_lpi_1_dfm_st_3 & (chn_inp_in_crt_sva_1_739_395_1[341])
      & or_11_cse;
  assign and_dcpl_1232 = (~ IsNaN_8U_23U_land_1_lpi_1_dfm_st_3) & (chn_inp_in_crt_sva_1_739_395_1[341])
      & or_11_cse;
  assign or_dcpl_660 = and_dcpl_78 | (~ main_stage_v_2);
  assign and_dcpl_1243 = (~ IsNaN_6U_10U_4_nor_tmp) & IsNaN_8U_23U_land_1_lpi_1_dfm_st_4;
  assign and_dcpl_1247 = (inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_4_0_1[4]) & (inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_4_0_1[0]);
  assign and_dcpl_1252 = inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_6_5_1 & (~ IsNaN_6U_10U_4_nor_1_tmp);
  assign and_dcpl_1256 = (inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_6_4_0_1[1:0]==2'b11);
  assign and_dcpl_1261 = inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_6_5_1 & (~ IsNaN_6U_10U_4_nor_2_tmp);
  assign and_dcpl_1265 = (inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_6_4_0_1[1:0]==2'b11);
  assign and_dcpl_1270 = inp_lookup_else_if_a0_15_10_lpi_1_dfm_6_5_1 & (~ IsNaN_6U_10U_4_nor_3_tmp);
  assign and_dcpl_1274 = (inp_lookup_else_if_a0_15_10_lpi_1_dfm_6_4_0_1[1:0]==2'b11);
  assign or_dcpl_699 = and_dcpl_78 | (~ main_stage_v_3);
  assign and_dcpl_1335 = FpAdd_6U_10U_1_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0 & or_11_cse;
  assign or_dcpl_727 = ~((~ FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_itm_10) & IsNaN_8U_23U_2_land_1_lpi_1_dfm_9);
  assign and_dcpl_1338 = or_dcpl_727 & (~ IsNaN_8U_23U_3_land_1_lpi_1_dfm_6) & (~
      (chn_inp_in_crt_sva_5_739_736_1[0])) & or_11_cse;
  assign and_dcpl_1348 = FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0 & or_11_cse;
  assign or_dcpl_732 = ~((~ FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_1_itm_10) &
      IsNaN_8U_23U_2_land_2_lpi_1_dfm_9);
  assign and_dcpl_1351 = or_dcpl_732 & (~ IsNaN_8U_23U_3_land_2_lpi_1_dfm_6) & (~
      (chn_inp_in_crt_sva_5_739_736_1[1])) & or_11_cse;
  assign and_dcpl_1361 = FpAdd_6U_10U_1_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0 & or_11_cse;
  assign or_dcpl_737 = ~((~ FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_2_itm_10) &
      IsNaN_8U_23U_2_land_3_lpi_1_dfm_9);
  assign and_dcpl_1364 = or_dcpl_737 & (~ IsNaN_8U_23U_3_land_3_lpi_1_dfm_6) & (~
      (chn_inp_in_crt_sva_5_739_736_1[2])) & or_11_cse;
  assign mux_tmp_1861 = MUX_s_1_2_2(nor_1130_cse, (~ IsNaN_8U_23U_2_land_lpi_1_dfm_st_8),
      FpAdd_6U_10U_1_is_a_greater_oif_aelse_acc_3_itm_10);
  assign and_dcpl_1373 = mux_tmp_1861 & IsNaN_8U_23U_2_land_lpi_1_dfm_9;
  assign and_dcpl_1374 = (and_dcpl_1373 | IsNaN_8U_23U_3_land_lpi_1_dfm_5) & or_11_cse;
  assign or_dcpl_742 = ~(mux_tmp_1861 & IsNaN_8U_23U_2_land_lpi_1_dfm_9);
  assign and_dcpl_1377 = or_dcpl_742 & (~ IsNaN_8U_23U_3_land_lpi_1_dfm_5) & (~ (chn_inp_in_crt_sva_5_739_736_1[3]))
      & or_11_cse;
  assign mux_tmp_1862 = MUX_s_1_2_2((chn_inp_in_crt_sva_7_739_736_1[2]), (chn_inp_in_crt_sva_6_739_736_1[2]),
      or_11_cse);
  assign and_dcpl_1404 = or_11_cse & IsNaN_6U_10U_land_1_lpi_1_dfm_5;
  assign and_dcpl_1415 = or_11_cse & IsNaN_6U_10U_land_2_lpi_1_dfm_5;
  assign and_dcpl_1426 = or_11_cse & IsNaN_6U_10U_land_3_lpi_1_dfm_5;
  assign and_dcpl_1437 = or_11_cse & IsNaN_6U_10U_land_lpi_1_dfm_5;
  assign and_dcpl_1448 = or_11_cse & (~ IsNaN_6U_10U_2_land_lpi_1_dfm_24);
  assign and_dcpl_1450 = or_11_cse & (~ IsNaN_6U_10U_2_land_3_lpi_1_dfm_24);
  assign and_dcpl_1452 = or_11_cse & (~ IsNaN_6U_10U_2_land_2_lpi_1_dfm_24);
  assign and_dcpl_1454 = or_11_cse & (~ IsNaN_6U_10U_2_land_1_lpi_1_dfm_24);
  assign and_dcpl_1473 = or_11_cse & (chn_inp_in_crt_sva_10_739_736_1[0]);
  assign and_dcpl_1481 = (~ mux_tmp_1835) & main_stage_v_10 & and_dcpl_927 & (~ reg_inp_lookup_1_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse)
      & and_dcpl_1473;
  assign and_dcpl_1484 = main_stage_v_10 & (cfg_precision_1_sva_st_101==2'b10);
  assign and_dcpl_1488 = and_dcpl_943 & and_dcpl_1484 & and_dcpl_941;
  assign and_dcpl_1497 = (~ mux_tmp_1837) & main_stage_v_10 & and_dcpl_947 & or_11_cse
      & (~ reg_inp_lookup_3_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse);
  assign and_dcpl_1504 = ~((cfg_precision_1_sva_st_91[0]) | (chn_inp_in_crt_sva_2_739_736_1[3]));
  assign and_dcpl_1534 = (chn_inp_in_rsci_d_mxwt[312:311]==2'b11);
  assign or_dcpl_818 = (chn_inp_in_rsci_d_mxwt[313:311]!=3'b111) | (~((chn_inp_in_rsci_d_mxwt[310])
      & (chn_inp_in_rsci_d_mxwt[314]) & IsDenorm_5U_10U_2_or_2_tmp));
  assign and_dcpl_1541 = (FpFractionToFloat_35U_6U_10U_1_mux_tmp[4:3]==2'b11);
  assign and_dcpl_1545 = (FpFractionToFloat_35U_6U_10U_1_mux_tmp[2:0]==3'b111);
  assign and_dcpl_1556 = (FpFractionToFloat_35U_6U_10U_1_mux_40_tmp[2:0]==3'b111);
  assign and_dcpl_1566 = (FpFractionToFloat_35U_6U_10U_1_mux_41_tmp[4]) & (FpFractionToFloat_35U_6U_10U_1_mux_41_tmp[2])
      & (FpFractionToFloat_35U_6U_10U_1_mux_41_tmp[0]);
  assign and_dcpl_1577 = (FpFractionToFloat_35U_6U_10U_1_mux_42_tmp[2:0]==3'b111);
  assign or_tmp_4282 = (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[0]) |
      (cfg_precision_1_sva_st_80!=2'b10) | IsNaN_6U_10U_7_land_1_lpi_1_dfm_6 | IsNaN_6U_10U_6_land_1_lpi_1_dfm_5;
  assign and_dcpl_1588 = (~ (chn_inp_in_crt_sva_2_739_736_1[1])) & main_stage_v_2
      & or_11_cse;
  assign and_dcpl_1596 = main_stage_v_2 & (~ (chn_inp_in_crt_sva_2_739_736_1[2]))
      & or_11_cse;
  assign and_dcpl_1617 = IsNaN_6U_10U_8_land_lpi_1_dfm_4 & (~ (chn_inp_in_crt_sva_5_739_736_1[3]))
      & or_11_cse;
  assign and_dcpl_1619 = (~ IsNaN_6U_10U_8_land_lpi_1_dfm_4) & (~ (chn_inp_in_crt_sva_5_739_736_1[3]))
      & or_11_cse;
  assign and_dcpl_1624 = IsNaN_6U_10U_8_land_3_lpi_1_dfm_4 & (~ (chn_inp_in_crt_sva_5_739_736_1[2]))
      & or_11_cse;
  assign and_dcpl_1626 = (~ IsNaN_6U_10U_8_land_3_lpi_1_dfm_4) & (~ (chn_inp_in_crt_sva_5_739_736_1[2]))
      & or_11_cse;
  assign and_dcpl_1632 = IsNaN_6U_10U_8_land_2_lpi_1_dfm_4 & (~ (chn_inp_in_crt_sva_5_739_736_1[1]))
      & or_11_cse;
  assign and_dcpl_1634 = (~ IsNaN_6U_10U_8_land_2_lpi_1_dfm_4) & (~ (chn_inp_in_crt_sva_5_739_736_1[1]))
      & or_11_cse;
  assign and_dcpl_1639 = IsNaN_6U_10U_8_land_1_lpi_1_dfm_6 & (~ (chn_inp_in_crt_sva_5_739_736_1[0]))
      & or_11_cse;
  assign and_dcpl_1641 = (~ IsNaN_6U_10U_8_land_1_lpi_1_dfm_6) & (~ (chn_inp_in_crt_sva_5_739_736_1[0]))
      & or_11_cse;
  assign or_dcpl_897 = or_2010_cse | (chn_inp_in_crt_sva_1_739_395_1[341]);
  assign or_dcpl_903 = or_2010_cse | (chn_inp_in_crt_sva_1_739_395_1[342]);
  assign or_dcpl_906 = and_dcpl_78 | (chn_inp_in_crt_sva_1_739_395_1[343]);
  assign or_dcpl_913 = and_dcpl_78 | (chn_inp_in_crt_sva_1_739_395_1[344]);
  assign and_dcpl_1722 = or_11_cse & (chn_inp_in_crt_sva_10_739_736_1[3]);
  assign and_dcpl_1731 = (~ mux_tmp_1838) & main_stage_v_10 & (~ reg_inp_lookup_4_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse)
      & (cfg_precision_1_sva_st_125==2'b10) & and_dcpl_1722;
  assign and_dcpl_1758 = (chn_inp_in_rsci_d_mxwt[346:342]==5'b11111) & IsDenorm_5U_10U_3_or_tmp;
  assign and_dcpl_1759 = and_dcpl_142 & chn_inp_in_rsci_bawt;
  assign and_dcpl_1760 = and_dcpl_1759 & and_dcpl_105;
  assign and_dcpl_1764 = and_dcpl_1759 & (~ (chn_inp_in_rsci_d_mxwt[736])) & chn_inp_out_rsci_bawt
      & reg_chn_inp_out_rsci_ld_core_psct_cse;
  assign and_dcpl_1772 = (chn_inp_in_rsci_d_mxwt[362:358]==5'b11111) & IsDenorm_5U_10U_3_or_1_tmp;
  assign and_dcpl_1773 = and_dcpl_1759 & and_dcpl_176;
  assign and_dcpl_1777 = and_dcpl_1759 & (~ (chn_inp_in_rsci_d_mxwt[737])) & chn_inp_out_rsci_bawt
      & reg_chn_inp_out_rsci_ld_core_psct_cse;
  assign and_dcpl_1785 = (chn_inp_in_rsci_d_mxwt[378:374]==5'b11111) & IsDenorm_5U_10U_3_or_2_tmp;
  assign and_dcpl_1786 = and_dcpl_1759 & and_dcpl_246;
  assign and_dcpl_1790 = and_dcpl_1759 & (~ (chn_inp_in_rsci_d_mxwt[738])) & chn_inp_out_rsci_bawt
      & reg_chn_inp_out_rsci_ld_core_psct_cse;
  assign and_dcpl_1798 = (chn_inp_in_rsci_d_mxwt[394:390]==5'b11111) & IsDenorm_5U_10U_3_or_3_tmp;
  assign and_dcpl_1799 = and_dcpl_1759 & and_dcpl_316;
  assign and_dcpl_1803 = and_dcpl_1759 & (~ (chn_inp_in_rsci_d_mxwt[739])) & chn_inp_out_rsci_bawt
      & reg_chn_inp_out_rsci_ld_core_psct_cse;
  assign and_dcpl_1852 = and_dcpl_142 & (chn_inp_in_rsci_d_mxwt[736]);
  assign and_dcpl_1853 = and_dcpl_1852 & or_11_cse;
  assign and_dcpl_1854 = (or_2_cse | (~ (chn_inp_in_rsci_d_mxwt[736]))) & or_11_cse;
  assign and_dcpl_1856 = and_dcpl_142 & (chn_inp_in_rsci_d_mxwt[737]) & or_11_cse;
  assign and_dcpl_1857 = (or_2_cse | (~ (chn_inp_in_rsci_d_mxwt[737]))) & or_11_cse;
  assign and_dcpl_1858 = and_dcpl_142 & (chn_inp_in_rsci_d_mxwt[738]);
  assign and_dcpl_1859 = and_dcpl_1858 & or_11_cse;
  assign and_dcpl_1860 = (or_2_cse | (~ (chn_inp_in_rsci_d_mxwt[738]))) & or_11_cse;
  assign and_dcpl_1862 = and_dcpl_142 & (chn_inp_in_rsci_d_mxwt[739]) & or_11_cse;
  assign and_dcpl_1863 = (or_2_cse | (~ (chn_inp_in_rsci_d_mxwt[739]))) & or_11_cse;
  assign or_dcpl_985 = (~(IsDenorm_5U_10U_or_tmp & (chn_inp_in_rsci_d_mxwt[407:406]==2'b11)))
      | (chn_inp_in_rsci_d_mxwt[410:408]!=3'b111);
  assign or_dcpl_990 = (chn_inp_in_rsci_d_mxwt[424:422]!=3'b111) | (~((chn_inp_in_rsci_d_mxwt[426:425]==2'b11)
      & IsDenorm_5U_10U_or_1_tmp));
  assign or_dcpl_995 = (~((chn_inp_in_rsci_d_mxwt[442]) & (chn_inp_in_rsci_d_mxwt[441])
      & (chn_inp_in_rsci_d_mxwt[438]))) | (~((chn_inp_in_rsci_d_mxwt[440]) & IsDenorm_5U_10U_or_2_tmp
      & (chn_inp_in_rsci_d_mxwt[439])));
  assign or_dcpl_1000 = (chn_inp_in_rsci_d_mxwt[456:454]!=3'b111) | (~((chn_inp_in_rsci_d_mxwt[458:457]==2'b11)
      & IsDenorm_5U_10U_or_3_tmp));
  assign or_dcpl_1005 = (chn_inp_in_rsci_d_mxwt[280:278]!=3'b111) | (~((chn_inp_in_rsci_d_mxwt[282:281]==2'b11)
      & IsDenorm_5U_10U_2_or_tmp));
  assign or_dcpl_1010 = (chn_inp_in_rsci_d_mxwt[296:294]!=3'b111) | (~((chn_inp_in_rsci_d_mxwt[298:297]==2'b11)
      & IsDenorm_5U_10U_2_or_1_tmp));
  assign and_dcpl_1927 = and_dcpl_1534 & (chn_inp_in_rsci_d_mxwt[313]) & (chn_inp_in_rsci_d_mxwt[310])
      & (chn_inp_in_rsci_d_mxwt[314]) & IsDenorm_5U_10U_2_or_2_tmp;
  assign or_dcpl_1015 = (~((chn_inp_in_rsci_d_mxwt[329]) & (chn_inp_in_rsci_d_mxwt[326])
      & (chn_inp_in_rsci_d_mxwt[327]))) | (~((chn_inp_in_rsci_d_mxwt[328]) & (chn_inp_in_rsci_d_mxwt[330])
      & IsDenorm_5U_10U_2_or_3_tmp));
  assign and_dcpl_1947 = (or_2_cse | (~ chn_inp_in_rsci_bawt) | (~ (chn_inp_in_rsci_d_mxwt[739])))
      & and_4210_cse;
  assign and_dcpl_1953 = and_dcpl_1759 & and_dcpl_65;
  assign and_dcpl_1957 = (chn_inp_in_rsci_d_mxwt[410:408]==3'b111);
  assign and_dcpl_1961 = and_dcpl_1759 & and_dcpl_38;
  assign and_dcpl_1979 = (chn_inp_in_rsci_d_mxwt[426:422]==5'b11111) & IsDenorm_5U_10U_or_1_tmp;
  assign and_dcpl_1980 = and_dcpl_1759 & and_dcpl_49;
  assign and_dcpl_1984 = and_dcpl_1759 & (chn_inp_in_rsci_d_mxwt[737]) & chn_inp_out_rsci_bawt
      & reg_chn_inp_out_rsci_ld_core_psct_cse;
  assign and_dcpl_1989 = (chn_inp_in_rsci_d_mxwt[440]) & IsDenorm_5U_10U_or_2_tmp
      & (chn_inp_in_rsci_d_mxwt[439]);
  assign and_dcpl_1993 = and_dcpl_1759 & and_dcpl_57;
  assign and_dcpl_2005 = and_dcpl_1759 & (chn_inp_in_rsci_d_mxwt[738]) & chn_inp_out_rsci_bawt
      & reg_chn_inp_out_rsci_ld_core_psct_cse;
  assign and_dcpl_2011 = (chn_inp_in_rsci_d_mxwt[458:454]==5'b11111) & IsDenorm_5U_10U_or_3_tmp;
  assign and_dcpl_2015 = and_dcpl_1759 & (chn_inp_in_rsci_d_mxwt[739]) & chn_inp_out_rsci_bawt
      & reg_chn_inp_out_rsci_ld_core_psct_cse;
  assign or_tmp_4339 = or_11_cse & chn_inp_in_rsci_bawt & (fsm_output[1]);
  assign nor_725_nl = ~((cfg_precision_1_sva_st_91[1]) | and_dcpl_633);
  assign or_4697_nl = (~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[3]) |
      (cfg_precision_1_sva_st_91[0]);
  assign mux_1920_nl = MUX_s_1_2_2((nor_725_nl), or_tmp_4220, or_4697_nl);
  assign mux_1921_nl = MUX_s_1_2_2(or_5809_cse, (mux_1920_nl), main_stage_v_3);
  assign or_4702_nl = main_stage_v_3 | (~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[3])
      | (cfg_precision_1_sva_st_91!=2'b10);
  assign mux_1922_nl = MUX_s_1_2_2((or_4702_nl), (mux_1921_nl), or_11_cse);
  assign or_tmp_4457 = (mux_1922_nl) | (fsm_output[0]);
  assign chn_inp_in_rsci_ld_core_psct_mx0c0 = main_stage_en_1 | (fsm_output[0]);
  assign chn_inp_out_rsci_d_0_mx0c1 = main_stage_v_12 & (~ (chn_inp_in_crt_sva_12_739_736_1[0]))
      & or_11_cse;
  assign chn_inp_out_rsci_d_32_mx0c1 = main_stage_v_12 & (~ (chn_inp_in_crt_sva_12_739_736_1[1]))
      & or_11_cse;
  assign chn_inp_out_rsci_d_64_mx0c1 = main_stage_v_12 & (~ (chn_inp_in_crt_sva_12_739_736_1[2]))
      & or_11_cse;
  assign chn_inp_out_rsci_d_96_mx0c1 = main_stage_v_12 & (~ (chn_inp_in_crt_sva_12_739_736_1[3]))
      & or_11_cse;
  assign main_stage_v_1_mx0c1 = (~ chn_inp_in_rsci_bawt) & main_stage_v_1 & or_11_cse;
  assign FpFractionToFloat_35U_6U_10U_1_o_mant_1_lpi_1_dfm_6_mx0c1 = (and_dcpl_173
      | inp_lookup_1_FpMantRNE_36U_11U_1_else_and_tmp) & or_11_cse;
  assign FpFractionToFloat_35U_6U_10U_1_o_mant_2_lpi_1_dfm_6_mx0c1 = (and_dcpl_243
      | inp_lookup_2_FpMantRNE_36U_11U_1_else_and_tmp) & or_11_cse;
  assign FpFractionToFloat_35U_6U_10U_1_o_mant_3_lpi_1_dfm_6_mx0c1 = (and_dcpl_313
      | inp_lookup_3_FpMantRNE_36U_11U_1_else_and_tmp) & or_11_cse;
  assign FpFractionToFloat_35U_6U_10U_1_o_mant_lpi_1_dfm_6_mx0c1 = (and_dcpl_383
      | inp_lookup_4_FpMantRNE_36U_11U_1_else_and_tmp) & or_11_cse;
  assign main_stage_v_2_mx0c1 = (~ main_stage_v_1) & main_stage_v_2 & or_11_cse;
  assign main_stage_v_3_mx0c1 = (~ main_stage_v_2) & main_stage_v_3 & or_11_cse;
  assign main_stage_v_4_mx0c1 = (~ main_stage_v_3) & main_stage_v_4 & or_11_cse;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_9_mx0c0 = and_dcpl_615
      & (cfg_precision_1_sva_st_80[1]) & IsNaN_6U_10U_5_land_3_lpi_1_dfm_5 & and_dcpl_613;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_9_mx0c2 = and_dcpl_615
      & (cfg_precision_1_sva_st_80[1]) & (~ IsNaN_6U_10U_5_land_3_lpi_1_dfm_5) &
      and_dcpl_613;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_9_mx0c3 = IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_15
      & (~ (cfg_precision_1_sva_st_80[0])) & and_dcpl_526 & and_dcpl_560;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_9_1_mx0c0 = and_dcpl_584
      & and_dcpl_642 & and_dcpl_560;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_9_1_mx0c2 = and_dcpl_584
      & and_dcpl_645 & and_dcpl_560;
  assign main_stage_v_5_mx0c1 = main_stage_v_5 & (~ main_stage_v_4) & or_11_cse;
  assign main_stage_v_6_mx0c1 = (~ main_stage_v_5) & main_stage_v_6 & or_11_cse;
  assign main_stage_v_7_mx0c1 = (~ main_stage_v_6) & main_stage_v_7 & or_11_cse;
  assign main_stage_v_8_mx0c1 = main_stage_v_8 & (~ main_stage_v_7) & or_11_cse;
  assign main_stage_v_9_mx0c1 = (~ main_stage_v_8) & main_stage_v_9 & or_11_cse;
  assign main_stage_v_10_mx0c1 = (~ main_stage_v_9) & main_stage_v_10 & or_11_cse;
  assign main_stage_v_11_mx0c1 = (~ main_stage_v_10) & main_stage_v_11 & or_11_cse;
  assign main_stage_v_12_mx0c1 = (~ main_stage_v_11) & main_stage_v_12 & or_11_cse;
  assign FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx0c0 = or_tmp_899 & main_stage_v_6
      & (cfg_precision_1_sva_st_83==2'b10) & nor_tmp_686;
  assign FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx0c1 = or_tmp_899 & main_stage_v_6
      & (cfg_precision_1_sva_st_83==2'b10) & (chn_inp_in_crt_sva_6_739_736_1[2])
      & (~ IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_4) & or_11_cse;
  assign FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx0c2 = main_stage_v_5 & (cfg_precision_1_sva_st_82==2'b10)
      & and_dcpl_712;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_3_mx0c1 = (or_dcpl_499
      & and_dcpl_1760 & (fsm_output[1])) | (or_dcpl_499 & and_dcpl_1764);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_3_mx0c1 = (or_dcpl_542
      & and_dcpl_1773 & (fsm_output[1])) | (or_dcpl_542 & and_dcpl_1777);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_3_lpi_1_dfm_3_mx0c1 = (or_dcpl_585
      & and_dcpl_1786 & (fsm_output[1])) | (or_dcpl_585 & and_dcpl_1790);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_3_mx0c1 = (or_dcpl_628
      & and_dcpl_1799 & (fsm_output[1])) | (or_dcpl_628 & and_dcpl_1803);
  assign FpAdd_8U_23U_o_sign_lpi_1_dfm_1_mx0c0 = and_dcpl_1947 & IsNaN_8U_23U_land_lpi_1_dfm_4
      & main_stage_v_1 & (chn_inp_in_crt_sva_1_739_395_1[344]) & or_11_cse;
  assign FpAdd_8U_23U_o_sign_lpi_1_dfm_1_mx0c1 = and_dcpl_1947 & (~ IsNaN_8U_23U_land_lpi_1_dfm_4)
      & main_stage_v_1 & (chn_inp_in_crt_sva_1_739_395_1[344]) & or_11_cse;
  assign FpAdd_8U_23U_o_sign_lpi_1_dfm_1_mx0c2 = and_dcpl_1953 & (fsm_output[1]);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_3_mx0c1 = (or_dcpl_985
      & and_dcpl_1961 & (fsm_output[1])) | (or_dcpl_985 & and_dcpl_1759 & (chn_inp_in_rsci_d_mxwt[736])
      & chn_inp_out_rsci_bawt & reg_chn_inp_out_rsci_ld_core_psct_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_3_mx0c1 = (or_dcpl_990
      & and_dcpl_1980 & (fsm_output[1])) | (or_dcpl_990 & and_dcpl_1984);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_3_mx0c1 = (or_dcpl_995
      & and_dcpl_1993 & (fsm_output[1])) | (or_dcpl_995 & and_dcpl_2005);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_3_mx0c1 = (or_dcpl_1000
      & and_dcpl_1953 & (fsm_output[1])) | (or_dcpl_1000 & and_dcpl_2015);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_3_mx0c1 = (or_dcpl_818
      & and_dcpl_1993 & (fsm_output[1])) | (or_dcpl_818 & and_dcpl_2005);
  assign nl_FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_nl = ({1'b1 , (chn_inp_in_crt_sva_3_127_0_1[22:0])})
      + conv_u2u_23_24(~ FpAdd_8U_23U_o_mant_1_lpi_1_dfm_2_mx2) + 24'b1;
  assign FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_nl = nl_FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_nl[23:0];
  assign FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_nl));
  assign nl_FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_1_nl = ({1'b1 , (chn_inp_in_crt_sva_3_127_0_1[54:32])})
      + conv_u2u_23_24(~ FpAdd_8U_23U_o_mant_2_lpi_1_dfm_2_mx2) + 24'b1;
  assign FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_1_nl = nl_FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_1_nl[23:0];
  assign FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_1_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_1_nl));
  assign nl_FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_2_nl = ({1'b1 , (chn_inp_in_crt_sva_3_127_0_1[86:64])})
      + conv_u2u_23_24(~ FpAdd_8U_23U_o_mant_3_lpi_1_dfm_2_mx2) + 24'b1;
  assign FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_2_nl = nl_FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_2_nl[23:0];
  assign FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_2_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_2_nl));
  assign nl_FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_3_nl = ({1'b1 , (chn_inp_in_crt_sva_3_127_0_1[118:96])})
      + conv_u2u_23_24(~ FpAdd_8U_23U_o_mant_lpi_1_dfm_2_mx2) + 24'b1;
  assign FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_3_nl = nl_FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_3_nl[23:0];
  assign FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_3_itm_23_1 = readslicef_24_1_23((FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_3_nl));
  assign nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_24})
      + conv_u2u_10_11(~ FpMul_6U_10U_o_mant_1_lpi_1_dfm_7) + 11'b1;
  assign FpAdd_6U_10U_is_a_greater_oif_aelse_acc_nl = nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_nl[10:0];
  assign FpAdd_6U_10U_is_a_greater_oif_aelse_acc_itm_10_1 = readslicef_11_1_10((FpAdd_6U_10U_is_a_greater_oif_aelse_acc_nl));
  assign nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_1_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_24})
      + conv_u2u_10_11(~ FpMul_6U_10U_o_mant_2_lpi_1_dfm_7) + 11'b1;
  assign FpAdd_6U_10U_is_a_greater_oif_aelse_acc_1_nl = nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_1_nl[10:0];
  assign FpAdd_6U_10U_is_a_greater_oif_aelse_acc_1_itm_10_1 = readslicef_11_1_10((FpAdd_6U_10U_is_a_greater_oif_aelse_acc_1_nl));
  assign nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_2_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_27})
      + conv_u2u_10_11(~ FpMul_6U_10U_o_mant_3_lpi_1_dfm_7) + 11'b1;
  assign FpAdd_6U_10U_is_a_greater_oif_aelse_acc_2_nl = nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_2_nl[10:0];
  assign FpAdd_6U_10U_is_a_greater_oif_aelse_acc_2_itm_10_1 = readslicef_11_1_10((FpAdd_6U_10U_is_a_greater_oif_aelse_acc_2_nl));
  assign nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_3_nl = ({1'b1 , FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_24})
      + conv_u2u_10_11(~ FpMul_6U_10U_o_mant_lpi_1_dfm_7) + 11'b1;
  assign FpAdd_6U_10U_is_a_greater_oif_aelse_acc_3_nl = nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_3_nl[10:0];
  assign FpAdd_6U_10U_is_a_greater_oif_aelse_acc_3_itm_10_1 = readslicef_11_1_10((FpAdd_6U_10U_is_a_greater_oif_aelse_acc_3_nl));
  assign inp_lookup_if_and_m1c_9 = (~ inp_lookup_if_unequal_tmp_1_mx0w0) & and_dcpl_1722;
  assign inp_lookup_if_and_m1c_10 = (~ IsNaN_6U_10U_2_land_lpi_1_dfm_24) & inp_lookup_if_and_m1c_9;
  assign inp_lookup_if_and_m1c_11 = (~ IsNaN_6U_10U_3_land_lpi_1_dfm_6) & inp_lookup_if_and_m1c_10;
  assign and_1942_m1c = or_11_cse & (chn_inp_in_crt_sva_10_739_736_1[2]);
  assign inp_lookup_if_and_m1c_6 = (~ inp_lookup_if_unequal_tmp_1_mx0w0) & and_1942_m1c;
  assign inp_lookup_if_and_m1c_7 = (~ IsNaN_6U_10U_2_land_3_lpi_1_dfm_24) & inp_lookup_if_and_m1c_6;
  assign inp_lookup_if_and_m1c_8 = (~ IsNaN_6U_10U_3_land_3_lpi_1_dfm_6) & inp_lookup_if_and_m1c_7;
  assign and_1944_m1c = or_11_cse & (chn_inp_in_crt_sva_10_739_736_1[1]);
  assign inp_lookup_if_and_m1c_3 = (~ inp_lookup_if_unequal_tmp_1_mx0w0) & and_1944_m1c;
  assign inp_lookup_if_and_m1c_4 = (~ IsNaN_6U_10U_2_land_2_lpi_1_dfm_24) & inp_lookup_if_and_m1c_3;
  assign inp_lookup_if_and_m1c_5 = (~ IsNaN_6U_10U_3_land_2_lpi_1_dfm_6) & inp_lookup_if_and_m1c_4;
  assign inp_lookup_if_and_m1c = (~ inp_lookup_if_unequal_tmp_1_mx0w0) & and_dcpl_1473;
  assign inp_lookup_if_and_m1c_1 = (~ IsNaN_6U_10U_2_land_1_lpi_1_dfm_24) & inp_lookup_if_and_m1c;
  assign inp_lookup_if_and_m1c_2 = (~ IsNaN_6U_10U_3_land_1_lpi_1_dfm_6) & inp_lookup_if_and_m1c_1;
  assign and_2307_m1c = (chn_inp_in_crt_sva_4_739_736_1[0]) & (~ IsNaN_6U_10U_5_land_1_lpi_1_dfm_6)
      & or_11_cse;
  assign and_m1c_3 = (~ FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_4) & and_2307_m1c;
  assign and_2311_m1c = (~ IsNaN_6U_10U_5_land_2_lpi_1_dfm_6) & (chn_inp_in_crt_sva_4_739_736_1[1])
      & or_11_cse;
  assign and_m1c_2 = (~ FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_4) & and_2311_m1c;
  assign and_2315_m1c = (chn_inp_in_crt_sva_4_739_736_1[2]) & (~ IsNaN_6U_10U_5_land_3_lpi_1_dfm_6)
      & or_11_cse;
  assign and_m1c_1 = (~ FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_4) & and_2315_m1c;
  assign and_2319_m1c = (chn_inp_in_crt_sva_4_739_736_1[3]) & (~ FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_4)
      & or_11_cse;
  assign and_m1c = (~ IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0) & and_2319_m1c;
  assign and_2321_m1c = (~ or_3384_cse) & or_11_cse;
  assign IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_6 = (~ IsNaN_6U_10U_8_land_lpi_1_dfm_4)
      & and_2321_m1c;
  assign IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_7 = (~ IsNaN_6U_10U_9_land_lpi_1_dfm_6)
      & IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_6;
  assign IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_4 = (~ IsNaN_6U_10U_8_land_3_lpi_1_dfm_4)
      & and_2321_m1c;
  assign IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_5 = (~ IsNaN_6U_10U_9_land_3_lpi_1_dfm_6)
      & IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_4;
  assign IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_2 = (~ IsNaN_6U_10U_8_land_2_lpi_1_dfm_4)
      & and_2321_m1c;
  assign IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_3 = (~ IsNaN_6U_10U_9_land_2_lpi_1_dfm_6)
      & IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_2;
  assign IntShiftRight_69U_6U_32U_obits_fixed_and_m1c = (~ IsNaN_6U_10U_8_land_1_lpi_1_dfm_6)
      & and_2321_m1c;
  assign IntShiftRight_69U_6U_32U_obits_fixed_and_m1c_1 = (~ IsNaN_6U_10U_9_land_1_lpi_1_dfm_6)
      & IntShiftRight_69U_6U_32U_obits_fixed_and_m1c;
  assign chn_inp_in_rsci_oswt_unreg = or_tmp_4339;
  assign chn_inp_out_rsci_oswt_unreg = chn_inp_out_rsci_bawt & reg_chn_inp_out_rsci_ld_core_psct_cse;
  assign not_tmp_2674 = ~(or_5882_cse & FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_6_1_1
      & FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_6_0_1 & (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_9==4'b1111));
  assign or_tmp_4611 = ((FpFractionToFloat_35U_6U_10U_1_mux_tmp[4:3]==2'b11) & (IntLeadZero_35U_1_leading_sign_35_0_rtn_1_sva_2[5])
      & inp_lookup_1_FpMantRNE_36U_11U_1_else_and_svs_2 & FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_st_2
      & (FpFractionToFloat_35U_6U_10U_1_mux_tmp[2:0]==3'b111)) | not_tmp_2674;
  assign or_tmp_4615 = (((FpFractionToFloat_35U_6U_10U_1_o_mant_1_lpi_1_dfm_6[8:0]!=9'b000000000))
      & (FpFractionToFloat_35U_6U_10U_1_mux_tmp[4:3]==2'b11) & (IntLeadZero_35U_1_leading_sign_35_0_rtn_1_sva_2[5])
      & inp_lookup_1_FpMantRNE_36U_11U_1_else_and_svs_2 & FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_st_2
      & (FpFractionToFloat_35U_6U_10U_1_mux_tmp[2:0]==3'b111)) | not_tmp_2674;
  assign or_tmp_4620 = inp_lookup_1_FpMul_6U_10U_2_oelse_1_acc_itm_7 | IsZero_6U_10U_7_IsZero_6U_10U_7_and_itm_2
      | IsZero_6U_10U_6_IsZero_6U_10U_6_nor_tmp | (~ inp_lookup_1_FpMul_6U_10U_2_else_2_if_acc_itm_6);
  assign nor_tmp_708 = FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_6_1_1
      & FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_6_0_1 & (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_9==4'b1111);
  assign or_tmp_4625 = (FpFractionToFloat_35U_6U_10U_1_o_mant_2_lpi_1_dfm_6!=10'b0000000000)
      | (~ nor_tmp_708);
  assign or_tmp_4637 = inp_lookup_4_FpMul_6U_10U_2_oelse_1_acc_itm_7 | IsZero_6U_10U_7_IsZero_6U_10U_7_and_3_itm_2
      | IsZero_6U_10U_6_IsZero_6U_10U_6_nor_3_tmp | (~ inp_lookup_4_FpMul_6U_10U_2_else_2_if_acc_itm_6);
  assign and_dcpl_2185 = main_stage_v_4 & core_wen;
  assign or_tmp_4675 = (FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_8!=10'b0000000000);
  assign or_tmp_4685 = (FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_8!=10'b0000000000);
  assign or_tmp_4698 = (~(FpAdd_6U_10U_1_is_a_greater_acc_2_itm_6 | (~ inp_lookup_3_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp)))
      | mux_500_cse;
  assign or_tmp_4703 = (FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_8!=10'b0000000000);
  assign and_dcpl_2279 = core_wen & main_stage_v_11;
  assign and_dcpl_2318 = core_wen & main_stage_v_1;
  assign or_tmp_4714 = ~((chn_inp_in_crt_sva_1_739_395_1[344]) & (cfg_precision_1_sva_st_90==2'b10)
      & or_5695_itm);
  assign or_tmp_4721 = (cfg_precision_1_sva_st_90!=2'b10) | (~((chn_inp_in_crt_sva_1_739_395_1[343])
      & or_5694_itm));
  assign or_tmp_4726 = (cfg_precision_1_sva_st_90[0]) | (~((cfg_precision_1_sva_st_90[1])
      & (chn_inp_in_crt_sva_1_739_395_1[341]) & or_6042_cse));
  assign or_tmp_4730 = ~((chn_inp_in_crt_sva_1_739_395_1[342]) & (cfg_precision_1_sva_st_90==2'b10)
      & or_5693_itm);
  assign or_tmp_4737 = (chn_inp_in_crt_sva_6_739_736_1[2]) | (~ or_tmp_2703);
  assign or_tmp_4741 = (chn_inp_in_crt_sva_6_739_736_1[0]) | (~ or_tmp_2723);
  assign or_tmp_4745 = (chn_inp_in_crt_sva_6_739_736_1[1]) | (~ or_tmp_2738);
  assign or_tmp_4753 = (chn_inp_in_crt_sva_6_739_736_1[3]) | (~ or_tmp_2695);
  assign and_dcpl_2461 = core_wen & main_stage_v_10;
  assign and_dcpl_2487 = core_wen & main_stage_v_5;
  assign and_dcpl_2500 = core_wen & main_stage_v_9;
  assign and_dcpl_2528 = core_wen & main_stage_v_8;
  assign FpAdd_8U_23U_else_2_and_tmp = (fsm_output[1]) & (~ inp_lookup_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_4);
  assign FpAdd_8U_23U_else_2_and_tmp_1 = (fsm_output[1]) & (~ inp_lookup_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_4);
  assign FpAdd_8U_23U_else_2_and_tmp_2 = (fsm_output[1]) & (~ inp_lookup_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_4);
  assign FpAdd_8U_23U_else_2_and_tmp_3 = (fsm_output[1]) & (~ inp_lookup_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_4);
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp = (fsm_output[1]) & (~ FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_5);
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp_1 = (fsm_output[1]) & (~ FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2);
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp_2 = (fsm_output[1]) & (~ FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_5);
  assign FpAdd_8U_23U_a_right_shift_qelse_and_tmp_3 = (fsm_output[1]) & (~ FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_5);
  assign FpAdd_6U_10U_1_if_4_if_and_tmp = (fsm_output[1]) & (~ (chn_inp_in_crt_sva_7_739_736_1[0]));
  assign FpAdd_6U_10U_1_if_4_if_and_tmp_1 = (fsm_output[1]) & (~ (chn_inp_in_crt_sva_7_739_736_1[1]));
  assign FpAdd_6U_10U_1_if_4_if_and_tmp_2 = (fsm_output[1]) & (~ (chn_inp_in_crt_sva_7_739_736_1[2]));
  assign FpAdd_6U_10U_1_if_4_if_and_tmp_3 = (fsm_output[1]) & (~ (chn_inp_in_crt_sva_7_739_736_1[3]));
  assign FpAdd_6U_10U_b_right_shift_qif_and_tmp = (fsm_output[1]) & FpAdd_6U_10U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0;
  assign FpAdd_6U_10U_b_right_shift_qif_and_tmp_1 = (fsm_output[1]) & FpAdd_6U_10U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0;
  assign FpAdd_6U_10U_b_right_shift_qif_and_tmp_2 = (fsm_output[1]) & FpAdd_6U_10U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0;
  assign FpAdd_6U_10U_b_right_shift_qif_and_tmp_3 = (fsm_output[1]) & FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_1_mx0w0;
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_and_tmp = (fsm_output[1]) & (chn_inp_in_rsci_d_mxwt[736]);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_if_1_if_and_tmp_1 = (fsm_output[1]) & (chn_inp_in_rsci_d_mxwt[738]);
  assign or_tmp_4811 = FpMul_6U_10U_2_lor_6_lpi_1_dfm_st_3 | IsNaN_6U_10U_7_land_1_lpi_1_dfm_5;
  assign or_tmp_4815 = (fsm_output[0]) | (~ or_4340_cse);
  assign mux_tmp = MUX_s_1_2_2(or_tmp_4815, (fsm_output[0]), or_6231_cse);
  assign not_tmp_3015 = ~((cfg_precision_1_sva_st_90[1]) | (~ (fsm_output[0])));
  assign or_tmp_4829 = (cfg_precision_1_sva_st_80[0]) | (~((cfg_precision_1_sva_st_80[1])
      & (chn_inp_in_crt_sva_3_739_736_1[1])));
  assign or_tmp_4830 = (fsm_output[0]) | (~ or_tmp_4829);
  assign mux_tmp_2075 = MUX_s_1_2_2(or_tmp_4830, (fsm_output[0]), or_6230_cse);
  assign or_tmp_4831 = FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_3 | IsNaN_6U_10U_7_land_2_lpi_1_dfm_5;
  assign or_tmp_4843 = FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_3 | IsNaN_6U_10U_7_land_3_lpi_1_dfm_5;
  assign or_tmp_4845 = (cfg_precision_1_sva_st_80[0]) | (~((cfg_precision_1_sva_st_80[1])
      & (chn_inp_in_crt_sva_3_739_736_1[2])));
  assign or_tmp_4846 = (fsm_output[0]) | (~ or_tmp_4845);
  assign mux_tmp_2091 = MUX_s_1_2_2(or_tmp_4846, (fsm_output[0]), or_6229_cse);
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_rsci_iswt0 <= 1'b0;
      chn_inp_out_rsci_iswt0 <= 1'b0;
    end
    else if ( core_wen ) begin
      chn_inp_in_rsci_iswt0 <= ~((~ main_stage_en_1) & (fsm_output[1]));
      chn_inp_out_rsci_iswt0 <= and_dcpl_96;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_rsci_ld_core_psct <= 1'b0;
    end
    else if ( core_wen & chn_inp_in_rsci_ld_core_psct_mx0c0 ) begin
      chn_inp_in_rsci_ld_core_psct <= chn_inp_in_rsci_ld_core_psct_mx0c0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_out_rsci_d_26_23 <= 4'b0;
      chn_inp_out_rsci_d_27 <= 1'b0;
      chn_inp_out_rsci_d_58_55 <= 4'b0;
      chn_inp_out_rsci_d_59 <= 1'b0;
      chn_inp_out_rsci_d_90_87 <= 4'b0;
      chn_inp_out_rsci_d_91 <= 1'b0;
      chn_inp_out_rsci_d_122_119 <= 4'b0;
      chn_inp_out_rsci_d_123 <= 1'b0;
      chn_inp_out_rsci_d_9_1 <= 9'b0;
      chn_inp_out_rsci_d_12_10 <= 3'b0;
      chn_inp_out_rsci_d_22_13 <= 10'b0;
      chn_inp_out_rsci_d_30_28 <= 3'b0;
      chn_inp_out_rsci_d_31 <= 1'b0;
      chn_inp_out_rsci_d_41_33 <= 9'b0;
      chn_inp_out_rsci_d_44_42 <= 3'b0;
      chn_inp_out_rsci_d_54_45 <= 10'b0;
      chn_inp_out_rsci_d_62_60 <= 3'b0;
      chn_inp_out_rsci_d_63 <= 1'b0;
      chn_inp_out_rsci_d_73_65 <= 9'b0;
      chn_inp_out_rsci_d_76_74 <= 3'b0;
      chn_inp_out_rsci_d_86_77 <= 10'b0;
      chn_inp_out_rsci_d_94_92 <= 3'b0;
      chn_inp_out_rsci_d_95 <= 1'b0;
      chn_inp_out_rsci_d_105_97 <= 9'b0;
      chn_inp_out_rsci_d_108_106 <= 3'b0;
      chn_inp_out_rsci_d_118_109 <= 10'b0;
      chn_inp_out_rsci_d_126_124 <= 3'b0;
      chn_inp_out_rsci_d_127 <= 1'b0;
    end
    else if ( chn_inp_out_and_cse ) begin
      chn_inp_out_rsci_d_26_23 <= MUX1HOT_v_4_4_2(FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_8_3_0_1,
          (signext_4_1(reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_10_17_1_itm[7])),
          (FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_4_nl),
          (IntSaturation_51U_32U_o_1_lpi_1_dfm_12_30_0_1[26:23]), {inp_lookup_and_8_m1c
          , inp_lookup_asn_106 , inp_lookup_and_10_m1c , inp_lookup_asn_110});
      chn_inp_out_rsci_d_27 <= MUX1HOT_s_1_4_2(FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_8_4_1,
          (reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_10_17_1_itm[7]),
          (FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_20_nl),
          (IntSaturation_51U_32U_o_1_lpi_1_dfm_12_30_0_1[27]), {inp_lookup_and_8_m1c
          , inp_lookup_asn_106 , inp_lookup_and_10_m1c , inp_lookup_asn_110});
      chn_inp_out_rsci_d_58_55 <= MUX1HOT_v_4_4_2(FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_8_3_0_1,
          (signext_4_1(reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_10_17_1_itm[7])),
          (FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_9_nl),
          (IntSaturation_51U_32U_o_2_lpi_1_dfm_12_30_0_1[26:23]), {inp_lookup_and_28_m1c
          , inp_lookup_asn_122 , inp_lookup_and_30_m1c , inp_lookup_asn_126});
      chn_inp_out_rsci_d_59 <= MUX1HOT_s_1_4_2(FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_8_4_1,
          (reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_10_17_1_itm[7]),
          (FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_21_nl),
          (IntSaturation_51U_32U_o_2_lpi_1_dfm_12_30_0_1[27]), {inp_lookup_and_28_m1c
          , inp_lookup_asn_122 , inp_lookup_and_30_m1c , inp_lookup_asn_126});
      chn_inp_out_rsci_d_90_87 <= MUX1HOT_v_4_4_2(FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_8_3_0_1,
          (signext_4_1(reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_10_17_1_itm[7])),
          (FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_14_nl),
          (IntSaturation_51U_32U_o_3_lpi_1_dfm_12_30_0_1[26:23]), {inp_lookup_and_48_m1c
          , inp_lookup_asn_114 , inp_lookup_and_50_m1c , inp_lookup_asn_118});
      chn_inp_out_rsci_d_91 <= MUX1HOT_s_1_4_2(FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_8_4_1,
          (reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_10_17_1_itm[7]),
          (FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_22_nl),
          (IntSaturation_51U_32U_o_3_lpi_1_dfm_12_30_0_1[27]), {inp_lookup_and_48_m1c
          , inp_lookup_asn_114 , inp_lookup_and_50_m1c , inp_lookup_asn_118});
      chn_inp_out_rsci_d_122_119 <= MUX1HOT_v_4_4_2(FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_8_3_0_1,
          (signext_4_1(reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_10_17_1_itm[7])),
          (FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_19_nl),
          (IntSaturation_51U_32U_o_lpi_1_dfm_12_30_0_1[26:23]), {inp_lookup_and_68_m1c
          , inp_lookup_asn_98 , inp_lookup_and_70_m1c , inp_lookup_asn_102});
      chn_inp_out_rsci_d_123 <= MUX1HOT_s_1_4_2(FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_8_4_1,
          (reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_10_17_1_itm[7]),
          (FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_23_nl),
          (IntSaturation_51U_32U_o_lpi_1_dfm_12_30_0_1[27]), {inp_lookup_and_68_m1c
          , inp_lookup_asn_98 , inp_lookup_and_70_m1c , inp_lookup_asn_102});
      chn_inp_out_rsci_d_9_1 <= MUX1HOT_v_9_3_2((FpExpoWidthInc_6U_8U_23U_0U_1U_o_mant_9_0_1_lpi_1_dfm_2_mx0[9:1]),
          (IntSaturation_51U_32U_o_1_lpi_1_dfm_12_30_0_1[9:1]), reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_10_17_1_1_itm,
          {(nor_1802_nl) , inp_lookup_asn_110 , or_5836_tmp});
      chn_inp_out_rsci_d_12_10 <= MUX1HOT_v_3_4_2(({{2{FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_4_itm_8}},
          FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_4_itm_8}),
          (reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_10_17_1_itm[2:0]),
          (signext_3_1(FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_4_nl)),
          (IntSaturation_51U_32U_o_1_lpi_1_dfm_12_30_0_1[12:10]), {inp_lookup_and_8_m1c
          , inp_lookup_asn_106 , inp_lookup_and_10_m1c , inp_lookup_asn_110});
      chn_inp_out_rsci_d_22_13 <= MUX1HOT_v_10_5_2(FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_1_lpi_1_dfm_12,
          (signext_10_5(reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_10_17_1_itm[7:3])),
          ({{9{IsInf_6U_23U_land_1_lpi_1_dfm_mx0w0}}, IsInf_6U_23U_land_1_lpi_1_dfm_mx0w0}),
          (IntSaturation_51U_32U_o_1_lpi_1_dfm_12_30_0_1[22:13]), FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_22_13_1_lpi_1_dfm,
          {(inp_lookup_or_nl) , inp_lookup_asn_106 , (inp_lookup_and_82_nl) , inp_lookup_asn_110
          , and_3545_tmp});
      chn_inp_out_rsci_d_30_28 <= MUX1HOT_v_3_4_2(FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_1_lpi_1_dfm_12,
          (signext_3_1(reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_10_17_1_itm[7])),
          (FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_3_nl),
          (IntSaturation_51U_32U_o_1_lpi_1_dfm_12_30_0_1[30:28]), {inp_lookup_and_8_m1c
          , inp_lookup_asn_106 , inp_lookup_and_10_m1c , inp_lookup_asn_110});
      chn_inp_out_rsci_d_31 <= inp_lookup_mux_259_itm_4;
      chn_inp_out_rsci_d_41_33 <= MUX1HOT_v_9_3_2((FpExpoWidthInc_6U_8U_23U_0U_1U_o_mant_9_0_2_lpi_1_dfm_2_mx0[9:1]),
          (IntSaturation_51U_32U_o_2_lpi_1_dfm_12_30_0_1[9:1]), reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_10_17_1_1_itm,
          {(nor_1803_nl) , inp_lookup_asn_126 , or_5838_tmp});
      chn_inp_out_rsci_d_44_42 <= MUX1HOT_v_3_4_2(({{2{FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_9_itm_8}},
          FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_9_itm_8}),
          (reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_10_17_1_itm[2:0]),
          (signext_3_1(FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_9_nl)),
          (IntSaturation_51U_32U_o_2_lpi_1_dfm_12_30_0_1[12:10]), {inp_lookup_and_28_m1c
          , inp_lookup_asn_122 , inp_lookup_and_30_m1c , inp_lookup_asn_126});
      chn_inp_out_rsci_d_54_45 <= MUX1HOT_v_10_5_2(FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_2_lpi_1_dfm_12,
          (signext_10_5(reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_10_17_1_itm[7:3])),
          ({{9{IsInf_6U_23U_land_2_lpi_1_dfm_mx0w0}}, IsInf_6U_23U_land_2_lpi_1_dfm_mx0w0}),
          (IntSaturation_51U_32U_o_2_lpi_1_dfm_12_30_0_1[22:13]), FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_22_13_2_lpi_1_dfm,
          {(inp_lookup_or_1_nl) , inp_lookup_asn_122 , (inp_lookup_and_86_nl) , inp_lookup_asn_126
          , and_3546_tmp});
      chn_inp_out_rsci_d_62_60 <= MUX1HOT_v_3_4_2(FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_2_lpi_1_dfm_12,
          (signext_3_1(reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_10_17_1_itm[7])),
          (FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_8_nl),
          (IntSaturation_51U_32U_o_2_lpi_1_dfm_12_30_0_1[30:28]), {inp_lookup_and_28_m1c
          , inp_lookup_asn_122 , inp_lookup_and_30_m1c , inp_lookup_asn_126});
      chn_inp_out_rsci_d_63 <= inp_lookup_mux_525_itm_4;
      chn_inp_out_rsci_d_73_65 <= MUX1HOT_v_9_3_2((FpExpoWidthInc_6U_8U_23U_0U_1U_o_mant_9_0_3_lpi_1_dfm_2_mx0[9:1]),
          (IntSaturation_51U_32U_o_3_lpi_1_dfm_12_30_0_1[9:1]), reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_10_17_1_1_itm,
          {(nor_1804_nl) , inp_lookup_asn_118 , or_5840_tmp});
      chn_inp_out_rsci_d_76_74 <= MUX1HOT_v_3_4_2(({{2{FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_14_itm_8}},
          FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_14_itm_8}),
          (reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_10_17_1_itm[2:0]),
          (signext_3_1(FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_14_nl)),
          (IntSaturation_51U_32U_o_3_lpi_1_dfm_12_30_0_1[12:10]), {inp_lookup_and_48_m1c
          , inp_lookup_asn_114 , inp_lookup_and_50_m1c , inp_lookup_asn_118});
      chn_inp_out_rsci_d_86_77 <= MUX1HOT_v_10_5_2(FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_3_lpi_1_dfm_12,
          (signext_10_5(reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_10_17_1_itm[7:3])),
          ({{9{IsInf_6U_23U_land_3_lpi_1_dfm_mx0w0}}, IsInf_6U_23U_land_3_lpi_1_dfm_mx0w0}),
          (IntSaturation_51U_32U_o_3_lpi_1_dfm_12_30_0_1[22:13]), FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_22_13_3_lpi_1_dfm,
          {(inp_lookup_or_2_nl) , inp_lookup_asn_114 , (inp_lookup_and_90_nl) , inp_lookup_asn_118
          , and_3547_tmp});
      chn_inp_out_rsci_d_94_92 <= MUX1HOT_v_3_4_2(FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_3_lpi_1_dfm_12,
          (signext_3_1(reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_10_17_1_itm[7])),
          (FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_13_nl),
          (IntSaturation_51U_32U_o_3_lpi_1_dfm_12_30_0_1[30:28]), {inp_lookup_and_48_m1c
          , inp_lookup_asn_114 , inp_lookup_and_50_m1c , inp_lookup_asn_118});
      chn_inp_out_rsci_d_95 <= inp_lookup_mux_791_itm_4;
      chn_inp_out_rsci_d_105_97 <= MUX1HOT_v_9_3_2((FpExpoWidthInc_6U_8U_23U_0U_1U_o_mant_9_0_lpi_1_dfm_2_mx0[9:1]),
          (IntSaturation_51U_32U_o_lpi_1_dfm_12_30_0_1[9:1]), reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_10_17_1_1_itm,
          {(nor_1805_nl) , inp_lookup_asn_102 , or_5842_tmp});
      chn_inp_out_rsci_d_108_106 <= MUX1HOT_v_3_4_2(({{2{FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_19_itm_8}},
          FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_19_itm_8}),
          (reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_10_17_1_itm[2:0]),
          (signext_3_1(FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_19_nl)),
          (IntSaturation_51U_32U_o_lpi_1_dfm_12_30_0_1[12:10]), {inp_lookup_and_68_m1c
          , inp_lookup_asn_98 , inp_lookup_and_70_m1c , inp_lookup_asn_102});
      chn_inp_out_rsci_d_118_109 <= MUX1HOT_v_10_5_2(FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_lpi_1_dfm_12,
          (signext_10_5(reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_10_17_1_itm[7:3])),
          ({{9{IsInf_6U_23U_land_lpi_1_dfm_mx0w0}}, IsInf_6U_23U_land_lpi_1_dfm_mx0w0}),
          (IntSaturation_51U_32U_o_lpi_1_dfm_12_30_0_1[22:13]), FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_22_13_lpi_1_dfm,
          {(inp_lookup_or_3_nl) , inp_lookup_asn_98 , (inp_lookup_and_94_nl) , inp_lookup_asn_102
          , and_3548_tmp});
      chn_inp_out_rsci_d_126_124 <= MUX1HOT_v_3_4_2(FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_lpi_1_dfm_12,
          (signext_3_1(reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_10_17_1_itm[7])),
          (FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_18_nl),
          (IntSaturation_51U_32U_o_lpi_1_dfm_12_30_0_1[30:28]), {inp_lookup_and_68_m1c
          , inp_lookup_asn_98 , inp_lookup_and_70_m1c , inp_lookup_asn_102});
      chn_inp_out_rsci_d_127 <= inp_lookup_mux_1057_itm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_out_rsci_d_0 <= 1'b0;
    end
    else if ( core_wen & ((main_stage_v_12 & (chn_inp_in_crt_sva_12_739_736_1[0])
        & or_11_cse) | chn_inp_out_rsci_d_0_mx0c1) ) begin
      chn_inp_out_rsci_d_0 <= MUX_s_1_2_2((inp_lookup_if_mux_600_nl), inp_lookup_else_mux_122_itm_8,
          chn_inp_out_rsci_d_0_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_out_rsci_d_32 <= 1'b0;
    end
    else if ( core_wen & ((main_stage_v_12 & (chn_inp_in_crt_sva_12_739_736_1[1])
        & or_11_cse) | chn_inp_out_rsci_d_32_mx0c1) ) begin
      chn_inp_out_rsci_d_32 <= MUX_s_1_2_2((inp_lookup_if_mux_601_nl), inp_lookup_else_mux_245_itm_8,
          chn_inp_out_rsci_d_32_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_out_rsci_d_64 <= 1'b0;
    end
    else if ( core_wen & ((main_stage_v_12 & (chn_inp_in_crt_sva_12_739_736_1[2])
        & or_11_cse) | chn_inp_out_rsci_d_64_mx0c1) ) begin
      chn_inp_out_rsci_d_64 <= MUX_s_1_2_2((inp_lookup_if_mux_602_nl), inp_lookup_else_mux_368_itm_8,
          chn_inp_out_rsci_d_64_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_out_rsci_d_96 <= 1'b0;
    end
    else if ( core_wen & ((main_stage_v_12 & (chn_inp_in_crt_sva_12_739_736_1[3])
        & or_11_cse) | chn_inp_out_rsci_d_96_mx0c1) ) begin
      chn_inp_out_rsci_d_96 <= MUX_s_1_2_2((inp_lookup_if_mux_603_nl), inp_lookup_else_mux_491_itm_8,
          chn_inp_out_rsci_d_96_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_out_rsci_ld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_96 | and_dcpl_98) ) begin
      reg_chn_inp_out_rsci_ld_core_psct_cse <= ~ and_dcpl_98;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_1 <= 1'b0;
    end
    else if ( core_wen & (or_tmp_4339 | main_stage_v_1_mx0c1) ) begin
      main_stage_v_1 <= ~ main_stage_v_1_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_3 <= 1'b0;
      inp_lookup_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3 <=
          1'b0;
      IsNaN_8U_23U_2_land_1_lpi_1_dfm_st_6 <= 1'b0;
      inp_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_5 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_aelse_and_cse ) begin
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_3 <= ~(IsNaN_8U_23U_nor_tmp | (chn_inp_in_rsci_d_mxwt[510:503]!=8'b11111111));
      inp_lookup_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3 <=
          ~((chn_inp_in_rsci_d_mxwt[511]) ^ (chn_inp_in_rsci_d_mxwt[639]));
      IsNaN_8U_23U_2_land_1_lpi_1_dfm_st_6 <= ~((~((chn_inp_in_rsci_d_mxwt[22:0]!=23'b00000000000000000000000)))
          | (chn_inp_in_rsci_d_mxwt[30:23]!=8'b11111111));
      inp_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_5 <= (chn_inp_in_rsci_d_mxwt[30:0]!=31'b0000000000000000000000000000000);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_st_2 <= 1'b0;
      IsZero_6U_10U_7_IsZero_6U_10U_7_and_itm_2 <= 1'b0;
      FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_5 <= 1'b0;
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_itm_7 <= 1'b0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_13 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_is_a_greater_oelse_and_cse ) begin
      FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_st_2 <= MUX_s_1_2_2(FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0,
          inp_lookup_else_if_unequal_tmp_mx0w1, and_dcpl_105);
      IsZero_6U_10U_7_IsZero_6U_10U_7_and_itm_2 <= MUX_s_1_2_2((IsZero_6U_10U_7_IsZero_6U_10U_7_and_nl),
          (inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_nl), and_dcpl_38);
      FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0,
          (chn_inp_in_rsci_d_mxwt[347]), and_dcpl_105);
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_itm_7 <= MUX_s_1_2_2((IsZero_6U_10U_1_IsZero_6U_10U_1_and_nl),
          (IsZero_6U_10U_5_IsZero_6U_10U_5_and_nl), and_dcpl_105);
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_13 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_1_lpi_1_dfm_mx0w0,
          inp_lookup_else_if_unequal_tmp_mx0w1, and_dcpl_105);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_35U_leading_sign_35_0_rtn_1_sva_2 <= 6'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_80_nl) ) begin
      IntLeadZero_35U_leading_sign_35_0_rtn_1_sva_2 <= libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_35U_1_leading_sign_35_0_rtn_1_sva_2 <= 6'b0;
      inp_lookup_1_FpMantRNE_36U_11U_1_else_and_svs_2 <= 1'b0;
    end
    else if ( IntLeadZero_35U_1_leading_sign_35_0_rtn_and_4_cse ) begin
      IntLeadZero_35U_1_leading_sign_35_0_rtn_1_sva_2 <= MUX_v_6_2_2(libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_12,
          IntLeadZero_35U_1_leading_sign_35_0_rtn_1_sva, and_dcpl_141);
      inp_lookup_1_FpMantRNE_36U_11U_1_else_and_svs_2 <= MUX_s_1_2_2(inp_lookup_1_FpMantRNE_36U_11U_1_else_and_tmp,
          inp_lookup_1_FpMantRNE_36U_11U_1_else_and_svs, and_dcpl_141);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_6_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_6_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_9 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_12_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_6_1_1 <= MUX_s_1_2_2((chn_inp_in_rsci_d_mxwt[346]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_3_1, and_dcpl_145);
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_6_0_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_3_0_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_3_0, and_dcpl_145);
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_3, and_dcpl_145);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFractionToFloat_35U_6U_10U_1_o_mant_1_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & ((and_dcpl_106 & (~ inp_lookup_1_FpMantRNE_36U_11U_1_else_and_tmp))
        | FpFractionToFloat_35U_6U_10U_1_o_mant_1_lpi_1_dfm_6_mx0c1) ) begin
      FpFractionToFloat_35U_6U_10U_1_o_mant_1_lpi_1_dfm_6 <= MUX1HOT_v_10_3_2((FpFractionToFloat_35U_6U_10U_1_if_else_else_FpFractionToFloat_35U_6U_10U_1_if_else_else_and_nl),
          (FpMantRNE_36U_11U_1_else_ac_int_cctor_2_sva_mx0w0[10:1]), reg_FpMantRNE_36U_11U_1_else_ac_int_cctor_2_tmp,
          {(~ FpFractionToFloat_35U_6U_10U_1_o_mant_1_lpi_1_dfm_6_mx0c1) , (FpFractionToFloat_35U_6U_10U_1_o_mant_and_nl)
          , (FpFractionToFloat_35U_6U_10U_1_o_mant_and_10_nl)});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFractionToFloat_35U_6U_10U_1_if_else_else_if_slc_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_5_mdf_1_sva_2
          <= 1'b0;
      inp_lookup_1_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_3 <= 35'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_6_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_6_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_8 <= 4'b0;
    end
    else if ( FpFractionToFloat_35U_6U_10U_1_if_else_else_and_cse ) begin
      FpFractionToFloat_35U_6U_10U_1_if_else_else_if_slc_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_5_mdf_1_sva_2
          <= inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_itm_5;
      inp_lookup_1_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_3 <= chn_inp_in_rsci_d_mxwt[162:128];
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_6_1_1 <= chn_inp_in_rsci_d_mxwt[282];
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_6_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_3_0_mx0w0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_8 <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_st_90 <= 2'b0;
      chn_inp_in_crt_sva_1_739_395_1 <= 345'b0;
      chn_inp_in_crt_sva_1_127_0_1 <= 128'b0;
      chn_inp_in_crt_sva_1_331_268_1 <= 64'b0;
      IsNaN_6U_10U_2_land_lpi_1_dfm_15 <= 1'b0;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_15 <= 1'b0;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_15 <= 1'b0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_15 <= 1'b0;
    end
    else if ( cfg_precision_and_cse ) begin
      cfg_precision_1_sva_st_90 <= cfg_precision_rsci_d;
      chn_inp_in_crt_sva_1_739_395_1 <= chn_inp_in_rsci_d_mxwt[739:395];
      chn_inp_in_crt_sva_1_127_0_1 <= chn_inp_in_rsci_d_mxwt[127:0];
      chn_inp_in_crt_sva_1_331_268_1 <= chn_inp_in_rsci_d_mxwt[331:268];
      IsNaN_6U_10U_2_land_lpi_1_dfm_15 <= IsNaN_6U_10U_2_land_lpi_1_dfm_mx0w0;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_15 <= IsNaN_6U_10U_2_land_3_lpi_1_dfm_mx0w0;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_15 <= IsNaN_6U_10U_2_land_2_lpi_1_dfm_mx0w0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_15 <= IsNaN_6U_10U_2_land_1_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_st_2 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_6_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_6_0_1 <= 1'b0;
      IsZero_6U_10U_5_IsZero_6U_10U_5_and_1_itm_2 <= 1'b0;
      FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_13 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_is_a_greater_oelse_and_1_cse ) begin
      FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_st_2 <= MUX_s_1_2_2(FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0,
          inp_lookup_else_if_unequal_tmp_1_mx0w1, and_dcpl_176);
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_6_1_1 <= MUX_s_1_2_2((chn_inp_in_rsci_d_mxwt[298]),
          inp_lookup_2_IsZero_6U_10U_5_IsZero_6U_10U_5_nor_mx0w1, and_dcpl_49);
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_6_0_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_3_0_mx0w0,
          (inp_lookup_2_IsZero_6U_10U_1_IsZero_6U_10U_1_nor_nl), and_dcpl_49);
      IsZero_6U_10U_5_IsZero_6U_10U_5_and_1_itm_2 <= MUX_s_1_2_2((IsZero_6U_10U_5_IsZero_6U_10U_5_and_1_nl),
          (inp_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_nl), and_dcpl_49);
      FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0,
          (chn_inp_in_rsci_d_mxwt[363]), and_dcpl_176);
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_13 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_2_lpi_1_dfm_mx0w0,
          inp_lookup_else_if_unequal_tmp_1_mx0w1, and_dcpl_176);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_35U_leading_sign_35_0_rtn_2_sva_2 <= 6'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_86_nl) ) begin
      IntLeadZero_35U_leading_sign_35_0_rtn_2_sva_2 <= libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_35U_1_leading_sign_35_0_rtn_2_sva_2 <= 6'b0;
      inp_lookup_2_FpMantRNE_36U_11U_1_else_and_svs_2 <= 1'b0;
    end
    else if ( IntLeadZero_35U_1_leading_sign_35_0_rtn_and_5_cse ) begin
      IntLeadZero_35U_1_leading_sign_35_0_rtn_2_sva_2 <= MUX_v_6_2_2(libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_13,
          IntLeadZero_35U_1_leading_sign_35_0_rtn_2_sva, and_dcpl_212);
      inp_lookup_2_FpMantRNE_36U_11U_1_else_and_svs_2 <= MUX_s_1_2_2(inp_lookup_2_FpMantRNE_36U_11U_1_else_and_tmp,
          inp_lookup_2_FpMantRNE_36U_11U_1_else_and_svs, and_dcpl_212);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_6_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_6_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_9 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_15_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_6_1_1 <= MUX_s_1_2_2((chn_inp_in_rsci_d_mxwt[362]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_3_1, and_dcpl_215);
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_6_0_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_3_0_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_3_0, and_dcpl_215);
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_3, and_dcpl_215);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_6U_10U_7_IsZero_6U_10U_7_and_1_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_is_a_greater_oelse_FpAdd_8U_23U_is_a_greater_oelse_or_19_cse
        & (~ (mux_92_nl)) ) begin
      IsZero_6U_10U_7_IsZero_6U_10U_7_and_1_itm_2 <= MUX_s_1_2_2((IsZero_6U_10U_7_IsZero_6U_10U_7_and_1_nl),
          (inp_lookup_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_nl), and_dcpl_49);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFractionToFloat_35U_6U_10U_1_o_mant_2_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & ((and_dcpl_177 & (~ inp_lookup_2_FpMantRNE_36U_11U_1_else_and_tmp))
        | FpFractionToFloat_35U_6U_10U_1_o_mant_2_lpi_1_dfm_6_mx0c1) ) begin
      FpFractionToFloat_35U_6U_10U_1_o_mant_2_lpi_1_dfm_6 <= MUX1HOT_v_10_3_2((FpFractionToFloat_35U_6U_10U_1_if_else_else_FpFractionToFloat_35U_6U_10U_1_if_else_else_and_1_nl),
          (FpMantRNE_36U_11U_1_else_ac_int_cctor_3_sva_mx0w0[10:1]), reg_FpMantRNE_36U_11U_1_else_ac_int_cctor_3_tmp,
          {(~ FpFractionToFloat_35U_6U_10U_1_o_mant_2_lpi_1_dfm_6_mx0c1) , (FpFractionToFloat_35U_6U_10U_1_o_mant_and_8_nl)
          , (FpFractionToFloat_35U_6U_10U_1_o_mant_and_9_nl)});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFractionToFloat_35U_6U_10U_1_if_else_else_if_slc_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_5_mdf_2_sva_2
          <= 1'b0;
      inp_lookup_2_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_3 <= 35'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_8 <= 4'b0;
    end
    else if ( FpFractionToFloat_35U_6U_10U_1_if_else_else_and_1_cse ) begin
      FpFractionToFloat_35U_6U_10U_1_if_else_else_if_slc_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_5_mdf_2_sva_2
          <= inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_itm_5;
      inp_lookup_2_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_3 <= chn_inp_in_rsci_d_mxwt[197:163];
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_8 <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_st_2 <= 1'b0;
      IsZero_6U_10U_7_IsZero_6U_10U_7_and_2_itm_2 <= 1'b0;
      FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_5 <= 1'b0;
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_itm_7 <= 1'b0;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_13 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_is_a_greater_oelse_and_2_cse ) begin
      FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_st_2 <= MUX_s_1_2_2(FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0,
          or_79_cse, and_dcpl_246);
      IsZero_6U_10U_7_IsZero_6U_10U_7_and_2_itm_2 <= MUX_s_1_2_2((IsZero_6U_10U_7_IsZero_6U_10U_7_and_2_nl),
          (inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_nl), and_dcpl_57);
      FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0,
          (chn_inp_in_rsci_d_mxwt[379]), and_dcpl_246);
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_itm_7 <= MUX_s_1_2_2((IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_nl),
          (IsZero_6U_10U_5_IsZero_6U_10U_5_and_2_nl), and_dcpl_246);
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_13 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_3_lpi_1_dfm_mx0w0,
          or_79_cse, and_dcpl_246);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_35U_leading_sign_35_0_rtn_3_sva_2 <= 6'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_94_nl) ) begin
      IntLeadZero_35U_leading_sign_35_0_rtn_3_sva_2 <= libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_35U_1_leading_sign_35_0_rtn_3_sva_2 <= 6'b0;
      inp_lookup_3_FpMantRNE_36U_11U_1_else_and_svs_2 <= 1'b0;
    end
    else if ( IntLeadZero_35U_1_leading_sign_35_0_rtn_and_6_cse ) begin
      IntLeadZero_35U_1_leading_sign_35_0_rtn_3_sva_2 <= MUX_v_6_2_2(libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_14,
          IntLeadZero_35U_1_leading_sign_35_0_rtn_3_sva, and_dcpl_282);
      inp_lookup_3_FpMantRNE_36U_11U_1_else_and_svs_2 <= MUX_s_1_2_2(inp_lookup_3_FpMantRNE_36U_11U_1_else_and_tmp,
          inp_lookup_3_FpMantRNE_36U_11U_1_else_and_svs, and_dcpl_282);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_6_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_6_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_3_lpi_1_dfm_9 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_18_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_6_1_1 <= MUX_s_1_2_2((chn_inp_in_rsci_d_mxwt[378]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_3_1, and_dcpl_285);
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_6_0_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_3_0_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_3_0, and_dcpl_285);
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_3_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_3_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_3_lpi_1_dfm_3, and_dcpl_285);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFractionToFloat_35U_6U_10U_1_o_mant_3_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & ((and_dcpl_247 & (~ inp_lookup_3_FpMantRNE_36U_11U_1_else_and_tmp))
        | FpFractionToFloat_35U_6U_10U_1_o_mant_3_lpi_1_dfm_6_mx0c1) ) begin
      FpFractionToFloat_35U_6U_10U_1_o_mant_3_lpi_1_dfm_6 <= MUX1HOT_v_10_3_2((FpFractionToFloat_35U_6U_10U_1_if_else_else_FpFractionToFloat_35U_6U_10U_1_if_else_else_and_2_nl),
          (FpMantRNE_36U_11U_1_else_ac_int_cctor_4_sva_mx0w0[10:1]), reg_FpMantRNE_36U_11U_1_else_ac_int_cctor_4_tmp,
          {(~ FpFractionToFloat_35U_6U_10U_1_o_mant_3_lpi_1_dfm_6_mx0c1) , (FpFractionToFloat_35U_6U_10U_1_o_mant_and_6_nl)
          , (FpFractionToFloat_35U_6U_10U_1_o_mant_and_7_nl)});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFractionToFloat_35U_6U_10U_1_if_else_else_if_slc_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_5_mdf_3_sva_2
          <= 1'b0;
      inp_lookup_3_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_3 <= 35'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_6_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_6_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_8 <= 4'b0;
    end
    else if ( FpFractionToFloat_35U_6U_10U_1_if_else_else_and_2_cse ) begin
      FpFractionToFloat_35U_6U_10U_1_if_else_else_if_slc_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_5_mdf_3_sva_2
          <= inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_itm_5;
      inp_lookup_3_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_3 <= chn_inp_in_rsci_d_mxwt[232:198];
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_6_1_1 <= chn_inp_in_rsci_d_mxwt[314];
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_6_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_3_0_mx0w0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_8 <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_6_0_1 <= 1'b0;
      IsZero_6U_10U_5_IsZero_6U_10U_5_and_3_itm_2 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_is_a_greater_oelse_and_3_cse ) begin
      FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2 <= MUX_s_1_2_2((FpAdd_8U_23U_is_a_greater_FpAdd_8U_23U_is_a_greater_or_3_nl),
          inp_lookup_else_if_unequal_tmp_3_mx0w1, and_dcpl_316);
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_6_0_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_3_0_mx0w0,
          inp_lookup_4_IsZero_6U_10U_5_IsZero_6U_10U_5_nor_mx0w1, and_dcpl_65);
      IsZero_6U_10U_5_IsZero_6U_10U_5_and_3_itm_2 <= MUX_s_1_2_2((IsZero_6U_10U_5_IsZero_6U_10U_5_and_3_nl),
          (inp_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_nl), and_dcpl_65);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_35U_leading_sign_35_0_rtn_sva_2 <= 6'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_99_nl) ) begin
      IntLeadZero_35U_leading_sign_35_0_rtn_sva_2 <= libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_11;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_35U_1_leading_sign_35_0_rtn_sva_2 <= 6'b0;
      inp_lookup_4_FpMantRNE_36U_11U_1_else_and_svs_2 <= 1'b0;
    end
    else if ( IntLeadZero_35U_1_leading_sign_35_0_rtn_and_7_cse ) begin
      IntLeadZero_35U_1_leading_sign_35_0_rtn_sva_2 <= MUX_v_6_2_2(libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_15,
          IntLeadZero_35U_1_leading_sign_35_0_rtn_sva, and_dcpl_352);
      inp_lookup_4_FpMantRNE_36U_11U_1_else_and_svs_2 <= MUX_s_1_2_2(inp_lookup_4_FpMantRNE_36U_11U_1_else_and_tmp,
          inp_lookup_4_FpMantRNE_36U_11U_1_else_and_svs, and_dcpl_352);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_6_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_6_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_9 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_21_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_6_1_1 <= MUX_s_1_2_2((chn_inp_in_rsci_d_mxwt[394]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_3_1, and_dcpl_355);
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_6_0_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_3_0_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_3_0, and_dcpl_355);
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_9 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_3, and_dcpl_355);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_6U_10U_7_IsZero_6U_10U_7_and_3_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_is_a_greater_oelse_FpAdd_8U_23U_is_a_greater_oelse_or_17_cse
        & (~ (mux_105_nl)) ) begin
      IsZero_6U_10U_7_IsZero_6U_10U_7_and_3_itm_2 <= MUX_s_1_2_2((IsZero_6U_10U_7_IsZero_6U_10U_7_and_3_nl),
          (inp_lookup_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_nl), and_dcpl_65);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFractionToFloat_35U_6U_10U_1_o_mant_lpi_1_dfm_6 <= 10'b0;
    end
    else if ( core_wen & ((and_dcpl_317 & (~ inp_lookup_4_FpMantRNE_36U_11U_1_else_and_tmp))
        | FpFractionToFloat_35U_6U_10U_1_o_mant_lpi_1_dfm_6_mx0c1) ) begin
      FpFractionToFloat_35U_6U_10U_1_o_mant_lpi_1_dfm_6 <= MUX1HOT_v_10_3_2((FpFractionToFloat_35U_6U_10U_1_if_else_else_FpFractionToFloat_35U_6U_10U_1_if_else_else_and_3_nl),
          (FpMantRNE_36U_11U_1_else_ac_int_cctor_sva_mx0w0[10:1]), reg_FpMantRNE_36U_11U_1_else_ac_int_cctor_tmp,
          {(~ FpFractionToFloat_35U_6U_10U_1_o_mant_lpi_1_dfm_6_mx0c1) , (FpFractionToFloat_35U_6U_10U_1_o_mant_and_4_nl)
          , (FpFractionToFloat_35U_6U_10U_1_o_mant_and_5_nl)});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFractionToFloat_35U_6U_10U_1_if_else_else_if_slc_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_5_mdf_sva_2
          <= 1'b0;
      inp_lookup_4_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_3 <= 35'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_6_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_8 <= 4'b0;
    end
    else if ( FpFractionToFloat_35U_6U_10U_1_if_else_else_and_3_cse ) begin
      FpFractionToFloat_35U_6U_10U_1_if_else_else_if_slc_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_5_mdf_sva_2
          <= inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_itm_5;
      inp_lookup_4_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_3 <= chn_inp_in_rsci_d_mxwt[267:233];
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_6_1_1 <= chn_inp_in_rsci_d_mxwt[330];
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_8 <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_2 <= 1'b0;
    end
    else if ( core_wen & ((or_11_cse & main_stage_v_1) | main_stage_v_2_mx0c1) )
        begin
      main_stage_v_2 <= ~ main_stage_v_2_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_addend_larger_qr_1_lpi_1_dfm_4 <= 49'b0;
      FpAdd_8U_23U_addend_smaller_qr_1_lpi_1_dfm_4 <= 49'b0;
    end
    else if ( FpAdd_8U_23U_addend_larger_and_cse ) begin
      FpAdd_8U_23U_addend_larger_qr_1_lpi_1_dfm_4 <= MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_1_sva,
          FpAdd_8U_23U_addend_larger_asn_19_mx0w1, and_dcpl_390);
      FpAdd_8U_23U_addend_smaller_qr_1_lpi_1_dfm_4 <= MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_19_mx0w1,
          FpAdd_8U_23U_a_int_mant_p1_1_sva, and_dcpl_390);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_4 <=
          1'b0;
      inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_11 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_is_addition_and_cse ) begin
      inp_lookup_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_4 <=
          inp_lookup_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3;
      inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_11 <= IsZero_6U_10U_7_IsZero_6U_10U_7_and_itm_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFractionToFloat_35U_6U_10U_if_else_mux_2_itm_2 <= 10'b0;
    end
    else if ( core_wen & ((or_11_cse & inp_lookup_1_FpMantRNE_36U_11U_else_and_tmp)
        | and_861_rgt) & (mux_111_nl) ) begin
      FpFractionToFloat_35U_6U_10U_if_else_mux_2_itm_2 <= MUX_v_10_2_2((FpMantRNE_36U_11U_else_ac_int_cctor_2_sva[10:1]),
          (FpFractionToFloat_35U_6U_10U_if_else_else_FpFractionToFloat_35U_6U_10U_if_else_else_and_nl),
          and_861_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFractionToFloat_35U_6U_10U_is_zero_1_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & FpFractionToFloat_35U_6U_10U_is_zero_FpFractionToFloat_35U_6U_10U_is_zero_or_3_cse
        & (mux_114_nl) ) begin
      FpFractionToFloat_35U_6U_10U_is_zero_1_lpi_1_dfm_5 <= MUX_s_1_2_2(FpFractionToFloat_35U_6U_10U_is_zero_1_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_2_land_1_lpi_1_dfm_st_6, and_dcpl_394);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_7_1_1 <= 1'b0;
      FpMul_6U_10U_2_lor_6_lpi_1_dfm_st_3 <= 1'b0;
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_4 <= 1'b0;
      chn_inp_in_crt_sva_2_347_1 <= 1'b0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_14 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_7_1_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_6_1_1,
          inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_mx0w1,
          and_dcpl_394);
      FpMul_6U_10U_2_lor_6_lpi_1_dfm_st_3 <= MUX_s_1_2_2(or_5873_cse, IsNaN_8U_23U_land_1_lpi_1_dfm_st_3,
          and_dcpl_394);
      IsNaN_8U_23U_land_1_lpi_1_dfm_st_4 <= MUX_s_1_2_2(IsNaN_8U_23U_land_1_lpi_1_dfm_st_3,
          IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_13, and_dcpl_393);
      chn_inp_in_crt_sva_2_347_1 <= MUX_s_1_2_2(FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_5,
          (chn_inp_in_crt_sva_1_739_395_1[16]), and_dcpl_394);
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_14 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_13,
          (IsNaN_6U_10U_6_IsNaN_6U_10U_6_nor_nl), and_dcpl_393);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_9 <= 4'b0;
      inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_5_1 <= 1'b0;
      inp_lookup_1_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_4 <= 35'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_17_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_9 <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_8;
      inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_5_1 <= (IntLeadZero_35U_leading_sign_35_0_rtn_1_sva_2[5])
          & (~(inp_lookup_1_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_itm_5_1
          & (~ inp_lookup_1_FpMantRNE_36U_11U_else_and_tmp))) & (~ FpFractionToFloat_35U_6U_10U_is_zero_1_lpi_1_dfm_mx0w0);
      inp_lookup_1_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_4 <= inp_lookup_1_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFractionToFloat_35U_6U_10U_1_o_mant_1_lpi_1_dfm_8 <= 10'b0;
      FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_6_5_1 <= 1'b0;
      FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_6_4_0_1 <= 5'b0;
    end
    else if ( FpFractionToFloat_35U_6U_10U_1_o_mant_and_12_cse ) begin
      FpFractionToFloat_35U_6U_10U_1_o_mant_1_lpi_1_dfm_8 <= FpFractionToFloat_35U_6U_10U_1_o_mant_1_lpi_1_dfm_3_mx0w0;
      FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_6_5_1 <= FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_3_5_mx0w0;
      FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_6_4_0_1 <= FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_3_4_0_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_7_itm <= 2'b0;
    end
    else if ( (~ (mux_2045_nl)) & core_wen & (cfg_precision_1_sva_st_90==2'b10) &
        main_stage_v_1 & (~(nor_1896_cse | (chn_inp_in_crt_sva_1_739_395_1[341])))
        ) begin
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_7_itm <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_mux1h_1_itm[9:8];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_7_1_itm <= 8'b0;
    end
    else if ( ((~ (mux_2047_nl)) | (chn_inp_in_crt_sva_1_739_395_1[341])) & core_wen
        & (cfg_precision_1_sva_st_90==2'b10) & or_11_cse & main_stage_v_1 ) begin
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_7_1_itm <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_mux1h_1_itm[7:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_4_0_1 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_127_nl)) ) begin
      inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_4_0_1 <= ~(MUX_v_5_2_2((FpFractionToFloat_35U_6U_10U_nor_nl),
          5'b11111, FpFractionToFloat_35U_6U_10U_is_zero_1_lpi_1_dfm_mx0w0));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_st_91 <= 2'b0;
      chn_inp_in_crt_sva_2_127_0_1 <= 128'b0;
      chn_inp_in_crt_sva_2_331_268_1 <= 64'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_7_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_7_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_16 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_7_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_7_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_16 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_7_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_7_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_16 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_7_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_7_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_16 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_16 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_16 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_16 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_16 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_7_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_7_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_19 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_7_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_7_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_19 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_19 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_7_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_7_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_19 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_7_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_7_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_19 <= 4'b0;
      IsNaN_6U_10U_2_land_lpi_1_dfm_16 <= 1'b0;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_16 <= 1'b0;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_16 <= 1'b0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_16 <= 1'b0;
      chn_inp_in_crt_sva_2_739_736_1 <= 4'b0;
    end
    else if ( cfg_precision_and_4_cse ) begin
      cfg_precision_1_sva_st_91 <= cfg_precision_1_sva_st_90;
      chn_inp_in_crt_sva_2_127_0_1 <= chn_inp_in_crt_sva_1_127_0_1;
      chn_inp_in_crt_sva_2_331_268_1 <= chn_inp_in_crt_sva_1_331_268_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_7_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_6_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_7_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_6_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_16 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_15;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_7_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_6_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_7_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_6_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_16 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_15;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_7_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_6_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_7_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_6_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_16 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_15;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_7_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_6_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_7_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_6_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_16 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_15;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_16 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_15;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_16 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_15;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_16 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_15;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_16 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_15;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_7_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_6_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_7_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_6_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_19 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_18;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_7_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_6_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_7_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_6_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_19 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_18;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_19 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_18;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_7_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_6_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_7_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_6_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_19 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_18;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_7_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_6_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_7_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_6_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_19 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_18;
      IsNaN_6U_10U_2_land_lpi_1_dfm_16 <= IsNaN_6U_10U_2_land_lpi_1_dfm_15;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_16 <= IsNaN_6U_10U_2_land_3_lpi_1_dfm_15;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_16 <= IsNaN_6U_10U_2_land_2_lpi_1_dfm_15;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_16 <= IsNaN_6U_10U_2_land_1_lpi_1_dfm_15;
      chn_inp_in_crt_sva_2_739_736_1 <= chn_inp_in_crt_sva_1_739_395_1[344:341];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_addend_larger_qr_2_lpi_1_dfm_4 <= 49'b0;
      FpAdd_8U_23U_addend_smaller_qr_2_lpi_1_dfm_4 <= 49'b0;
    end
    else if ( FpAdd_8U_23U_addend_larger_and_1_cse ) begin
      FpAdd_8U_23U_addend_larger_qr_2_lpi_1_dfm_4 <= MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_2_sva,
          FpAdd_8U_23U_addend_larger_asn_13_mx0w1, and_dcpl_398);
      FpAdd_8U_23U_addend_smaller_qr_2_lpi_1_dfm_4 <= MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_13_mx0w1,
          FpAdd_8U_23U_a_int_mant_p1_2_sva, and_dcpl_398);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_4 <=
          1'b0;
      inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_10 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_is_addition_and_2_cse ) begin
      inp_lookup_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_4 <=
          inp_lookup_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3;
      inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_10 <= ~(inp_lookup_2_IsZero_6U_10U_2_aif_IsZero_6U_10U_2_aelse_nor_itm_2
          & FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_6_1_1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFractionToFloat_35U_6U_10U_if_else_mux_6_itm_2 <= 10'b0;
    end
    else if ( core_wen & ((or_11_cse & inp_lookup_2_FpMantRNE_36U_11U_else_and_tmp)
        | and_869_rgt) & (mux_134_nl) ) begin
      FpFractionToFloat_35U_6U_10U_if_else_mux_6_itm_2 <= MUX_v_10_2_2((FpMantRNE_36U_11U_else_ac_int_cctor_3_sva[10:1]),
          (FpFractionToFloat_35U_6U_10U_if_else_else_FpFractionToFloat_35U_6U_10U_if_else_else_and_1_nl),
          and_869_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFractionToFloat_35U_6U_10U_is_zero_2_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & FpFractionToFloat_35U_6U_10U_is_zero_FpFractionToFloat_35U_6U_10U_is_zero_or_2_cse
        & (mux_137_nl) ) begin
      FpFractionToFloat_35U_6U_10U_is_zero_2_lpi_1_dfm_5 <= MUX_s_1_2_2(FpFractionToFloat_35U_6U_10U_is_zero_2_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_2_land_2_lpi_1_dfm_st_6, and_dcpl_402);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_7_1_1 <= 1'b0;
      FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_3 <= 1'b0;
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_4 <= 1'b0;
      chn_inp_in_crt_sva_2_363_1 <= 1'b0;
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_1_itm_6 <= 1'b0;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_14 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_18_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_7_1_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_6_1_1,
          inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_mx0w1,
          and_dcpl_402);
      FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_3 <= MUX_s_1_2_2(or_5890_cse, IsNaN_8U_23U_land_2_lpi_1_dfm_4,
          and_dcpl_402);
      IsNaN_8U_23U_land_2_lpi_1_dfm_st_4 <= MUX_s_1_2_2(IsNaN_8U_23U_land_2_lpi_1_dfm_4,
          IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_13, and_dcpl_401);
      chn_inp_in_crt_sva_2_363_1 <= MUX_s_1_2_2(FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_5,
          (chn_inp_in_crt_sva_1_739_395_1[32]), and_dcpl_402);
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_1_itm_6 <= MUX_s_1_2_2((IsZero_6U_10U_1_IsZero_6U_10U_1_and_1_nl),
          IsZero_6U_10U_5_IsZero_6U_10U_5_and_1_itm_2, and_dcpl_401);
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_14 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_13,
          (IsNaN_6U_10U_6_IsNaN_6U_10U_6_nor_1_nl), and_dcpl_401);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_9 <= 4'b0;
      inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_6_5_1 <= 1'b0;
      inp_lookup_2_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_4 <= 35'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_19_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_9 <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_8;
      inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_6_5_1 <= (IntLeadZero_35U_leading_sign_35_0_rtn_2_sva_2[5])
          & (~(inp_lookup_2_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_itm_5_1
          & (~ inp_lookup_2_FpMantRNE_36U_11U_else_and_tmp))) & (~ FpFractionToFloat_35U_6U_10U_is_zero_2_lpi_1_dfm_mx0w0);
      inp_lookup_2_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_4 <= inp_lookup_2_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFractionToFloat_35U_6U_10U_1_o_mant_2_lpi_1_dfm_8 <= 10'b0;
      FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_6_5_1 <= 1'b0;
      FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_6_4_0_1 <= 5'b0;
    end
    else if ( FpFractionToFloat_35U_6U_10U_1_o_mant_and_13_cse ) begin
      FpFractionToFloat_35U_6U_10U_1_o_mant_2_lpi_1_dfm_8 <= FpFractionToFloat_35U_6U_10U_1_o_mant_2_lpi_1_dfm_3_mx0w0;
      FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_6_5_1 <= FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_3_5_mx0w0;
      FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_6_4_0_1 <= FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_3_4_0_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_7_itm <= 2'b0;
    end
    else if ( (~ (mux_2050_nl)) & core_wen & (cfg_precision_1_sva_st_90==2'b10) &
        main_stage_v_1 & (~(nor_1896_cse | (chn_inp_in_crt_sva_1_739_395_1[342])))
        ) begin
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_7_itm <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_mux1h_3_itm[9:8];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_7_1_itm <= 8'b0;
    end
    else if ( ((~ (mux_2051_nl)) | (chn_inp_in_crt_sva_1_739_395_1[342])) & core_wen
        & (cfg_precision_1_sva_st_90==2'b10) & or_11_cse & main_stage_v_1 ) begin
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_7_1_itm <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_mux1h_3_itm[7:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_6_4_0_1 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_149_nl)) ) begin
      inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_6_4_0_1 <= ~(MUX_v_5_2_2((FpFractionToFloat_35U_6U_10U_nor_1_nl),
          5'b11111, FpFractionToFloat_35U_6U_10U_is_zero_2_lpi_1_dfm_mx0w0));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_addend_larger_qr_3_lpi_1_dfm_4 <= 49'b0;
      FpAdd_8U_23U_addend_smaller_qr_3_lpi_1_dfm_4 <= 49'b0;
    end
    else if ( FpAdd_8U_23U_addend_larger_and_2_cse ) begin
      FpAdd_8U_23U_addend_larger_qr_3_lpi_1_dfm_4 <= MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_3_sva,
          FpAdd_8U_23U_addend_larger_asn_7_mx0w1, and_dcpl_406);
      FpAdd_8U_23U_addend_smaller_qr_3_lpi_1_dfm_4 <= MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_7_mx0w1,
          FpAdd_8U_23U_a_int_mant_p1_3_sva, and_dcpl_406);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_4 <=
          1'b0;
      inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_11 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_is_addition_and_4_cse ) begin
      inp_lookup_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_4 <=
          inp_lookup_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3;
      inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_11 <= IsZero_6U_10U_7_IsZero_6U_10U_7_and_2_itm_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFractionToFloat_35U_6U_10U_if_else_mux_10_itm_2 <= 10'b0;
    end
    else if ( core_wen & ((or_11_cse & inp_lookup_3_FpMantRNE_36U_11U_else_and_tmp)
        | and_877_rgt) & (mux_156_nl) ) begin
      FpFractionToFloat_35U_6U_10U_if_else_mux_10_itm_2 <= MUX_v_10_2_2((FpMantRNE_36U_11U_else_ac_int_cctor_4_sva[10:1]),
          (FpFractionToFloat_35U_6U_10U_if_else_else_FpFractionToFloat_35U_6U_10U_if_else_else_and_2_nl),
          and_877_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFractionToFloat_35U_6U_10U_is_zero_3_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & FpFractionToFloat_35U_6U_10U_is_zero_FpFractionToFloat_35U_6U_10U_is_zero_or_1_cse
        & (mux_159_nl) ) begin
      FpFractionToFloat_35U_6U_10U_is_zero_3_lpi_1_dfm_5 <= MUX_s_1_2_2(FpFractionToFloat_35U_6U_10U_is_zero_3_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_2_land_3_lpi_1_dfm_st_6, and_dcpl_410);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_7_1_1 <= 1'b0;
      FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_3 <= 1'b0;
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_4 <= 1'b0;
      chn_inp_in_crt_sva_2_379_1 <= 1'b0;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_14 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_20_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_7_1_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_6_1_1,
          inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_mx0w1,
          and_dcpl_410);
      FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_3 <= MUX_s_1_2_2(FpMul_6U_10U_2_if_2_FpMul_6U_10U_2_if_2_or_5_tmp,
          IsNaN_8U_23U_land_3_lpi_1_dfm_4, and_dcpl_410);
      IsNaN_8U_23U_land_3_lpi_1_dfm_st_4 <= MUX_s_1_2_2(IsNaN_8U_23U_land_3_lpi_1_dfm_4,
          IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_13, and_dcpl_409);
      chn_inp_in_crt_sva_2_379_1 <= MUX_s_1_2_2(FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_5,
          (chn_inp_in_crt_sva_1_739_395_1[48]), and_dcpl_410);
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_14 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_13,
          (IsNaN_6U_10U_6_IsNaN_6U_10U_6_nor_2_nl), and_dcpl_409);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_9 <= 4'b0;
      inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_6_5_1 <= 1'b0;
      inp_lookup_3_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_4 <= 35'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_21_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_9 <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_8;
      inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_6_5_1 <= (IntLeadZero_35U_leading_sign_35_0_rtn_3_sva_2[5])
          & (~(inp_lookup_3_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_itm_5_1
          & (~ inp_lookup_3_FpMantRNE_36U_11U_else_and_tmp))) & (~ FpFractionToFloat_35U_6U_10U_is_zero_3_lpi_1_dfm_mx0w0);
      inp_lookup_3_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_4 <= inp_lookup_3_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFractionToFloat_35U_6U_10U_1_o_mant_3_lpi_1_dfm_8 <= 10'b0;
      FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_6_5_1 <= 1'b0;
      FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_6_4_0_1 <= 5'b0;
    end
    else if ( FpFractionToFloat_35U_6U_10U_1_o_mant_and_14_cse ) begin
      FpFractionToFloat_35U_6U_10U_1_o_mant_3_lpi_1_dfm_8 <= FpFractionToFloat_35U_6U_10U_1_o_mant_3_lpi_1_dfm_3_mx0w0;
      FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_6_5_1 <= FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_3_5_mx0w0;
      FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_6_4_0_1 <= FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_3_4_0_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_3_lpi_1_dfm_9 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_7_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_3_lpi_1_dfm_10 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_and_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_3_lpi_1_dfm_9 <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_3_lpi_1_dfm_8;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_7_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_6_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_3_lpi_1_dfm_10 <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_3_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_6_4_0_1 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_169_nl)) ) begin
      inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_6_4_0_1 <= ~(MUX_v_5_2_2((FpFractionToFloat_35U_6U_10U_nor_2_nl),
          5'b11111, FpFractionToFloat_35U_6U_10U_is_zero_3_lpi_1_dfm_mx0w0));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_addend_larger_qr_lpi_1_dfm_4 <= 49'b0;
      FpAdd_8U_23U_addend_smaller_qr_lpi_1_dfm_4 <= 49'b0;
    end
    else if ( FpAdd_8U_23U_addend_larger_and_3_cse ) begin
      FpAdd_8U_23U_addend_larger_qr_lpi_1_dfm_4 <= MUX_v_49_2_2(FpAdd_8U_23U_a_int_mant_p1_sva,
          FpAdd_8U_23U_addend_larger_asn_1_mx0w1, and_dcpl_412);
      FpAdd_8U_23U_addend_smaller_qr_lpi_1_dfm_4 <= MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_asn_1_mx0w1,
          FpAdd_8U_23U_a_int_mant_p1_sva, and_dcpl_412);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_4 <=
          1'b0;
      inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_10 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_is_addition_and_6_cse ) begin
      inp_lookup_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_4 <=
          inp_lookup_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3;
      inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_10 <= ~(inp_lookup_4_IsZero_6U_10U_2_aif_IsZero_6U_10U_2_aelse_nor_itm_2
          & FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_6_0_1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFractionToFloat_35U_6U_10U_if_else_mux_14_itm_2 <= 10'b0;
    end
    else if ( core_wen & ((or_11_cse & inp_lookup_4_FpMantRNE_36U_11U_else_and_tmp)
        | and_883_rgt) & (mux_175_nl) ) begin
      FpFractionToFloat_35U_6U_10U_if_else_mux_14_itm_2 <= MUX_v_10_2_2((FpMantRNE_36U_11U_else_ac_int_cctor_sva[10:1]),
          (FpFractionToFloat_35U_6U_10U_if_else_else_FpFractionToFloat_35U_6U_10U_if_else_else_and_3_nl),
          and_883_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFractionToFloat_35U_6U_10U_is_zero_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & FpFractionToFloat_35U_6U_10U_is_zero_FpFractionToFloat_35U_6U_10U_is_zero_or_cse
        & (mux_177_nl) ) begin
      FpFractionToFloat_35U_6U_10U_is_zero_lpi_1_dfm_5 <= MUX_s_1_2_2(FpFractionToFloat_35U_6U_10U_is_zero_lpi_1_dfm_mx0w0,
          IsNaN_8U_23U_2_land_lpi_1_dfm_st_6, and_dcpl_416);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_7_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_7_0_1 <= 1'b0;
      FpMul_6U_10U_2_lor_1_lpi_1_dfm_st_3 <= 1'b0;
      IsNaN_8U_23U_land_lpi_1_dfm_st_4 <= 1'b0;
      chn_inp_in_crt_sva_2_395_1 <= 1'b0;
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_3_itm_6 <= 1'b0;
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_14 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_22_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_7_1_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_6_1_1,
          inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_mx0w1,
          and_dcpl_416);
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_7_0_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_6_0_1,
          inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_mx0w1,
          and_dcpl_416);
      FpMul_6U_10U_2_lor_1_lpi_1_dfm_st_3 <= MUX_s_1_2_2(FpMul_6U_10U_2_if_2_FpMul_6U_10U_2_if_2_or_7_tmp,
          IsNaN_8U_23U_land_lpi_1_dfm_4, and_dcpl_416);
      IsNaN_8U_23U_land_lpi_1_dfm_st_4 <= MUX_s_1_2_2(IsNaN_8U_23U_land_lpi_1_dfm_4,
          FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2, and_dcpl_415);
      chn_inp_in_crt_sva_2_395_1 <= MUX_s_1_2_2((chn_inp_in_crt_sva_1_739_395_1[0]),
          (chn_inp_in_crt_sva_1_739_395_1[64]), and_dcpl_416);
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_3_itm_6 <= MUX_s_1_2_2((IsZero_6U_10U_1_IsZero_6U_10U_1_and_3_nl),
          IsZero_6U_10U_5_IsZero_6U_10U_5_and_3_itm_2, and_dcpl_415);
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_14 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_lpi_1_dfm_st_13,
          (IsNaN_6U_10U_6_IsNaN_6U_10U_6_nor_3_nl), and_dcpl_415);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_9 <= 4'b0;
      inp_lookup_else_if_a0_15_10_lpi_1_dfm_6_5_1 <= 1'b0;
      inp_lookup_4_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_4 <= 35'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_24_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_9 <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_8;
      inp_lookup_else_if_a0_15_10_lpi_1_dfm_6_5_1 <= (IntLeadZero_35U_leading_sign_35_0_rtn_sva_2[5])
          & (~(inp_lookup_4_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_itm_5_1
          & (~ inp_lookup_4_FpMantRNE_36U_11U_else_and_tmp))) & (~ FpFractionToFloat_35U_6U_10U_is_zero_lpi_1_dfm_mx0w0);
      inp_lookup_4_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_4 <= inp_lookup_4_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFractionToFloat_35U_6U_10U_1_o_mant_lpi_1_dfm_8 <= 10'b0;
      FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_6_5_1 <= 1'b0;
      FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_6_4_0_1 <= 5'b0;
    end
    else if ( FpFractionToFloat_35U_6U_10U_1_o_mant_and_15_cse ) begin
      FpFractionToFloat_35U_6U_10U_1_o_mant_lpi_1_dfm_8 <= FpFractionToFloat_35U_6U_10U_1_o_mant_lpi_1_dfm_3_mx0w0;
      FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_6_5_1 <= FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_3_5_mx0w0;
      FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_6_4_0_1 <= FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_3_4_0_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_7_itm <= 2'b0;
    end
    else if ( (~ (mux_2053_nl)) & core_wen & (cfg_precision_1_sva_st_90==2'b10) &
        main_stage_v_1 & (~(nor_1896_cse | (chn_inp_in_crt_sva_1_739_395_1[344])))
        ) begin
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_7_itm <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_mux1h_6_itm[9:8];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_7_1_itm <= 8'b0;
    end
    else if ( ((~ (mux_2054_nl)) | (chn_inp_in_crt_sva_1_739_395_1[344])) & core_wen
        & (cfg_precision_1_sva_st_90==2'b10) & or_11_cse & main_stage_v_1 ) begin
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_7_1_itm <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_mux1h_6_itm[7:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_if_a0_15_10_lpi_1_dfm_6_4_0_1 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_187_nl) ) begin
      inp_lookup_else_if_a0_15_10_lpi_1_dfm_6_4_0_1 <= ~(MUX_v_5_2_2((FpFractionToFloat_35U_6U_10U_nor_3_nl),
          5'b11111, FpFractionToFloat_35U_6U_10U_is_zero_lpi_1_dfm_mx0w0));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_3 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_419 | main_stage_v_3_mx0c1) ) begin
      main_stage_v_3 <= ~ main_stage_v_3_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_int_mant_2_sva_5 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_189_nl) ) begin
      FpAdd_8U_23U_int_mant_2_sva_5 <= inp_lookup_1_FpNormalize_8U_49U_else_lshift_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_3_127_0_1 <= 128'b0;
      cfg_precision_1_sva_st_80 <= 2'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_8_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_8_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_17 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_8_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_8_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_17 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_8_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_8_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_17 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_8_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_8_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_17 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_17 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_17 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_17 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_17 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_8_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_8_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_20 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_8_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_8_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_20 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_20 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_8_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_8_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_20 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_8_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_8_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_20 <= 4'b0;
      FpAdd_8U_23U_o_sign_lpi_1_dfm_8 <= 1'b0;
      FpMul_6U_10U_2_o_sign_lpi_1_dfm_6 <= 1'b0;
      FpMul_6U_10U_2_o_sign_3_lpi_1_dfm_6 <= 1'b0;
      FpMul_6U_10U_2_o_sign_2_lpi_1_dfm_6 <= 1'b0;
      FpMul_6U_10U_2_o_sign_1_lpi_1_dfm_6 <= 1'b0;
      FpMul_6U_10U_1_o_sign_lpi_1_dfm_6 <= 1'b0;
      IsNaN_6U_10U_2_land_lpi_1_dfm_17 <= 1'b0;
      FpMul_6U_10U_1_o_sign_3_lpi_1_dfm_6 <= 1'b0;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_17 <= 1'b0;
      FpMul_6U_10U_1_o_sign_2_lpi_1_dfm_6 <= 1'b0;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_17 <= 1'b0;
      FpMul_6U_10U_1_o_sign_1_lpi_1_dfm_6 <= 1'b0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_17 <= 1'b0;
      chn_inp_in_crt_sva_3_739_736_1 <= 4'b0;
    end
    else if ( and_3624_cse ) begin
      chn_inp_in_crt_sva_3_127_0_1 <= chn_inp_in_crt_sva_2_127_0_1;
      cfg_precision_1_sva_st_80 <= cfg_precision_1_sva_st_91;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_8_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_7_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_8_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_7_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_17 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_16;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_8_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_7_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_8_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_7_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_17 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_16;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_8_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_7_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_8_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_7_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_17 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_16;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_8_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_7_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_8_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_7_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_17 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_16;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_17 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_16;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_17 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_16;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_17 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_16;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_17 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_16;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_8_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_7_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_8_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_7_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_20 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_19;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_8_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_7_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_8_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_7_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_20 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_19;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_20 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_19;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_8_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_7_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_8_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_7_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_20 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_19;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_8_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_7_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_8_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_7_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_20 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_19;
      FpAdd_8U_23U_o_sign_lpi_1_dfm_8 <= FpAdd_8U_23U_o_sign_lpi_1_dfm_7;
      FpMul_6U_10U_2_o_sign_lpi_1_dfm_6 <= FpMul_6U_10U_2_o_sign_lpi_1_dfm_mx0w0;
      FpMul_6U_10U_2_o_sign_3_lpi_1_dfm_6 <= FpMul_6U_10U_2_o_sign_3_lpi_1_dfm_mx0w0;
      FpMul_6U_10U_2_o_sign_2_lpi_1_dfm_6 <= FpMul_6U_10U_2_o_sign_2_lpi_1_dfm_mx0w0;
      FpMul_6U_10U_2_o_sign_1_lpi_1_dfm_6 <= FpMul_6U_10U_2_o_sign_1_lpi_1_dfm_mx0w0;
      FpMul_6U_10U_1_o_sign_lpi_1_dfm_6 <= FpMul_6U_10U_1_o_sign_lpi_1_dfm_mx0w0;
      IsNaN_6U_10U_2_land_lpi_1_dfm_17 <= IsNaN_6U_10U_2_land_lpi_1_dfm_16;
      FpMul_6U_10U_1_o_sign_3_lpi_1_dfm_6 <= FpMul_6U_10U_1_o_sign_3_lpi_1_dfm_mx0w0;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_17 <= IsNaN_6U_10U_2_land_3_lpi_1_dfm_16;
      FpMul_6U_10U_1_o_sign_2_lpi_1_dfm_6 <= FpMul_6U_10U_1_o_sign_2_lpi_1_dfm_mx0w0;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_17 <= IsNaN_6U_10U_2_land_2_lpi_1_dfm_16;
      FpMul_6U_10U_1_o_sign_1_lpi_1_dfm_6 <= FpMul_6U_10U_1_o_sign_1_lpi_1_dfm_mx0w0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_17 <= IsNaN_6U_10U_2_land_1_lpi_1_dfm_16;
      chn_inp_in_crt_sva_3_739_736_1 <= chn_inp_in_crt_sva_2_739_736_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_3_510_480_reg <= 8'b0;
    end
    else if ( and_3463_cse & (~((~ (mux_1870_nl)) & and_dcpl_78)) ) begin
      reg_chn_inp_in_crt_sva_3_510_480_reg <= reg_chn_inp_in_crt_sva_2_510_480_itm[11:4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_3_510_480_1_reg <= 23'b0;
    end
    else if ( (mux_2225_nl) & core_wen ) begin
      reg_chn_inp_in_crt_sva_3_510_480_1_reg <= MUX_v_23_2_2((and_3421_nl), ({(reg_chn_inp_in_crt_sva_2_510_480_itm[3:0])
          , reg_chn_inp_in_crt_sva_2_510_480_1_itm}), and_894_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_3_49_1_1 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_196_nl)) ) begin
      FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_3_49_1_1 <= z_out[49:1];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_2 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_427 | and_899_rgt | and_901_rgt | and_903_rgt)
        & (~ mux_197_itm) ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_1_sva_2 <= MUX1HOT_s_1_4_2(inp_lookup_1_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1,
          inp_lookup_1_FpMantRNE_22U_11U_2_else_and_tmp, FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_7_0_1,
          FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_6_5_1, {and_dcpl_427
          , and_899_rgt , and_901_rgt , and_903_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_o_expo_1_lpi_1_dfm_10 <= 8'b0;
    end
    else if ( FpAdd_8U_23U_o_expo_and_cse & (and_907_rgt | and_912_rgt | and_915_rgt
        | and_918_rgt) & (mux_200_nl) ) begin
      FpAdd_8U_23U_o_expo_1_lpi_1_dfm_10 <= MUX1HOT_v_8_4_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_nl),
          FpAdd_8U_23U_o_expo_1_lpi_1_dfm_7_mx1w1, (inp_lookup_1_FpAdd_8U_23U_if_3_if_acc_nl),
          reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_7_1_itm, {and_907_rgt
          , and_912_rgt , and_915_rgt , and_918_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_3_331_268_1 <= 64'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_201_nl) ) begin
      chn_inp_in_crt_sva_3_331_268_1 <= chn_inp_in_crt_sva_2_331_268_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_itm_2
          <= 1'b0;
      inp_lookup_1_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_itm_2
          <= 30'b0;
    end
    else if ( IntSignedShiftRight_50U_5U_32U_obits_fixed_and_cse ) begin
      inp_lookup_1_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_itm_2
          <= ~((~((IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_1_sva[31])
          | IntSignedShiftRight_50U_5U_32U_obits_fixed_and_unfl_1_sva)) | IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_ovfl_1_sva);
      inp_lookup_1_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_itm_2
          <= ~(MUX_v_30_2_2((inp_lookup_1_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_nl),
          30'b111111111111111111111111111111, IntSignedShiftRight_50U_5U_32U_obits_fixed_and_unfl_1_sva));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_itm_2
          <= 1'b0;
    end
    else if ( core_wen & ((or_tmp_439 & or_11_cse) | and_920_rgt) & (mux_208_nl)
        ) begin
      inp_lookup_1_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_itm_2
          <= MUX_s_1_2_2((inp_lookup_1_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_nl),
          inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_3_5_mx0w1, and_920_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_if_a0_9_0_1_lpi_1_dfm_10 <= 10'b0;
      inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_7_4_0_1 <= 5'b0;
    end
    else if ( inp_lookup_else_if_a0_and_8_cse ) begin
      inp_lookup_else_if_a0_9_0_1_lpi_1_dfm_10 <= inp_lookup_else_if_a0_9_0_1_lpi_1_dfm_3_mx0w0;
      inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_7_4_0_1 <= inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_3_4_0_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_else_2_else_if_if_slc_FpMul_6U_10U_2_else_2_else_if_if_acc_1_5_mdf_1_sva_st_1
          <= 1'b0;
    end
    else if ( FpAdd_8U_23U_o_expo_and_cse & FpMul_6U_10U_2_else_2_else_if_FpMul_6U_10U_2_else_2_else_if_or_3_cse
        & (mux_224_nl) ) begin
      FpMul_6U_10U_2_else_2_else_if_if_slc_FpMul_6U_10U_2_else_2_else_if_if_acc_1_5_mdf_1_sva_st_1
          <= MUX_s_1_2_2(inp_lookup_1_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1,
          FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_3_5_mx1w1, and_dcpl_458);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpMul_6U_10U_2_else_2_else_slc_FpMul_6U_10U_2_p_mant_p1_21_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_226_nl)) ) begin
      inp_lookup_1_FpMul_6U_10U_2_else_2_else_slc_FpMul_6U_10U_2_p_mant_p1_21_itm_2
          <= inp_lookup_1_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_228_nl)) ) begin
      inp_lookup_1_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4
          <= inp_lookup_1_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_lor_6_lpi_1_dfm_st_4 <= 1'b0;
      FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_3 <= 1'b0;
      IsNaN_6U_10U_6_land_1_lpi_1_dfm_5 <= 1'b0;
      inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4
          <= 1'b0;
      inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4
          <= 1'b0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_15 <= 1'b0;
    end
    else if ( FpMul_6U_10U_2_oelse_1_and_4_cse ) begin
      FpMul_6U_10U_2_lor_6_lpi_1_dfm_st_4 <= MUX_s_1_2_2(FpMul_6U_10U_2_lor_6_lpi_1_dfm_st_3,
          inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_11, and_dcpl_427);
      FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_3 <= MUX_s_1_2_2(or_457_cse, FpMul_6U_10U_2_lor_6_lpi_1_dfm_5,
          and_dcpl_427);
      IsNaN_6U_10U_6_land_1_lpi_1_dfm_5 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_14,
          FpMul_6U_10U_2_lor_6_lpi_1_dfm_st_3, and_dcpl_427);
      inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4
          <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_7_1_1,
          inp_lookup_1_FpMantRNE_22U_11U_2_else_and_tmp, and_dcpl_459);
      inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4
          <= MUX_s_1_2_2(inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0,
          (z_out[49]), and_dcpl_427);
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_15 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_14,
          IsNaN_6U_10U_4_land_1_lpi_1_dfm_mx0w1, and_dcpl_459);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_int_mant_3_sva_5 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_230_nl)) ) begin
      FpAdd_8U_23U_int_mant_3_sva_5 <= inp_lookup_2_FpNormalize_8U_49U_else_lshift_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_3_542_512_reg <= 8'b0;
    end
    else if ( and_3463_cse & (~((~ (mux_1874_nl)) & and_dcpl_78)) ) begin
      reg_chn_inp_in_crt_sva_3_542_512_reg <= reg_chn_inp_in_crt_sva_2_542_512_itm[11:4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_3_542_512_1_reg <= 23'b0;
    end
    else if ( (mux_2241_nl) & core_wen ) begin
      reg_chn_inp_in_crt_sva_3_542_512_1_reg <= MUX_v_23_2_2((and_3422_nl), ({(reg_chn_inp_in_crt_sva_2_542_512_itm[3:0])
          , reg_chn_inp_in_crt_sva_2_542_512_1_itm}), and_931_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_3_49_1_1 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_236_nl)) ) begin
      FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_3_49_1_1 <= z_out_1[49:1];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_2 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_464 | and_936_rgt | and_939_rgt | and_941_rgt)
        & (~ mux_197_itm) ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_2_sva_2 <= MUX1HOT_s_1_4_2(inp_lookup_2_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1,
          inp_lookup_2_FpMantRNE_22U_11U_2_else_and_tmp, FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_7_0_1,
          FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_6_5_1, {and_dcpl_464
          , and_936_rgt , and_939_rgt , and_941_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_o_expo_2_lpi_1_dfm_10 <= 8'b0;
    end
    else if ( FpAdd_8U_23U_o_expo_and_cse & (and_945_rgt | and_950_rgt | and_953_rgt
        | and_956_rgt) & (mux_238_nl) ) begin
      FpAdd_8U_23U_o_expo_2_lpi_1_dfm_10 <= MUX1HOT_v_8_4_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_2_nl),
          FpAdd_8U_23U_o_expo_2_lpi_1_dfm_7_mx1w1, (inp_lookup_2_FpAdd_8U_23U_if_3_if_acc_nl),
          reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_7_1_itm, {and_945_rgt
          , and_950_rgt , and_953_rgt , and_956_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_itm_2
          <= 1'b0;
      inp_lookup_2_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_itm_2
          <= 30'b0;
    end
    else if ( IntSignedShiftRight_50U_5U_32U_obits_fixed_and_3_cse ) begin
      inp_lookup_2_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_itm_2
          <= ~((~((IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_2_sva[31])
          | IntSignedShiftRight_50U_5U_32U_obits_fixed_and_unfl_2_sva)) | IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_ovfl_2_sva);
      inp_lookup_2_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_itm_2
          <= ~(MUX_v_30_2_2((inp_lookup_2_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_nl),
          30'b111111111111111111111111111111, IntSignedShiftRight_50U_5U_32U_obits_fixed_and_unfl_2_sva));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_itm_2
          <= 1'b0;
    end
    else if ( core_wen & IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_2_cse
        & (mux_246_nl) ) begin
      inp_lookup_2_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_itm_2
          <= MUX_s_1_2_2((inp_lookup_2_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_nl),
          inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_3_5_mx0w1, and_dcpl_488);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_if_a0_9_0_2_lpi_1_dfm_10 <= 10'b0;
      inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_7_4_0_1 <= 5'b0;
    end
    else if ( inp_lookup_else_if_a0_and_9_cse ) begin
      inp_lookup_else_if_a0_9_0_2_lpi_1_dfm_10 <= inp_lookup_else_if_a0_9_0_2_lpi_1_dfm_3_mx0w0;
      inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_7_4_0_1 <= inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_3_4_0_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_else_2_else_if_if_slc_FpMul_6U_10U_2_else_2_else_if_if_acc_1_5_mdf_2_sva_st_1
          <= 1'b0;
    end
    else if ( FpAdd_8U_23U_o_expo_and_cse & FpMul_6U_10U_2_else_2_else_if_FpMul_6U_10U_2_else_2_else_if_or_2_cse
        & (mux_263_nl) ) begin
      FpMul_6U_10U_2_else_2_else_if_if_slc_FpMul_6U_10U_2_else_2_else_if_if_acc_1_5_mdf_2_sva_st_1
          <= MUX_s_1_2_2(inp_lookup_2_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1,
          FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_3_5_mx1w1, and_dcpl_495);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpMul_6U_10U_2_else_2_else_slc_FpMul_6U_10U_2_p_mant_p1_21_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_264_nl)) ) begin
      inp_lookup_2_FpMul_6U_10U_2_else_2_else_slc_FpMul_6U_10U_2_p_mant_p1_21_itm_2
          <= inp_lookup_2_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_265_nl) ) begin
      inp_lookup_2_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4
          <= inp_lookup_2_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_4 <= 1'b0;
      FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_3 <= 1'b0;
      IsNaN_6U_10U_6_land_2_lpi_1_dfm_5 <= 1'b0;
      inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4
          <= 1'b0;
      inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4
          <= 1'b0;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_15 <= 1'b0;
    end
    else if ( FpMul_6U_10U_2_oelse_1_and_5_cse ) begin
      FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_4 <= MUX_s_1_2_2(FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_3,
          inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_10, and_dcpl_464);
      FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_3 <= MUX_s_1_2_2(or_519_cse, FpMul_6U_10U_2_lor_7_lpi_1_dfm_5,
          and_dcpl_464);
      IsNaN_6U_10U_6_land_2_lpi_1_dfm_5 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_14,
          FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_3, and_dcpl_464);
      inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4
          <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_7_1_1,
          inp_lookup_2_FpMantRNE_22U_11U_2_else_and_tmp, and_dcpl_488);
      inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4
          <= MUX_s_1_2_2(inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0,
          (z_out_1[49]), and_dcpl_464);
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_15 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_14,
          IsNaN_6U_10U_4_land_2_lpi_1_dfm_mx0w1, and_dcpl_488);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_int_mant_4_sva_5 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_267_nl)) ) begin
      FpAdd_8U_23U_int_mant_4_sva_5 <= inp_lookup_3_FpNormalize_8U_49U_else_lshift_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_3_574_544_reg <= 8'b0;
    end
    else if ( and_3463_cse & (~((~ (mux_1880_nl)) & and_dcpl_78)) ) begin
      reg_chn_inp_in_crt_sva_3_574_544_reg <= reg_chn_inp_in_crt_sva_2_574_544_itm[11:4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_3_574_544_1_reg <= 23'b0;
    end
    else if ( (mux_2258_nl) & core_wen ) begin
      reg_chn_inp_in_crt_sva_3_574_544_1_reg <= MUX_v_23_2_2((and_3423_nl), ({(reg_chn_inp_in_crt_sva_2_574_544_itm[3:0])
          , reg_chn_inp_in_crt_sva_2_574_544_1_itm}), and_969_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_3_49_1_1 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_273_nl)) ) begin
      FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_3_49_1_1 <= z_out_2[49:1];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_2 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_496 | and_973_rgt | and_976_rgt | and_978_rgt)
        & (~ mux_197_itm) ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_3_sva_2 <= MUX1HOT_s_1_4_2(inp_lookup_3_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1,
          inp_lookup_3_FpMantRNE_22U_11U_2_else_and_tmp, FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_7_0_1,
          FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_6_5_1, {and_dcpl_496
          , and_973_rgt , and_976_rgt , and_978_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_o_expo_3_lpi_1_dfm_10 <= 8'b0;
    end
    else if ( FpAdd_8U_23U_o_expo_and_cse & (and_982_rgt | and_987_rgt | and_990_rgt
        | and_993_rgt) & (mux_276_nl) ) begin
      FpAdd_8U_23U_o_expo_3_lpi_1_dfm_10 <= MUX1HOT_v_8_4_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_4_nl),
          FpAdd_8U_23U_o_expo_3_lpi_1_dfm_7_mx1w1, (inp_lookup_3_FpAdd_8U_23U_if_3_if_acc_nl),
          reg_FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_7_1_itm, {and_982_rgt
          , and_987_rgt , and_990_rgt , and_993_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_itm_2
          <= 1'b0;
      inp_lookup_3_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_itm_2
          <= 30'b0;
    end
    else if ( IntSignedShiftRight_50U_5U_32U_obits_fixed_and_6_cse ) begin
      inp_lookup_3_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_itm_2
          <= ~((~((IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_3_sva[31])
          | IntSignedShiftRight_50U_5U_32U_obits_fixed_and_unfl_3_sva)) | IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_ovfl_3_sva);
      inp_lookup_3_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_itm_2
          <= ~(MUX_v_30_2_2((inp_lookup_3_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_nl),
          30'b111111111111111111111111111111, IntSignedShiftRight_50U_5U_32U_obits_fixed_and_unfl_3_sva));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_itm_2
          <= 1'b0;
    end
    else if ( core_wen & IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_1_cse
        & (mux_284_nl) ) begin
      inp_lookup_3_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_itm_2
          <= MUX_s_1_2_2((inp_lookup_3_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_nl),
          inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_3_5_mx0w1, and_dcpl_524);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_if_a0_9_0_3_lpi_1_dfm_10 <= 10'b0;
      inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_7_4_0_1 <= 5'b0;
    end
    else if ( inp_lookup_else_if_a0_and_10_cse ) begin
      inp_lookup_else_if_a0_9_0_3_lpi_1_dfm_10 <= inp_lookup_else_if_a0_9_0_3_lpi_1_dfm_3_mx0w0;
      inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_7_4_0_1 <= inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_3_4_0_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_10 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_8_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_10 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_and_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_10 <= MUX_v_10_2_2(({reg_FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_7_itm
          , reg_FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_7_1_itm}), FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_3_mx1w1,
          and_dcpl_530);
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_8_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_7_1_1,
          FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_3_4_mx0w0, and_dcpl_530);
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_10 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_9,
          FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_3_3_0_mx0w0, and_dcpl_530);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_else_2_else_if_if_slc_FpMul_6U_10U_2_else_2_else_if_if_acc_1_5_mdf_3_sva_st_1
          <= 1'b0;
    end
    else if ( FpAdd_8U_23U_o_expo_and_cse & FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_or_cse
        & (mux_308_nl) ) begin
      FpMul_6U_10U_2_else_2_else_if_if_slc_FpMul_6U_10U_2_else_2_else_if_if_acc_1_5_mdf_3_sva_st_1
          <= MUX_s_1_2_2(inp_lookup_3_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1,
          FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_3_5_mx1w1, and_dcpl_530);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpMul_6U_10U_2_else_2_else_slc_FpMul_6U_10U_2_p_mant_p1_21_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_310_nl)) ) begin
      inp_lookup_3_FpMul_6U_10U_2_else_2_else_slc_FpMul_6U_10U_2_p_mant_p1_21_itm_2
          <= inp_lookup_3_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_312_nl)) ) begin
      inp_lookup_3_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4
          <= inp_lookup_3_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_4 <= 1'b0;
      FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_3 <= 1'b0;
      IsNaN_6U_10U_6_land_3_lpi_1_dfm_5 <= 1'b0;
      inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4
          <= 1'b0;
      inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4
          <= 1'b0;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_15 <= 1'b0;
    end
    else if ( FpMul_6U_10U_2_oelse_1_and_6_cse ) begin
      FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_4 <= MUX_s_1_2_2(FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_3,
          inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_11, and_dcpl_496);
      FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_3 <= MUX_s_1_2_2(or_593_cse, FpMul_6U_10U_2_lor_8_lpi_1_dfm_5,
          and_dcpl_496);
      IsNaN_6U_10U_6_land_3_lpi_1_dfm_5 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_14,
          FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_3, and_dcpl_496);
      inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4
          <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_7_1_1,
          inp_lookup_3_FpMantRNE_22U_11U_2_else_and_tmp, and_dcpl_524);
      inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4
          <= MUX_s_1_2_2(inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0,
          (z_out_2[49]), and_dcpl_496);
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_15 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_14,
          IsNaN_6U_10U_4_land_3_lpi_1_dfm_mx0w1, and_dcpl_524);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_int_mant_1_sva_5 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_313_nl) ) begin
      FpAdd_8U_23U_int_mant_1_sva_5 <= inp_lookup_4_FpNormalize_8U_49U_else_lshift_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_3_606_576_reg <= 8'b0;
    end
    else if ( (cfg_precision_1_sva_st_91==2'b10) & or_11_cse & (chn_inp_in_crt_sva_2_739_736_1[3])
        & main_stage_v_2 & core_wen ) begin
      reg_chn_inp_in_crt_sva_3_606_576_reg <= mux_1993_rgt[30:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_3_606_576_1_reg <= 23'b0;
    end
    else if ( (((~(((~ main_stage_v_3) | (~ (chn_inp_in_crt_sva_3_739_736_1[3]))
        | (cfg_precision_1_sva_st_80!=2'b10) | IsNaN_6U_10U_6_land_lpi_1_dfm_5) &
        nand_701_cse)) & or_11_cse) | (fsm_output[0])) & core_wen ) begin
      reg_chn_inp_in_crt_sva_3_606_576_1_reg <= mux_1993_rgt[22:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_3_49_1_1 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_314_nl)) ) begin
      FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_3_49_1_1 <= z_out_3[49:1];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_sva_2 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_535 | nor_1743_rgt | and_1012_rgt | and_1014_rgt)
        & (~ mux_197_itm) ) begin
      FpAdd_8U_23U_if_3_if_slc_FpAdd_8U_23U_if_3_if_acc_1_7_mdf_sva_2 <= MUX1HOT_s_1_4_2(inp_lookup_4_FpAdd_8U_23U_if_3_if_acc_1_itm_7_1,
          inp_lookup_4_FpMantRNE_22U_11U_2_else_and_tmp, FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_7_0_1,
          FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_6_5_1, {and_dcpl_535 ,
          nor_1743_rgt , and_1012_rgt , and_1014_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_o_expo_lpi_1_dfm_10 <= 8'b0;
    end
    else if ( FpAdd_8U_23U_o_expo_and_cse & (and_1018_rgt | and_1023_rgt | and_1026_rgt
        | and_1029_rgt) & (mux_319_nl) ) begin
      FpAdd_8U_23U_o_expo_lpi_1_dfm_10 <= MUX1HOT_v_8_4_2((FpNormalize_8U_49U_FpNormalize_8U_49U_and_6_nl),
          FpAdd_8U_23U_o_expo_lpi_1_dfm_7_mx1w1, (inp_lookup_4_FpAdd_8U_23U_if_3_if_acc_nl),
          reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_7_1_itm, {and_1018_rgt
          , and_1023_rgt , and_1026_rgt , and_1029_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_itm_2
          <= 1'b0;
      inp_lookup_4_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_itm_2
          <= 30'b0;
    end
    else if ( IntSignedShiftRight_50U_5U_32U_obits_fixed_and_9_cse ) begin
      inp_lookup_4_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_itm_2
          <= ~((~((IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_sva[31]) |
          IntSignedShiftRight_50U_5U_32U_obits_fixed_and_unfl_sva)) | IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_ovfl_sva);
      inp_lookup_4_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_itm_2
          <= ~(MUX_v_30_2_2((inp_lookup_4_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_nl),
          30'b111111111111111111111111111111, IntSignedShiftRight_50U_5U_32U_obits_fixed_and_unfl_sva));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_itm_2
          <= 1'b0;
    end
    else if ( core_wen & IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_cse
        & (mux_335_nl) ) begin
      inp_lookup_4_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_itm_2
          <= MUX_s_1_2_2((inp_lookup_4_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_nl),
          inp_lookup_else_if_a0_15_10_lpi_1_dfm_3_5_mx0w1, and_dcpl_559);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_if_a0_9_0_lpi_1_dfm_10 <= 10'b0;
      inp_lookup_else_if_a0_15_10_lpi_1_dfm_7_4_0_1 <= 5'b0;
    end
    else if ( inp_lookup_else_if_a0_and_11_cse ) begin
      inp_lookup_else_if_a0_9_0_lpi_1_dfm_10 <= inp_lookup_else_if_a0_9_0_lpi_1_dfm_3_mx0w0;
      inp_lookup_else_if_a0_15_10_lpi_1_dfm_7_4_0_1 <= inp_lookup_else_if_a0_15_10_lpi_1_dfm_3_4_0_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_else_2_else_if_if_slc_FpMul_6U_10U_2_else_2_else_if_if_acc_1_5_mdf_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_cse
        & (mux_347_nl) ) begin
      FpMul_6U_10U_2_else_2_else_if_if_slc_FpMul_6U_10U_2_else_2_else_if_if_acc_1_5_mdf_sva_st_2
          <= MUX_s_1_2_2(inp_lookup_4_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_7_0_1, and_dcpl_535);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpMul_6U_10U_2_else_2_else_slc_FpMul_6U_10U_2_p_mant_p1_21_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_348_nl)) ) begin
      inp_lookup_4_FpMul_6U_10U_2_else_2_else_slc_FpMul_6U_10U_2_p_mant_p1_21_itm_2
          <= inp_lookup_4_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_349_nl) ) begin
      inp_lookup_4_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4
          <= inp_lookup_4_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_lor_1_lpi_1_dfm_st_4 <= 1'b0;
      FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_3 <= 1'b0;
      inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4
          <= 1'b0;
      IsNaN_6U_10U_6_land_lpi_1_dfm_5 <= 1'b0;
      inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4
          <= 1'b0;
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_15 <= 1'b0;
    end
    else if ( FpMul_6U_10U_2_oelse_1_and_7_cse ) begin
      FpMul_6U_10U_2_lor_1_lpi_1_dfm_st_4 <= MUX_s_1_2_2(FpMul_6U_10U_2_lor_1_lpi_1_dfm_st_3,
          inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_10, and_dcpl_535);
      FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_3 <= MUX_s_1_2_2(or_648_cse, FpMul_6U_10U_2_lor_1_lpi_1_dfm_5,
          and_dcpl_535);
      inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4
          <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_7_1_1,
          inp_lookup_4_FpMantRNE_22U_11U_2_else_and_tmp, and_dcpl_559);
      IsNaN_6U_10U_6_land_lpi_1_dfm_5 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_lpi_1_dfm_st_14,
          FpMul_6U_10U_2_lor_1_lpi_1_dfm_st_3, and_dcpl_535);
      inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4
          <= MUX_s_1_2_2(inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0,
          (z_out_3[49]), and_dcpl_535);
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_15 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_lpi_1_dfm_st_14,
          IsNaN_6U_10U_4_land_lpi_1_dfm_mx0w1, and_dcpl_559);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_4 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_560 | main_stage_v_4_mx0c1) ) begin
      main_stage_v_4 <= ~ main_stage_v_4_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5
          <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_or_6_cse
        & (mux_351_nl) ) begin
      inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5
          <= MUX_s_1_2_2(inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4,
          inp_lookup_1_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs,
          and_dcpl_565);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_1_st_2 <= 1'b0;
      FpMul_6U_10U_1_lor_6_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_1_is_a_greater_oelse_and_cse ) begin
      FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_1_st_2 <= MUX_s_1_2_2(FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0,
          (FpMul_6U_10U_1_FpMul_6U_10U_1_and_nl), and_dcpl_565);
      FpMul_6U_10U_1_lor_6_lpi_1_dfm_6 <= MUX_s_1_2_2(FpMul_6U_10U_1_lor_6_lpi_1_dfm_5,
          FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_3, and_dcpl_564);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_st_81 <= 2'b0;
      chn_inp_in_crt_sva_4_127_0_1 <= 128'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_9_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_9_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_18 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_9_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_9_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_18 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_9_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_9_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_18 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_9_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_9_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_18 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_18 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_18 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_18 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_18 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_9_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_9_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_21 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_9_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_9_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_21 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_21 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_9_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_9_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_21 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_9_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_9_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_21 <= 4'b0;
      FpMul_6U_10U_2_o_sign_lpi_1_dfm_7 <= 1'b0;
      FpMul_6U_10U_2_o_sign_3_lpi_1_dfm_7 <= 1'b0;
      FpMul_6U_10U_2_o_sign_2_lpi_1_dfm_7 <= 1'b0;
      FpMul_6U_10U_2_o_sign_1_lpi_1_dfm_7 <= 1'b0;
      FpMul_6U_10U_1_o_sign_lpi_1_dfm_7 <= 1'b0;
      IsNaN_6U_10U_2_land_lpi_1_dfm_18 <= 1'b0;
      FpMul_6U_10U_1_o_sign_3_lpi_1_dfm_7 <= 1'b0;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_18 <= 1'b0;
      FpMul_6U_10U_1_o_sign_2_lpi_1_dfm_7 <= 1'b0;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_18 <= 1'b0;
      FpMul_6U_10U_1_o_sign_1_lpi_1_dfm_7 <= 1'b0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_18 <= 1'b0;
      chn_inp_in_crt_sva_4_739_736_1 <= 4'b0;
    end
    else if ( cfg_precision_and_12_cse ) begin
      cfg_precision_1_sva_st_81 <= cfg_precision_1_sva_st_80;
      chn_inp_in_crt_sva_4_127_0_1 <= chn_inp_in_crt_sva_3_127_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_9_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_8_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_9_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_8_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_18 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_17;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_9_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_8_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_9_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_8_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_18 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_17;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_9_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_8_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_9_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_8_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_18 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_17;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_9_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_8_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_9_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_8_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_18 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_17;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_18 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_17;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_18 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_17;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_18 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_17;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_18 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_17;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_9_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_8_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_9_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_8_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_21 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_20;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_9_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_8_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_9_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_8_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_21 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_20;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_21 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_20;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_9_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_8_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_9_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_8_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_21 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_20;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_9_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_8_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_9_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_8_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_21 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_20;
      FpMul_6U_10U_2_o_sign_lpi_1_dfm_7 <= FpMul_6U_10U_2_o_sign_lpi_1_dfm_6;
      FpMul_6U_10U_2_o_sign_3_lpi_1_dfm_7 <= FpMul_6U_10U_2_o_sign_3_lpi_1_dfm_6;
      FpMul_6U_10U_2_o_sign_2_lpi_1_dfm_7 <= FpMul_6U_10U_2_o_sign_2_lpi_1_dfm_6;
      FpMul_6U_10U_2_o_sign_1_lpi_1_dfm_7 <= FpMul_6U_10U_2_o_sign_1_lpi_1_dfm_6;
      FpMul_6U_10U_1_o_sign_lpi_1_dfm_7 <= FpMul_6U_10U_1_o_sign_lpi_1_dfm_6;
      IsNaN_6U_10U_2_land_lpi_1_dfm_18 <= IsNaN_6U_10U_2_land_lpi_1_dfm_17;
      FpMul_6U_10U_1_o_sign_3_lpi_1_dfm_7 <= FpMul_6U_10U_1_o_sign_3_lpi_1_dfm_6;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_18 <= IsNaN_6U_10U_2_land_3_lpi_1_dfm_17;
      FpMul_6U_10U_1_o_sign_2_lpi_1_dfm_7 <= FpMul_6U_10U_1_o_sign_2_lpi_1_dfm_6;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_18 <= IsNaN_6U_10U_2_land_2_lpi_1_dfm_17;
      FpMul_6U_10U_1_o_sign_1_lpi_1_dfm_7 <= FpMul_6U_10U_1_o_sign_1_lpi_1_dfm_6;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_18 <= IsNaN_6U_10U_2_land_1_lpi_1_dfm_17;
      chn_inp_in_crt_sva_4_739_736_1 <= chn_inp_in_crt_sva_3_739_736_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_5_1 <= 1'b0;
      FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_4_1 <= 1'b0;
      FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_3_0_1 <= 4'b0;
      FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_8 <= 10'b0;
    end
    else if ( FpMul_6U_10U_2_o_expo_and_cse ) begin
      FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_5_1 <= MUX_s_1_2_2(FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_3_5_mx1w1,
          FpMul_6U_10U_2_else_2_else_if_if_slc_FpMul_6U_10U_2_else_2_else_if_if_acc_1_5_mdf_1_sva_st_1,
          and_dcpl_575);
      FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_4_1 <= MUX_s_1_2_2(FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_3_4_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_8_1, and_dcpl_575);
      FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_3_0_1 <= MUX_v_4_2_2(FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_3_3_0_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_10, and_dcpl_575);
      FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_8 <= MUX_v_10_2_2(FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_3_mx0w0,
          ({reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_8_reg , reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_8_1_reg}),
          and_dcpl_575);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_8_5_1 <= 1'b0;
      inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_8_4_0_1 <= 5'b0;
    end
    else if ( inp_lookup_else_if_a0_and_12_cse ) begin
      inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_8_5_1 <= inp_lookup_1_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_itm_2;
      inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_8_4_0_1 <= inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_7_4_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_9_1 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_o_expo_and_cse & (and_1049_rgt | and_dcpl_573 | and_1052_rgt)
        & (mux_370_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_9_1 <= MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_8_1,
          FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_3_4_mx1w1, inp_lookup_1_FpMantRNE_22U_11U_1_else_and_tmp,
          {and_1049_rgt , and_dcpl_573 , and_1052_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_o_expo_and_cse & ((and_dcpl_567 & and_dcpl_560) | and_dcpl_573)
        & (mux_380_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_11 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_10,
          FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_3_3_0_mx1w1, and_dcpl_573);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_5_land_1_lpi_1_dfm_6 <= 1'b0;
      IsNaN_6U_10U_5_land_2_lpi_1_dfm_6 <= 1'b0;
      IsNaN_6U_10U_5_land_3_lpi_1_dfm_6 <= 1'b0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_16 <= 1'b0;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_16 <= 1'b0;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_16 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_5_aelse_and_4_cse ) begin
      IsNaN_6U_10U_5_land_1_lpi_1_dfm_6 <= IsNaN_6U_10U_5_land_1_lpi_1_dfm_5;
      IsNaN_6U_10U_5_land_2_lpi_1_dfm_6 <= IsNaN_6U_10U_5_land_2_lpi_1_dfm_5;
      IsNaN_6U_10U_5_land_3_lpi_1_dfm_6 <= IsNaN_6U_10U_5_land_3_lpi_1_dfm_5;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_16 <= IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_15;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_16 <= IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_15;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_16 <= IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_15;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_4 <= 1'b0;
      inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5
          <= 1'b0;
      inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5
          <= 1'b0;
      chn_inp_in_crt_sva_4_411_1 <= 1'b0;
    end
    else if ( FpMul_6U_10U_1_oelse_1_and_5_cse ) begin
      FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_4 <= MUX_s_1_2_2(FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_3,
          IsNaN_8U_23U_3_IsNaN_8U_23U_3_nor_tmp, and_dcpl_564);
      inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5
          <= MUX_s_1_2_2(inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4,
          inp_lookup_1_FpMantRNE_22U_11U_1_else_and_tmp, and_dcpl_565);
      inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5
          <= MUX_s_1_2_2(inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4,
          FpMul_6U_10U_2_lor_6_lpi_1_dfm_st_4, and_dcpl_564);
      chn_inp_in_crt_sva_4_411_1 <= MUX_s_1_2_2(FpMul_6U_10U_2_lor_6_lpi_1_dfm_6,
          inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4,
          and_dcpl_565);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5
          <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_or_5_cse
        & (mux_382_nl) ) begin
      inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5
          <= MUX_s_1_2_2(inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4,
          inp_lookup_2_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs,
          and_dcpl_583);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_1_st_2 <= 1'b0;
      FpMul_6U_10U_1_lor_7_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_1_is_a_greater_oelse_and_1_cse ) begin
      FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_1_st_2 <= MUX_s_1_2_2(FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0,
          (FpMul_6U_10U_1_FpMul_6U_10U_1_and_16_nl), and_dcpl_583);
      FpMul_6U_10U_1_lor_7_lpi_1_dfm_6 <= MUX_s_1_2_2(FpMul_6U_10U_1_lor_7_lpi_1_dfm_5,
          FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_3, and_dcpl_582);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_5_1 <= 1'b0;
      FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_4_1 <= 1'b0;
      FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_3_0_1 <= 4'b0;
      FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_8 <= 10'b0;
    end
    else if ( FpMul_6U_10U_2_o_expo_and_3_cse ) begin
      FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_5_1 <= MUX_s_1_2_2(FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_3_5_mx1w1,
          FpMul_6U_10U_2_else_2_else_if_if_slc_FpMul_6U_10U_2_else_2_else_if_if_acc_1_5_mdf_2_sva_st_1,
          and_dcpl_593);
      FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_4_1 <= MUX_s_1_2_2(FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_3_4_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_8_1, and_dcpl_593);
      FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_3_0_1 <= MUX_v_4_2_2(FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_3_3_0_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_10, and_dcpl_593);
      FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_8 <= MUX_v_10_2_2(FpMul_6U_10U_2_FpMul_6U_10U_2_FpMul_6U_10U_2_nor_5_itm,
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_10, FpMul_6U_10U_2_o_mant_or_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_8_5_1 <= 1'b0;
      inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_8_4_0_1 <= 5'b0;
    end
    else if ( inp_lookup_else_if_a0_and_14_cse ) begin
      inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_8_5_1 <= inp_lookup_2_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_itm_2;
      inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_8_4_0_1 <= inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_7_4_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_9_1 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_o_expo_and_cse & (and_1068_rgt | and_dcpl_591 | and_1071_rgt)
        & (mux_410_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_9_1 <= MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_8_1,
          FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_3_4_mx1w1, inp_lookup_2_FpMantRNE_22U_11U_1_else_and_tmp,
          {and_1068_rgt , and_dcpl_591 , and_1071_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_o_expo_and_cse & ((and_dcpl_585 & and_dcpl_560) | and_dcpl_591)
        & (mux_420_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_11 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_10,
          FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_3_3_0_mx1w1, and_dcpl_591);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_4 <= 1'b0;
      inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5
          <= 1'b0;
      inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5
          <= 1'b0;
      chn_inp_in_crt_sva_4_427_1 <= 1'b0;
    end
    else if ( FpMul_6U_10U_1_oelse_1_and_7_cse ) begin
      FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_4 <= MUX_s_1_2_2(FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_3,
          IsNaN_8U_23U_3_IsNaN_8U_23U_3_nor_1_tmp, and_dcpl_582);
      inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5
          <= MUX_s_1_2_2(inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4,
          inp_lookup_2_FpMantRNE_22U_11U_1_else_and_tmp, and_dcpl_583);
      inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5
          <= MUX_s_1_2_2(inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4,
          FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_4, and_dcpl_582);
      chn_inp_in_crt_sva_4_427_1 <= MUX_s_1_2_2(FpMul_6U_10U_2_lor_7_lpi_1_dfm_6,
          inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4,
          and_dcpl_583);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5
          <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_or_4_cse
        & (mux_422_nl) ) begin
      inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5
          <= MUX_s_1_2_2(inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4,
          inp_lookup_3_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs,
          and_dcpl_601);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_1_st_2 <= 1'b0;
      FpMul_6U_10U_1_lor_8_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_1_is_a_greater_oelse_and_2_cse ) begin
      FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_1_st_2 <= MUX_s_1_2_2(FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0,
          (FpMul_6U_10U_1_FpMul_6U_10U_1_and_17_nl), and_dcpl_601);
      FpMul_6U_10U_1_lor_8_lpi_1_dfm_6 <= MUX_s_1_2_2(FpMul_6U_10U_1_lor_8_lpi_1_dfm_5,
          FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_3, and_dcpl_600);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_5_1 <= 1'b0;
      FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_4_1 <= 1'b0;
      FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_3_0_1 <= 4'b0;
      FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_8 <= 10'b0;
    end
    else if ( FpMul_6U_10U_2_o_expo_and_6_cse ) begin
      FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_5_1 <= MUX_s_1_2_2(FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_3_5_mx1w1,
          FpMul_6U_10U_2_else_2_else_if_if_slc_FpMul_6U_10U_2_else_2_else_if_if_acc_1_5_mdf_3_sva_st_1,
          and_dcpl_611);
      FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_4_1 <= MUX_s_1_2_2(FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_3_4_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_8_1, and_dcpl_611);
      FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_3_0_1 <= MUX_v_4_2_2(FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_3_3_0_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_10, and_dcpl_611);
      FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_8 <= MUX_v_10_2_2(FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_3_mx1w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_10, and_dcpl_611);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_11 <= 10'b0;
    end
    else if ( core_wen & (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_9_mx0c0
        | and_dcpl_609 | FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_9_mx0c2
        | FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_9_mx0c3) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_11 <= MUX1HOT_v_10_4_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_10,
          FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_3_mx0w1, (FpMul_6U_10U_1_p_mant_20_1_3_lpi_1_dfm_3_mx0[19:10]),
          inp_lookup_else_if_a0_9_0_3_lpi_1_dfm_10, {FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_9_mx0c0
          , and_dcpl_609 , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_9_mx0c2
          , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_9_mx0c3});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_8_5_1 <= 1'b0;
      inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_8_4_0_1 <= 5'b0;
    end
    else if ( inp_lookup_else_if_a0_and_16_cse ) begin
      inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_8_5_1 <= inp_lookup_3_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_itm_2;
      inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_8_4_0_1 <= inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_7_4_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_9_1 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_o_expo_and_cse & (and_1099_rgt | and_dcpl_609 | and_1102_rgt)
        & (mux_449_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_9_1 <= MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_8_1,
          FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_4_mx1w1, inp_lookup_3_FpMantRNE_22U_11U_1_else_and_tmp,
          {and_1099_rgt , and_dcpl_609 , and_1102_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( FpAdd_8U_23U_o_expo_and_cse & ((and_dcpl_603 & and_dcpl_560) | and_dcpl_609)
        & (mux_459_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_11 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_10,
          FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_3_0_mx1w1, and_dcpl_609);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_4 <= 1'b0;
      inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5
          <= 1'b0;
      inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5
          <= 1'b0;
      chn_inp_in_crt_sva_4_443_1 <= 1'b0;
    end
    else if ( FpMul_6U_10U_1_oelse_1_and_9_cse ) begin
      FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_4 <= MUX_s_1_2_2(FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_3,
          IsNaN_8U_23U_3_IsNaN_8U_23U_3_nor_2_tmp, and_dcpl_600);
      inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5
          <= MUX_s_1_2_2(inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4,
          inp_lookup_3_FpMantRNE_22U_11U_1_else_and_tmp, and_dcpl_601);
      inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5
          <= MUX_s_1_2_2(inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4,
          FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_4, and_dcpl_600);
      chn_inp_in_crt_sva_4_443_1 <= MUX_s_1_2_2(FpMul_6U_10U_2_lor_8_lpi_1_dfm_6,
          inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4,
          and_dcpl_601);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_2_land_lpi_1_dfm_st_7 <= 1'b0;
      FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_4 <= 1'b0;
      inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4
          <= 1'b0;
      chn_inp_in_crt_sva_4_459_1 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_2_aelse_and_cse ) begin
      IsNaN_8U_23U_2_land_lpi_1_dfm_st_7 <= MUX_s_1_2_2(FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_3,
          inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4,
          and_dcpl_631);
      FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_4 <= MUX_s_1_2_2(FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_3,
          IsNaN_6U_10U_5_land_lpi_1_dfm_5, and_dcpl_630);
      inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4
          <= MUX_s_1_2_2(FpMul_6U_10U_2_else_2_else_if_if_slc_FpMul_6U_10U_2_else_2_else_if_if_acc_1_5_mdf_sva_st_2,
          inp_lookup_4_FpMantRNE_22U_11U_1_else_and_tmp, and_dcpl_631);
      chn_inp_in_crt_sva_4_459_1 <= MUX_s_1_2_2(FpMul_6U_10U_2_lor_1_lpi_1_dfm_6,
          inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4,
          and_dcpl_631);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5
          <= 1'b0;
    end
    else if ( core_wen & FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_4_cse & (~
        (mux_464_nl)) ) begin
      inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5
          <= MUX_s_1_2_2(inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4,
          inp_lookup_4_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs,
          and_dcpl_631);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_1_st_2 <= 1'b0;
      FpMul_6U_10U_1_lor_1_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_1_is_a_greater_oelse_and_3_cse ) begin
      FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_1_st_2 <= MUX_s_1_2_2(FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_1_mx0w0,
          (FpMul_6U_10U_1_FpMul_6U_10U_1_and_18_nl), and_dcpl_631);
      FpMul_6U_10U_1_lor_1_lpi_1_dfm_6 <= MUX_s_1_2_2(FpMul_6U_10U_1_lor_1_lpi_1_dfm_5,
          IsNaN_6U_10U_2_land_lpi_1_dfm_st_15, and_dcpl_630);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_5_1 <= 1'b0;
      FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_4_1 <= 1'b0;
      FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_3_0_1 <= 4'b0;
      FpMul_6U_10U_2_o_mant_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( FpMul_6U_10U_2_o_expo_and_9_cse ) begin
      FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_5_1 <= MUX_s_1_2_2(FpMul_6U_10U_2_o_expo_lpi_1_dfm_3_5_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_8_1, and_dcpl_641);
      FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_4_1 <= MUX_s_1_2_2(FpMul_6U_10U_2_o_expo_lpi_1_dfm_3_4_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_8_0, and_dcpl_641);
      FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_3_0_1 <= MUX_v_4_2_2(FpMul_6U_10U_2_o_expo_lpi_1_dfm_3_3_0_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_10, and_dcpl_641);
      FpMul_6U_10U_2_o_mant_lpi_1_dfm_7 <= MUX_v_10_2_2(FpMul_6U_10U_2_o_mant_lpi_1_dfm_3_mx0w0,
          ({reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_8_reg , reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_8_1_reg}),
          and_dcpl_641);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_4_land_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_5_land_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_4_aelse_and_cse ) begin
      IsNaN_6U_10U_4_land_lpi_1_dfm_5 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_lpi_1_dfm_st_15,
          IsNaN_8U_23U_3_IsNaN_8U_23U_3_nand_3_tmp, and_dcpl_630);
      IsNaN_6U_10U_5_land_lpi_1_dfm_6 <= MUX_s_1_2_2(IsNaN_6U_10U_5_land_lpi_1_dfm_5,
          IsNaN_8U_23U_3_nor_3_tmp, and_dcpl_630);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_if_a0_15_10_lpi_1_dfm_8_5_1 <= 1'b0;
      inp_lookup_else_if_a0_15_10_lpi_1_dfm_8_4_0_1 <= 5'b0;
    end
    else if ( inp_lookup_else_if_a0_and_18_cse ) begin
      inp_lookup_else_if_a0_15_10_lpi_1_dfm_8_5_1 <= inp_lookup_4_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_itm_2;
      inp_lookup_else_if_a0_15_10_lpi_1_dfm_8_4_0_1 <= inp_lookup_else_if_a0_15_10_lpi_1_dfm_7_4_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_9_1 <= 1'b0;
    end
    else if ( core_wen & (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_9_1_mx0c0
        | and_dcpl_639 | FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_9_1_mx0c2)
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_9_1 <= MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_8_1,
          FpMul_6U_10U_1_o_expo_lpi_1_dfm_3_4_mx0w1, inp_lookup_4_FpMantRNE_22U_11U_1_else_and_tmp,
          {FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_9_1_mx0c0 , and_dcpl_639
          , FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_9_1_mx0c2});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & ((and_dcpl_633 & and_dcpl_560) | and_dcpl_639) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_11 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_10,
          FpMul_6U_10U_1_o_expo_lpi_1_dfm_3_3_0_mx0w1, and_dcpl_639);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_5 <= 1'b0;
    end
    else if ( core_wen & ((or_11_cse & main_stage_v_4) | main_stage_v_5_mx0c1) )
        begin
      main_stage_v_5 <= ~ main_stage_v_5_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_2_land_1_lpi_1_dfm_st_7 <= 1'b0;
    end
    else if ( core_wen & FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_3_cse & (mux_471_nl)
        ) begin
      IsNaN_8U_23U_2_land_1_lpi_1_dfm_st_7 <= MUX_s_1_2_2(FpMul_6U_10U_1_lor_6_lpi_1_dfm_6,
          inp_lookup_1_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp, and_dcpl_655);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_int_mant_p1_1_sva_3 <= 50'b0;
    end
    else if ( core_wen & ((or_11_cse & (~ inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5))
        | and_1131_rgt) & (~ (mux_474_nl)) ) begin
      FpAdd_8U_23U_1_int_mant_p1_1_sva_3 <= MUX_v_50_2_2((inp_lookup_1_FpAdd_8U_23U_1_else_2_acc_nl),
          (inp_lookup_1_FpAdd_8U_23U_1_if_2_acc_nl), and_1131_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_st_82 <= 2'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_10_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_10_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_19 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_10_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_10_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_19 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_10_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_10_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_19 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_10_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_10_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_19 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_19 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_19 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_19 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_19 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_10_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_10_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_22 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_10_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_10_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_22 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_22 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_10_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_10_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_22 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_10_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_10_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_22 <= 4'b0;
      IsNaN_6U_10U_2_land_lpi_1_dfm_19 <= 1'b0;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_19 <= 1'b0;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_19 <= 1'b0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_19 <= 1'b0;
      chn_inp_in_crt_sva_5_739_736_1 <= 4'b0;
    end
    else if ( cfg_precision_and_16_cse ) begin
      cfg_precision_1_sva_st_82 <= cfg_precision_1_sva_st_81;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_10_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_9_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_10_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_9_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_19 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_18;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_10_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_9_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_10_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_9_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_19 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_18;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_10_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_9_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_10_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_9_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_19 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_18;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_10_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_9_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_10_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_9_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_19 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_18;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_19 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_18;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_19 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_18;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_19 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_18;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_19 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_18;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_10_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_9_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_10_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_9_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_22 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_21;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_10_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_9_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_10_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_9_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_22 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_21;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_22 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_21;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_10_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_9_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_10_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_9_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_22 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_21;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_10_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_9_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_10_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_9_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_22 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_21;
      IsNaN_6U_10U_2_land_lpi_1_dfm_19 <= IsNaN_6U_10U_2_land_lpi_1_dfm_18;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_19 <= IsNaN_6U_10U_2_land_3_lpi_1_dfm_18;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_19 <= IsNaN_6U_10U_2_land_2_lpi_1_dfm_18;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_19 <= IsNaN_6U_10U_2_land_1_lpi_1_dfm_18;
      chn_inp_in_crt_sva_5_739_736_1 <= chn_inp_in_crt_sva_4_739_736_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_7_itm <= 2'b0;
    end
    else if ( (((mux_2073_nl) & (FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_3_0_1==4'b1111)
        & FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_4_1 & FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_5_1)
        | and_3637_cse | xnor_6_cse) & (cfg_precision_1_sva_st_81==2'b10) & and_dcpl_2185
        & (~(nor_1896_cse | (chn_inp_in_crt_sva_4_739_736_1[0]))) ) begin
      reg_FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_7_itm <= FpMul_6U_10U_2_o_mant_mux1h_1_itm[9:8];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_7_1_itm <= 8'b0;
    end
    else if ( (((mux_2078_nl) & (FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_3_0_1==4'b1111)
        & FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_4_1 & FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_5_1)
        | and_3637_cse | xnor_6_cse | (chn_inp_in_crt_sva_4_739_736_1[0])) & (cfg_precision_1_sva_st_81[1])
        & main_stage_v_4 & core_wen & nor_1883_cse ) begin
      reg_FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_7_1_itm <= FpMul_6U_10U_2_o_mant_mux1h_1_itm[7:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_2_land_2_lpi_1_dfm_st_7 <= 1'b0;
    end
    else if ( core_wen & FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_2_cse & (mux_481_nl)
        ) begin
      IsNaN_8U_23U_2_land_2_lpi_1_dfm_st_7 <= MUX_s_1_2_2(FpMul_6U_10U_1_lor_7_lpi_1_dfm_6,
          inp_lookup_2_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp, and_dcpl_663);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_int_mant_p1_2_sva_3 <= 50'b0;
    end
    else if ( core_wen & ((or_11_cse & (~ inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5))
        | and_1139_rgt) & (~ (mux_484_nl)) ) begin
      FpAdd_8U_23U_1_int_mant_p1_2_sva_3 <= MUX_v_50_2_2((inp_lookup_2_FpAdd_8U_23U_1_else_2_acc_nl),
          (inp_lookup_2_FpAdd_8U_23U_1_if_2_acc_nl), and_1139_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_7_itm <= 2'b0;
    end
    else if ( (((mux_2082_nl) & (FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_3_0_1==4'b1111)
        & FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_4_1 & FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_5_1)
        | and_3663_cse | xnor_4_cse) & (cfg_precision_1_sva_st_81==2'b10) & and_dcpl_2185
        & (~(nor_1896_cse | (chn_inp_in_crt_sva_4_739_736_1[1]))) ) begin
      reg_FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_7_itm <= FpMul_6U_10U_2_o_mant_mux1h_3_itm[9:8];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_7_1_itm <= 8'b0;
    end
    else if ( (((mux_2087_nl) & (FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_3_0_1==4'b1111)
        & FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_4_1 & FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_5_1)
        | and_3663_cse | xnor_4_cse | (chn_inp_in_crt_sva_4_739_736_1[1])) & (cfg_precision_1_sva_st_81[1])
        & main_stage_v_4 & core_wen & nor_1883_cse ) begin
      reg_FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_7_1_itm <= FpMul_6U_10U_2_o_mant_mux1h_3_itm[7:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_2_land_3_lpi_1_dfm_st_7 <= 1'b0;
    end
    else if ( core_wen & FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_1_cse & (~
        (mux_492_nl)) ) begin
      IsNaN_8U_23U_2_land_3_lpi_1_dfm_st_7 <= MUX_s_1_2_2(FpMul_6U_10U_1_lor_8_lpi_1_dfm_6,
          inp_lookup_3_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp, and_dcpl_671);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_int_mant_p1_3_sva_3 <= 50'b0;
    end
    else if ( core_wen & ((or_11_cse & (~ inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5))
        | and_1147_rgt) & (~ (mux_499_nl)) ) begin
      FpAdd_8U_23U_1_int_mant_p1_3_sva_3 <= MUX_v_50_2_2((inp_lookup_3_FpAdd_8U_23U_1_else_2_acc_nl),
          (inp_lookup_3_FpAdd_8U_23U_1_if_2_acc_nl), and_1147_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_6_itm <= 2'b0;
    end
    else if ( ((or_5985_cse & (mux_2089_nl) & (FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_3_0_mx1w1==4'b1111))
        | and_3689_cse | xnor_2_cse) & core_wen & (cfg_precision_1_sva_st_81==2'b10)
        & main_stage_v_4 & nor_1877_cse ) begin
      reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_6_itm <= FpMul_6U_10U_1_o_mant_mux1h_1_itm[9:8];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_6_1_itm <= 8'b0;
    end
    else if ( (mux_2094_nl) & core_wen & (cfg_precision_1_sva_st_81==2'b10) & or_11_cse
        & main_stage_v_4 ) begin
      reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_6_1_itm <= FpMul_6U_10U_1_o_mant_mux1h_1_itm[7:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_7_itm <= 2'b0;
    end
    else if ( (((mux_2098_nl) & (FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_3_0_1==4'b1111)
        & FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_4_1 & FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_5_1)
        | and_3689_cse | xnor_2_cse) & (cfg_precision_1_sva_st_81==2'b10) & and_dcpl_2185
        & nor_1877_cse ) begin
      reg_FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_7_itm <= FpMul_6U_10U_2_o_mant_mux1h_5_itm[9:8];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_7_1_itm <= 8'b0;
    end
    else if ( (((mux_2103_nl) & (FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_3_0_1==4'b1111)
        & FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_4_1 & FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_5_1)
        | and_3689_cse | xnor_2_cse | (chn_inp_in_crt_sva_4_739_736_1[2])) & (cfg_precision_1_sva_st_81[1])
        & main_stage_v_4 & core_wen & nor_1883_cse ) begin
      reg_FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_7_1_itm <= FpMul_6U_10U_2_o_mant_mux1h_5_itm[7:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_2_land_lpi_1_dfm_st_8 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_2_aelse_IsNaN_8U_23U_2_aelse_or_cse & (mux_510_nl)
        ) begin
      IsNaN_8U_23U_2_land_lpi_1_dfm_st_8 <= MUX_s_1_2_2(IsNaN_8U_23U_2_land_lpi_1_dfm_st_7,
          inp_lookup_4_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp, and_dcpl_679);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_int_mant_p1_sva_3 <= 50'b0;
    end
    else if ( core_wen & ((or_11_cse & (~ inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4))
        | and_1155_rgt) & (~ (mux_513_nl)) ) begin
      FpAdd_8U_23U_1_int_mant_p1_sva_3 <= MUX_v_50_2_2((inp_lookup_4_FpAdd_8U_23U_1_else_2_acc_nl),
          (inp_lookup_4_FpAdd_8U_23U_1_if_2_acc_nl), and_1155_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_6U_10U_2_o_mant_lpi_1_dfm_7_reg <= 2'b0;
    end
    else if ( or_11_cse & core_wen & (~ (chn_inp_in_crt_sva_4_739_736_1[3])) ) begin
      reg_FpMul_6U_10U_2_o_mant_lpi_1_dfm_7_reg <= FpMul_6U_10U_2_o_mant_FpMul_6U_10U_2_o_mant_mux_rgt[9:8];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_6U_10U_2_o_mant_lpi_1_dfm_7_1_reg <= 8'b0;
      reg_chn_inp_in_crt_sva_6_30_0_1_reg <= 23'b0;
      reg_chn_inp_in_crt_sva_6_62_32_1_reg <= 23'b0;
      reg_chn_inp_in_crt_sva_6_94_64_1_reg <= 23'b0;
      reg_chn_inp_in_crt_sva_6_126_96_1_reg <= 23'b0;
      reg_FpAdd_8U_23U_o_expo_1_lpi_1_dfm_11_1_reg <= 6'b0;
      reg_FpAdd_8U_23U_o_expo_2_lpi_1_dfm_11_1_reg <= 6'b0;
      reg_FpAdd_8U_23U_o_expo_3_lpi_1_dfm_11_1_reg <= 6'b0;
      reg_FpAdd_8U_23U_o_expo_lpi_1_dfm_11_1_reg <= 6'b0;
      reg_inp_lookup_1_else_else_a0_acc_2_reg <= 34'b0;
      reg_inp_lookup_2_else_else_a0_acc_2_reg <= 34'b0;
      reg_inp_lookup_3_else_else_a0_acc_2_reg <= 34'b0;
      reg_inp_lookup_4_else_else_a0_acc_2_reg <= 34'b0;
    end
    else if ( and_3483_cse ) begin
      reg_FpMul_6U_10U_2_o_mant_lpi_1_dfm_7_1_reg <= FpMul_6U_10U_2_o_mant_FpMul_6U_10U_2_o_mant_mux_rgt[7:0];
      reg_chn_inp_in_crt_sva_6_30_0_1_reg <= MUX1HOT_v_23_3_2(inp_lookup_1_FpAdd_6U_10U_1_a_int_mant_p1_lshift_itm,
          reg_chn_inp_in_crt_sva_5_30_0_1_itm, (FpAdd_8U_23U_1_int_mant_2_lpi_1_dfm_2_mx0[47:25]),
          {and_dcpl_691 , (or_6170_nl) , (and_1172_nl)});
      reg_chn_inp_in_crt_sva_6_62_32_1_reg <= MUX1HOT_v_23_3_2(inp_lookup_2_FpAdd_6U_10U_1_a_int_mant_p1_lshift_itm,
          reg_chn_inp_in_crt_sva_5_62_32_1_itm, (FpAdd_8U_23U_1_int_mant_3_lpi_1_dfm_2_mx0[47:25]),
          {and_dcpl_702 , (or_6171_nl) , (and_1183_nl)});
      reg_chn_inp_in_crt_sva_6_94_64_1_reg <= MUX1HOT_v_23_3_2(inp_lookup_3_FpAdd_6U_10U_1_a_int_mant_p1_lshift_itm,
          (FpAdd_8U_23U_1_int_mant_4_lpi_1_dfm_2_mx0[47:25]), reg_chn_inp_in_crt_sva_5_94_64_1_itm,
          {(nor_1910_nl) , (and_4169_nl) , mux_1903_tmp});
      reg_chn_inp_in_crt_sva_6_126_96_1_reg <= MUX1HOT_v_23_3_2(inp_lookup_4_FpAdd_6U_10U_1_a_int_mant_p1_lshift_itm,
          reg_chn_inp_in_crt_sva_5_126_96_1_itm, (FpAdd_8U_23U_1_int_mant_1_lpi_1_dfm_2_mx0[47:25]),
          {and_dcpl_720 , (or_6172_nl) , (and_1201_nl)});
      reg_FpAdd_8U_23U_o_expo_1_lpi_1_dfm_11_1_reg <= FpAdd_8U_23U_o_expo_FpAdd_8U_23U_o_expo_mux_rgt[5:0];
      reg_FpAdd_8U_23U_o_expo_2_lpi_1_dfm_11_1_reg <= FpAdd_8U_23U_o_expo_FpAdd_8U_23U_o_expo_mux_1_rgt[5:0];
      reg_FpAdd_8U_23U_o_expo_3_lpi_1_dfm_11_1_reg <= FpAdd_8U_23U_o_expo_FpAdd_8U_23U_o_expo_mux_2_rgt[5:0];
      reg_FpAdd_8U_23U_o_expo_lpi_1_dfm_11_1_reg <= FpAdd_8U_23U_o_expo_FpAdd_8U_23U_o_expo_mux_3_rgt[5:0];
      reg_inp_lookup_1_else_else_a0_acc_2_reg <= inp_lookup_else_else_a0_mux1h_rgt[33:0];
      reg_inp_lookup_2_else_else_a0_acc_2_reg <= inp_lookup_else_else_a0_mux1h_1_rgt[33:0];
      reg_inp_lookup_3_else_else_a0_acc_2_reg <= inp_lookup_else_else_a0_mux1h_2_rgt[33:0];
      reg_inp_lookup_4_else_else_a0_acc_2_reg <= inp_lookup_else_else_a0_mux1h_3_rgt[33:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_6 <= 1'b0;
    end
    else if ( core_wen & ((or_11_cse & main_stage_v_5) | main_stage_v_6_mx0c1) )
        begin
      main_stage_v_6 <= ~ main_stage_v_6_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_12 <= 8'b0;
    end
    else if ( core_wen & (and_dcpl_688 | and_1163_rgt) & (mux_515_nl) ) begin
      FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_12 <= MUX_v_8_2_2(FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_2_mx0w0,
          ({reg_FpAdd_8U_23U_o_expo_1_lpi_1_dfm_12_tmp , reg_FpAdd_8U_23U_o_expo_1_lpi_1_dfm_12_tmp_1}),
          and_1163_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_3_land_1_lpi_1_dfm_7 <= 1'b0;
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_itm_11 <= 1'b0;
      IsNaN_6U_10U_8_land_1_lpi_1_dfm_st_3 <= 1'b0;
      IsNaN_6U_10U_9_land_1_lpi_1_dfm_7 <= 1'b0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_18 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_3_aelse_and_cse ) begin
      IsNaN_8U_23U_3_land_1_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_1_lpi_1_dfm_6,
          inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5,
          and_dcpl_691);
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_itm_11 <= MUX_s_1_2_2(IsZero_6U_10U_1_IsZero_6U_10U_1_and_itm_10,
          inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6,
          and_dcpl_691);
      IsNaN_6U_10U_8_land_1_lpi_1_dfm_st_3 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_17,
          IsNaN_8U_23U_2_land_1_lpi_1_dfm_9, and_dcpl_690);
      IsNaN_6U_10U_9_land_1_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_6U_10U_9_land_1_lpi_1_dfm_6,
          IsNaN_8U_23U_2_land_1_lpi_1_dfm_st_7, and_dcpl_690);
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_18 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_17,
          IsNaN_6U_10U_8_land_1_lpi_1_dfm_6, and_dcpl_691);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_6_30_0_reg <= 8'b0;
    end
    else if ( or_11_cse & core_wen & (chn_inp_in_crt_sva_5_739_736_1[0]) & IsNaN_8U_23U_2_land_1_lpi_1_dfm_9
        ) begin
      reg_chn_inp_in_crt_sva_6_30_0_reg <= reg_chn_inp_in_crt_sva_5_30_0_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpMantRNE_49U_24U_1_else_and_svs_2 <= 1'b0;
      chn_inp_in_crt_sva_6_411_1 <= 1'b0;
      inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_12 <= 1'b0;
    end
    else if ( FpMantRNE_49U_24U_1_else_and_cse ) begin
      inp_lookup_1_FpMantRNE_49U_24U_1_else_and_svs_2 <= inp_lookup_1_FpMantRNE_49U_24U_1_else_and_tmp;
      chn_inp_in_crt_sva_6_411_1 <= chn_inp_in_crt_sva_5_411_1;
      inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_12 <= inp_lookup_1_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_st_83 <= 2'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_11_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_11_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_20 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_11_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_11_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_20 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_11_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_11_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_20 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_11_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_11_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_20 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_20 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_20 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_20 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_20 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_11_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_11_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_23 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_11_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_11_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_23 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_23 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_11_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_11_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_23 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_11_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_11_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_23 <= 4'b0;
      IsNaN_6U_10U_2_land_lpi_1_dfm_20 <= 1'b0;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_20 <= 1'b0;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_20 <= 1'b0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_20 <= 1'b0;
      inp_lookup_else_unequal_tmp_32 <= 1'b0;
      chn_inp_in_crt_sva_6_739_736_1 <= 4'b0;
    end
    else if ( cfg_precision_and_20_cse ) begin
      cfg_precision_1_sva_st_83 <= cfg_precision_1_sva_st_82;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_11_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_10_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_11_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_10_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_20 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_19;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_11_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_10_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_11_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_10_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_20 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_19;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_11_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_10_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_11_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_10_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_20 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_19;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_11_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_10_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_11_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_10_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_20 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_19;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_20 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_19;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_20 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_19;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_20 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_19;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_20 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_19;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_11_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_10_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_11_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_10_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_23 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_22;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_11_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_10_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_11_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_10_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_23 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_22;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_23 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_22;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_11_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_10_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_11_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_10_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_23 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_22;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_11_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_10_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_11_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_10_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_23 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_22;
      IsNaN_6U_10U_2_land_lpi_1_dfm_20 <= IsNaN_6U_10U_2_land_lpi_1_dfm_19;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_20 <= IsNaN_6U_10U_2_land_3_lpi_1_dfm_19;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_20 <= IsNaN_6U_10U_2_land_2_lpi_1_dfm_19;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_20 <= IsNaN_6U_10U_2_land_1_lpi_1_dfm_19;
      inp_lookup_else_unequal_tmp_32 <= ~((cfg_precision_1_sva_st_82==2'b10));
      chn_inp_in_crt_sva_6_739_736_1 <= chn_inp_in_crt_sva_5_739_736_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_b_int_mant_p1_1_sva_2 <= 23'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_521_nl) ) begin
      FpAdd_6U_10U_1_b_int_mant_p1_1_sva_2 <= inp_lookup_1_FpAdd_6U_10U_1_b_int_mant_p1_lshift_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_is_a_greater_lor_1_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_4_cse & (~
        (mux_526_nl)) ) begin
      FpAdd_6U_10U_1_is_a_greater_lor_1_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_6U_10U_1_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0,
          nor_126_cse, and_dcpl_690);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_13 <= 8'b0;
    end
    else if ( core_wen & (and_dcpl_699 | and_1174_rgt) & (mux_529_nl) ) begin
      FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_13 <= MUX_v_8_2_2(FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_2_mx0w0,
          ({reg_FpAdd_8U_23U_o_expo_2_lpi_1_dfm_12_tmp , reg_FpAdd_8U_23U_o_expo_2_lpi_1_dfm_12_tmp_1}),
          and_1174_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_3_land_2_lpi_1_dfm_7 <= 1'b0;
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_1_itm_9 <= 1'b0;
      IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_4 <= 1'b0;
      IsNaN_6U_10U_9_land_2_lpi_1_dfm_7 <= 1'b0;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_18 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_3_aelse_and_1_cse ) begin
      IsNaN_8U_23U_3_land_2_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_2_lpi_1_dfm_6,
          inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5,
          and_dcpl_702);
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_1_itm_9 <= MUX_s_1_2_2(IsZero_6U_10U_1_IsZero_6U_10U_1_and_1_itm_8,
          inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6,
          and_dcpl_702);
      IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_4 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_17,
          IsNaN_8U_23U_2_land_2_lpi_1_dfm_9, and_dcpl_701);
      IsNaN_6U_10U_9_land_2_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_6U_10U_9_land_2_lpi_1_dfm_6,
          IsNaN_8U_23U_2_land_2_lpi_1_dfm_st_7, and_dcpl_701);
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_18 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_17,
          IsNaN_6U_10U_8_land_2_lpi_1_dfm_4, and_dcpl_702);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_6_62_32_reg <= 8'b0;
    end
    else if ( or_11_cse & core_wen & (chn_inp_in_crt_sva_5_739_736_1[1]) & IsNaN_8U_23U_2_land_2_lpi_1_dfm_9
        ) begin
      reg_chn_inp_in_crt_sva_6_62_32_reg <= reg_chn_inp_in_crt_sva_5_62_32_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpMantRNE_49U_24U_1_else_and_svs_2 <= 1'b0;
      chn_inp_in_crt_sva_6_427_1 <= 1'b0;
      inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_11 <= 1'b0;
    end
    else if ( FpMantRNE_49U_24U_1_else_and_2_cse ) begin
      inp_lookup_2_FpMantRNE_49U_24U_1_else_and_svs_2 <= inp_lookup_2_FpMantRNE_49U_24U_1_else_and_tmp;
      chn_inp_in_crt_sva_6_427_1 <= chn_inp_in_crt_sva_5_427_1;
      inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_11 <= inp_lookup_2_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_b_int_mant_p1_2_sva_2 <= 23'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_534_nl) ) begin
      FpAdd_6U_10U_1_b_int_mant_p1_2_sva_2 <= inp_lookup_2_FpAdd_6U_10U_1_b_int_mant_p1_lshift_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_3_cse & (~
        (mux_539_nl)) ) begin
      FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0,
          FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_1_cse, and_dcpl_701);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_3_land_3_lpi_1_dfm_7 <= 1'b0;
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_itm_11 <= 1'b0;
      IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_4 <= 1'b0;
      IsNaN_6U_10U_9_land_3_lpi_1_dfm_7 <= 1'b0;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_18 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_3_aelse_and_2_cse ) begin
      IsNaN_8U_23U_3_land_3_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_3_lpi_1_dfm_6,
          inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5,
          and_dcpl_713);
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_itm_11 <= MUX_s_1_2_2(IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_itm_10,
          inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6,
          and_dcpl_713);
      IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_4 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_17,
          IsNaN_8U_23U_2_land_3_lpi_1_dfm_9, and_dcpl_712);
      IsNaN_6U_10U_9_land_3_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_6U_10U_9_land_3_lpi_1_dfm_6,
          IsNaN_8U_23U_2_land_3_lpi_1_dfm_st_7, and_dcpl_712);
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_18 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_17,
          IsNaN_6U_10U_8_land_3_lpi_1_dfm_4, and_dcpl_713);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_6_94_64_reg <= 8'b0;
    end
    else if ( or_11_cse & core_wen & (chn_inp_in_crt_sva_5_739_736_1[2]) & IsNaN_8U_23U_2_land_3_lpi_1_dfm_9
        ) begin
      reg_chn_inp_in_crt_sva_6_94_64_reg <= reg_chn_inp_in_crt_sva_5_94_64_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_inp_lookup_3_FpMantRNE_49U_24U_1_else_and_svs_1_cse <= 1'b0;
      chn_inp_in_crt_sva_6_443_1 <= 1'b0;
      inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_12 <= 1'b0;
    end
    else if ( FpMantRNE_49U_24U_1_else_and_4_cse ) begin
      reg_inp_lookup_3_FpMantRNE_49U_24U_1_else_and_svs_1_cse <= inp_lookup_3_FpMantRNE_49U_24U_1_else_and_tmp;
      chn_inp_in_crt_sva_6_443_1 <= chn_inp_in_crt_sva_5_443_1;
      inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_12 <= inp_lookup_3_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_b_int_mant_p1_3_sva_2 <= 23'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_544_nl) ) begin
      FpAdd_6U_10U_1_b_int_mant_p1_3_sva_2 <= inp_lookup_3_FpAdd_6U_10U_1_b_int_mant_p1_lshift_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_is_a_greater_lor_3_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_2_cse & (~
        (mux_547_nl)) ) begin
      FpAdd_6U_10U_1_is_a_greater_lor_3_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_6U_10U_1_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0,
          FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_2_cse, and_dcpl_712);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_o_expo_lpi_1_dfm_13 <= 8'b0;
    end
    else if ( core_wen & (and_dcpl_717 | and_1192_rgt) & (mux_550_nl) ) begin
      FpAdd_8U_23U_1_o_expo_lpi_1_dfm_13 <= MUX_v_8_2_2(FpAdd_8U_23U_1_o_expo_lpi_1_dfm_2_mx0w0,
          ({reg_FpAdd_8U_23U_o_expo_lpi_1_dfm_12_tmp , reg_FpAdd_8U_23U_o_expo_lpi_1_dfm_12_tmp_1}),
          and_1192_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_3_land_lpi_1_dfm_6 <= 1'b0;
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_3_itm_9 <= 1'b0;
      IsNaN_6U_10U_8_land_lpi_1_dfm_st_4 <= 1'b0;
      IsNaN_6U_10U_9_land_lpi_1_dfm_7 <= 1'b0;
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_17 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_3_aelse_and_3_cse ) begin
      IsNaN_8U_23U_3_land_lpi_1_dfm_6 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_lpi_1_dfm_5,
          inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5,
          and_dcpl_720);
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_3_itm_9 <= MUX_s_1_2_2(IsZero_6U_10U_1_IsZero_6U_10U_1_and_3_itm_8,
          inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5,
          and_dcpl_720);
      IsNaN_6U_10U_8_land_lpi_1_dfm_st_4 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_lpi_1_dfm_st_16,
          IsNaN_8U_23U_2_land_lpi_1_dfm_9, and_dcpl_719);
      IsNaN_6U_10U_9_land_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_6U_10U_9_land_lpi_1_dfm_6,
          IsNaN_8U_23U_2_land_lpi_1_dfm_st_8, and_dcpl_719);
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_17 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_lpi_1_dfm_st_16,
          IsNaN_6U_10U_8_land_lpi_1_dfm_4, and_dcpl_720);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_6_126_96_reg <= 8'b0;
    end
    else if ( or_11_cse & core_wen & (chn_inp_in_crt_sva_5_739_736_1[3]) & IsNaN_8U_23U_2_land_lpi_1_dfm_9
        ) begin
      reg_chn_inp_in_crt_sva_6_126_96_reg <= reg_chn_inp_in_crt_sva_5_126_96_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpMantRNE_49U_24U_1_else_and_svs_2 <= 1'b0;
      chn_inp_in_crt_sva_6_459_1 <= 1'b0;
      inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_12 <= 1'b0;
    end
    else if ( FpMantRNE_49U_24U_1_else_and_6_cse ) begin
      inp_lookup_4_FpMantRNE_49U_24U_1_else_and_svs_2 <= inp_lookup_4_FpMantRNE_49U_24U_1_else_and_tmp;
      chn_inp_in_crt_sva_6_459_1 <= chn_inp_in_crt_sva_5_459_1;
      inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_12 <= inp_lookup_4_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_b_int_mant_p1_sva_2 <= 23'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_555_nl) ) begin
      FpAdd_6U_10U_1_b_int_mant_p1_sva_2 <= inp_lookup_4_FpAdd_6U_10U_1_b_int_mant_p1_lshift_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_is_a_greater_lor_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_3_aelse_IsNaN_8U_23U_3_aelse_or_1_cse & (~
        (mux_558_nl)) ) begin
      FpAdd_6U_10U_1_is_a_greater_lor_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_6U_10U_1_is_a_greater_lor_lpi_1_dfm_1_mx0w0,
          nor_136_cse, and_dcpl_719);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_7 <= 1'b0;
    end
    else if ( core_wen & ((or_11_cse & main_stage_v_6) | main_stage_v_7_mx0c1) )
        begin
      main_stage_v_7 <= ~ main_stage_v_7_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_2
          <= 1'b0;
      inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2
          <= 1'b0;
      inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_13 <= 1'b0;
    end
    else if ( FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_and_cse ) begin
      inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_2
          <= inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8;
      inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2
          <= inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8;
      inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_13 <= inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_12;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpMantRNE_24U_11U_else_and_svs_2 <= 1'b0;
    end
    else if ( core_wen & ((inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8
        & (~ inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7) & inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8
        & or_11_cse) | and_1209_rgt) & (~ mux_559_itm) ) begin
      inp_lookup_1_FpMantRNE_24U_11U_else_and_svs_2 <= MUX_s_1_2_2(inp_lookup_1_FpMantRNE_24U_11U_else_and_svs_mx0w0,
          inp_lookup_1_FpMantRNE_24U_11U_else_and_svs, and_1209_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((or_11_cse & IsNaN_6U_10U_8_land_1_lpi_1_dfm_st_3) | and_1211_rgt)
        & (mux_562_nl) ) begin
      FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_6 <= MUX_v_23_2_2(reg_chn_inp_in_crt_sva_6_30_0_1_reg,
          FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_4_itm, and_4221_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_1_sva_2 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_563_nl) ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_1_sva_2 <= nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_1_sva_2[4:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_565_nl) ) begin
      inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2
          <= inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2
          <= 1'b0;
    end
    else if ( core_wen & ((or_11_cse & inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8)
        | and_1213_rgt) & (~ mux_559_itm) ) begin
      inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2
          <= MUX_s_1_2_2(inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7,
          inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs,
          and_1213_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_st_84 <= 2'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_12_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_12_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_21 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_12_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_12_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_21 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_12_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_12_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_21 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_12_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_12_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_21 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_21 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_21 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_21 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_21 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_12_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_12_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_24 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_12_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_12_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_24 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_24 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_12_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_12_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_24 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_12_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_12_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_24 <= 4'b0;
      IsNaN_6U_10U_2_land_lpi_1_dfm_21 <= 1'b0;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_21 <= 1'b0;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_21 <= 1'b0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_21 <= 1'b0;
      inp_lookup_else_unequal_tmp_33 <= 1'b0;
      chn_inp_in_crt_sva_7_739_736_1 <= 4'b0;
    end
    else if ( cfg_precision_and_24_cse ) begin
      cfg_precision_1_sva_st_84 <= cfg_precision_1_sva_st_83;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_12_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_11_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_12_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_11_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_21 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_20;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_12_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_11_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_12_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_11_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_21 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_20;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_12_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_11_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_12_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_11_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_21 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_20;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_12_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_11_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_12_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_11_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_21 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_20;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_21 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_20;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_21 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_20;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_21 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_20;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_21 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_20;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_12_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_11_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_12_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_11_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_24 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_23;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_12_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_11_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_12_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_11_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_24 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_23;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_24 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_23;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_12_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_11_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_12_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_11_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_24 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_23;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_12_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_11_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_12_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_11_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_24 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_23;
      IsNaN_6U_10U_2_land_lpi_1_dfm_21 <= IsNaN_6U_10U_2_land_lpi_1_dfm_20;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_21 <= IsNaN_6U_10U_2_land_3_lpi_1_dfm_20;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_21 <= IsNaN_6U_10U_2_land_2_lpi_1_dfm_20;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_21 <= IsNaN_6U_10U_2_land_1_lpi_1_dfm_20;
      inp_lookup_else_unequal_tmp_33 <= inp_lookup_else_unequal_tmp_32;
      chn_inp_in_crt_sva_7_739_736_1 <= chn_inp_in_crt_sva_6_739_736_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_2_lpi_1_dfm_5 <= 6'b0;
    end
    else if ( core_wen & (and_dcpl_740 | FpAdd_6U_10U_1_and_47_rgt | (or_4591_tmp
        & and_dcpl_741)) & (mux_569_nl) ) begin
      FpAdd_6U_10U_1_qr_2_lpi_1_dfm_5 <= MUX_v_6_2_2(({FpAdd_6U_10U_1_qr_2_lpi_1_dfm_3_5_1
          , FpAdd_6U_10U_1_qr_2_lpi_1_dfm_3_4_1 , FpAdd_6U_10U_1_qr_2_lpi_1_dfm_3_3_0_1}),
          (FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_7_mx0w0[5:0]), FpAdd_6U_10U_1_and_47_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_4 <= 24'b0;
    end
    else if ( core_wen & ((or_11_cse & IsNaN_8U_23U_3_land_1_lpi_1_dfm_7) | and_1217_rgt)
        & (~ (mux_570_nl)) ) begin
      FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_4 <= MUX_v_24_2_2(FpAdd_6U_10U_1_int_mant_p1_1_sva,
          FpAdd_6U_10U_1_int_mant_p1_1_sva_1, and_1217_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_6U_23U_1_if_or_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpNormalize_6U_23U_1_if_FpNormalize_6U_23U_1_if_or_3_cse
        & (~ (mux_572_nl)) ) begin
      FpNormalize_6U_23U_1_if_or_itm_2 <= MUX_s_1_2_2((FpNormalize_6U_23U_1_if_or_nl),
          IsZero_6U_10U_1_IsZero_6U_10U_1_and_itm_11, and_dcpl_741);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpMantRNE_24U_11U_else_and_svs_2 <= 1'b0;
    end
    else if ( core_wen & ((inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8
        & (~ inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7) & inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8
        & or_11_cse) | and_1221_rgt) & (~ mux_573_itm) ) begin
      inp_lookup_2_FpMantRNE_24U_11U_else_and_svs_2 <= MUX_s_1_2_2(inp_lookup_2_FpMantRNE_24U_11U_else_and_svs_mx0w0,
          inp_lookup_2_FpMantRNE_24U_11U_else_and_svs, and_1221_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((or_11_cse & IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_4) | and_1223_rgt)
        & (mux_575_nl) ) begin
      FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_6 <= MUX_v_23_2_2(reg_chn_inp_in_crt_sva_6_62_32_1_reg,
          FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_5_itm, and_4220_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_2_sva_2 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_576_nl) ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_2_sva_2 <= nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_2_sva_2[4:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_578_nl) ) begin
      inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2
          <= inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2
          <= 1'b0;
    end
    else if ( core_wen & ((or_11_cse & inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8)
        | and_1225_rgt) & (~ mux_573_itm) ) begin
      inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2
          <= MUX_s_1_2_2(inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7,
          inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs,
          and_1225_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2
          <= 1'b0;
      inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_12 <= 1'b0;
    end
    else if ( FpWidthDec_8U_23U_6U_10U_0U_1U_if_and_2_cse ) begin
      inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2
          <= inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8;
      inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_12 <= inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_11;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_3_lpi_1_dfm_5 <= 6'b0;
    end
    else if ( core_wen & FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_14_cse & (mux_581_nl) )
        begin
      FpAdd_6U_10U_1_qr_3_lpi_1_dfm_5 <= MUX_v_6_2_2(({FpAdd_6U_10U_1_qr_3_lpi_1_dfm_3_5_1
          , FpAdd_6U_10U_1_qr_3_lpi_1_dfm_3_4_1 , FpAdd_6U_10U_1_qr_3_lpi_1_dfm_3_3_0_1}),
          (FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_7[5:0]), and_dcpl_753);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_4 <= 24'b0;
    end
    else if ( core_wen & ((or_11_cse & IsNaN_8U_23U_3_land_2_lpi_1_dfm_7) | and_1229_rgt)
        & (~ (mux_582_nl)) ) begin
      FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_4 <= MUX_v_24_2_2(FpAdd_6U_10U_1_int_mant_p1_2_sva,
          FpAdd_6U_10U_1_int_mant_p1_2_sva_1, and_1229_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_6U_23U_1_if_or_1_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_14_cse & (~ (mux_585_nl))
        ) begin
      FpNormalize_6U_23U_1_if_or_1_itm_2 <= MUX_s_1_2_2((FpNormalize_6U_23U_1_if_or_1_nl),
          IsZero_6U_10U_1_IsZero_6U_10U_1_and_1_itm_9, and_dcpl_753);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_5 <= 1'b0;
      IsNaN_6U_10U_9_land_2_lpi_1_dfm_8 <= 1'b0;
      chn_inp_in_crt_sva_7_427_1 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_8_aelse_and_cse ) begin
      IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_5 <= MUX_s_1_2_2(IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_4,
          IsNaN_8U_23U_4_IsNaN_8U_23U_4_nor_1_tmp, and_dcpl_753);
      IsNaN_6U_10U_9_land_2_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_6U_10U_9_land_2_lpi_1_dfm_7,
          inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8, and_dcpl_753);
      chn_inp_in_crt_sva_7_427_1 <= MUX_s_1_2_2(chn_inp_in_crt_sva_6_427_1, (FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_mx0[23]),
          and_dcpl_752);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpMantRNE_24U_11U_else_and_svs_2 <= 1'b0;
    end
    else if ( core_wen & ((inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8
        & (~ inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7) & inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8
        & or_11_cse) | and_1233_rgt) & (~ mux_587_itm) ) begin
      inp_lookup_3_FpMantRNE_24U_11U_else_and_svs_2 <= MUX_s_1_2_2(inp_lookup_3_FpMantRNE_24U_11U_else_and_svs_mx0w0,
          inp_lookup_3_FpMantRNE_24U_11U_else_and_svs, and_1233_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((or_11_cse & IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_4) | and_1235_rgt)
        & (mux_590_nl) ) begin
      FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_6 <= MUX_v_23_2_2(reg_chn_inp_in_crt_sva_6_94_64_1_reg,
          FpAdd_8U_23U_1_asn_40_mx0w1, and_1235_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_592_nl) ) begin
      inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2
          <= inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2
          <= 1'b0;
    end
    else if ( core_wen & ((or_11_cse & inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8)
        | and_1237_rgt) & (~ mux_587_itm) ) begin
      inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2
          <= MUX_s_1_2_2(inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7,
          inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs,
          and_1237_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2
          <= 1'b0;
      inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_13 <= 1'b0;
    end
    else if ( FpWidthDec_8U_23U_6U_10U_0U_1U_if_and_4_cse ) begin
      inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2
          <= inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8;
      inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_13 <= inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_12;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_4_lpi_1_dfm_5 <= 6'b0;
    end
    else if ( core_wen & FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_13_cse & (~ (mux_595_nl))
        ) begin
      FpAdd_6U_10U_1_qr_4_lpi_1_dfm_5 <= MUX_v_6_2_2(({FpAdd_6U_10U_1_qr_4_lpi_1_dfm_3_5_1
          , FpAdd_6U_10U_1_qr_4_lpi_1_dfm_3_4_1 , FpAdd_6U_10U_1_qr_4_lpi_1_dfm_3_3_0_1}),
          (FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_7[5:0]), and_dcpl_765);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_4 <= 24'b0;
    end
    else if ( core_wen & ((or_11_cse & IsNaN_8U_23U_3_land_3_lpi_1_dfm_7) | and_1241_rgt)
        & (~ (mux_596_nl)) ) begin
      FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_4 <= MUX_v_24_2_2(FpAdd_6U_10U_1_int_mant_p1_3_sva,
          FpAdd_6U_10U_1_int_mant_p1_3_sva_1, and_1241_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_6U_23U_1_if_or_2_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_13_cse & (mux_597_nl) )
        begin
      FpNormalize_6U_23U_1_if_or_2_itm_2 <= MUX_s_1_2_2((FpNormalize_6U_23U_1_if_or_2_nl),
          IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_itm_11, and_dcpl_765);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_5 <= 1'b0;
      IsNaN_6U_10U_9_land_3_lpi_1_dfm_8 <= 1'b0;
      chn_inp_in_crt_sva_7_443_1 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_8_aelse_and_1_cse ) begin
      IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_5 <= MUX_s_1_2_2(IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_4,
          IsNaN_8U_23U_4_IsNaN_8U_23U_4_nor_2_tmp, and_dcpl_765);
      IsNaN_6U_10U_9_land_3_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_6U_10U_9_land_3_lpi_1_dfm_7,
          inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8, and_dcpl_765);
      chn_inp_in_crt_sva_7_443_1 <= MUX_s_1_2_2(chn_inp_in_crt_sva_6_443_1, (FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_mx0[23]),
          and_dcpl_764);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpMantRNE_24U_11U_else_and_svs_2 <= 1'b0;
    end
    else if ( core_wen & ((inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8
        & (~ inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7) & inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8
        & or_11_cse) | and_1245_rgt) & (~ mux_599_itm) ) begin
      inp_lookup_4_FpMantRNE_24U_11U_else_and_svs_2 <= MUX_s_1_2_2(inp_lookup_4_FpMantRNE_24U_11U_else_and_svs_mx0w0,
          inp_lookup_4_FpMantRNE_24U_11U_else_and_svs, and_1245_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_o_mant_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((or_11_cse & IsNaN_6U_10U_8_land_lpi_1_dfm_st_4) | and_1247_rgt)
        & (mux_601_nl) ) begin
      FpAdd_8U_23U_1_o_mant_lpi_1_dfm_6 <= MUX_v_23_2_2(reg_chn_inp_in_crt_sva_6_126_96_1_reg,
          FpAdd_8U_23U_1_FpAdd_8U_23U_1_or_7_itm, and_4219_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva_2 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_602_nl) ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva_2 <= nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva_2[4:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_604_nl) ) begin
      inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2
          <= inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2
          <= 1'b0;
    end
    else if ( core_wen & ((or_11_cse & inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8)
        | and_1249_rgt) & (~ mux_599_itm) ) begin
      inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2
          <= MUX_s_1_2_2(inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7,
          inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs,
          and_1249_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2
          <= 1'b0;
      inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_13 <= 1'b0;
    end
    else if ( FpWidthDec_8U_23U_6U_10U_0U_1U_if_and_6_cse ) begin
      inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2
          <= inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8;
      inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_13 <= inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_12;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_lpi_1_dfm_5 <= 6'b0;
    end
    else if ( core_wen & FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_12_cse & (~ (mux_609_nl))
        ) begin
      FpAdd_6U_10U_1_qr_lpi_1_dfm_5 <= MUX_v_6_2_2(({FpAdd_6U_10U_1_qr_lpi_1_dfm_3_5_1
          , FpAdd_6U_10U_1_qr_lpi_1_dfm_3_4_1 , FpAdd_6U_10U_1_qr_lpi_1_dfm_3_3_0_1}),
          (FpAdd_8U_23U_1_o_expo_lpi_1_dfm_7[5:0]), and_dcpl_777);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_4 <= 24'b0;
    end
    else if ( core_wen & ((or_11_cse & IsNaN_8U_23U_3_land_lpi_1_dfm_6) | and_1253_rgt)
        & (~ (mux_610_nl)) ) begin
      FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_4 <= MUX_v_24_2_2(FpAdd_6U_10U_1_int_mant_p1_sva,
          FpAdd_6U_10U_1_int_mant_p1_sva_1, and_1253_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_6U_23U_1_if_or_3_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_12_cse & (mux_611_nl) )
        begin
      FpNormalize_6U_23U_1_if_or_3_itm_2 <= MUX_s_1_2_2((FpNormalize_6U_23U_1_if_or_3_nl),
          IsZero_6U_10U_1_IsZero_6U_10U_1_and_3_itm_9, and_dcpl_777);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_8_land_lpi_1_dfm_st_5 <= 1'b0;
      IsNaN_6U_10U_9_land_lpi_1_dfm_8 <= 1'b0;
      chn_inp_in_crt_sva_7_459_1 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_8_aelse_and_2_cse ) begin
      IsNaN_6U_10U_8_land_lpi_1_dfm_st_5 <= MUX_s_1_2_2(IsNaN_6U_10U_8_land_lpi_1_dfm_st_4,
          IsNaN_8U_23U_4_IsNaN_8U_23U_4_nor_3_tmp, and_dcpl_777);
      IsNaN_6U_10U_9_land_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_6U_10U_9_land_lpi_1_dfm_7,
          inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8, and_dcpl_777);
      chn_inp_in_crt_sva_7_459_1 <= MUX_s_1_2_2(chn_inp_in_crt_sva_6_459_1, (FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_mx0[23]),
          and_dcpl_776);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_8 <= 1'b0;
    end
    else if ( core_wen & ((or_11_cse & main_stage_v_7) | main_stage_v_8_mx0c1) )
        begin
      main_stage_v_8 <= ~ main_stage_v_8_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_10_5_1 <= 1'b0;
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_10_4_0_1 <= 5'b0;
    end
    else if ( FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_and_cse ) begin
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_10_5_1 <= FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_7_5_mx0w0;
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_10_4_0_1 <= FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_7_4_0_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_13_1_1 <= 1'b0;
      FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_5_1 <= 1'b0;
      FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_3_0_1 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_12_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_13_1_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_12_1_1,
          (inp_lookup_1_IsInf_6U_23U_1_IsInf_6U_23U_1_and_nl), and_dcpl_785);
      FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_5_1 <= MUX_s_1_2_2(FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_5_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_12_0_1, and_dcpl_784);
      FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_3_0_1 <= MUX_v_4_2_2(FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_3_0_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_21, and_dcpl_784);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_oelse_1_acc_itm_2 <= 7'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_620_nl) ) begin
      FpMul_6U_10U_oelse_1_acc_itm_2 <= z_out_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_6U_10U_lor_3_lpi_1_dfm_3_cse <= 1'b0;
      inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_14 <= 1'b0;
    end
    else if ( FpMul_6U_10U_oelse_and_cse ) begin
      reg_FpMul_6U_10U_lor_3_lpi_1_dfm_3_cse <= FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_tmp;
      inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_14 <= inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_13;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_st_85 <= 2'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_13_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_13_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_25 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_13_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_13_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_25 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_25 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_13_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_13_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_25 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_13_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_13_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_25 <= 4'b0;
      inp_lookup_else_unequal_tmp_55 <= 1'b0;
      IsNaN_6U_10U_2_land_lpi_1_dfm_22 <= 1'b0;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_22 <= 1'b0;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_22 <= 1'b0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_22 <= 1'b0;
      chn_inp_in_crt_sva_8_739_736_1 <= 4'b0;
    end
    else if ( cfg_precision_and_28_cse ) begin
      cfg_precision_1_sva_st_85 <= cfg_precision_1_sva_st_84;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_13_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_12_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_13_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_12_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_25 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_24;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_13_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_12_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_13_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_12_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_25 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_24;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_25 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_24;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_13_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_12_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_13_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_12_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_25 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_24;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_13_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_12_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_13_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_12_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_25 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_24;
      inp_lookup_else_unequal_tmp_55 <= inp_lookup_else_unequal_tmp_33;
      IsNaN_6U_10U_2_land_lpi_1_dfm_22 <= IsNaN_6U_10U_2_land_lpi_1_dfm_21;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_22 <= IsNaN_6U_10U_2_land_3_lpi_1_dfm_21;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_22 <= IsNaN_6U_10U_2_land_2_lpi_1_dfm_21;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_22 <= IsNaN_6U_10U_2_land_1_lpi_1_dfm_21;
      chn_inp_in_crt_sva_8_739_736_1 <= chn_inp_in_crt_sva_7_739_736_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_4_1 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_785 | and_dcpl_787 | and_1270_rgt | and_1273_rgt)
        & (~ mux_623_itm) ) begin
      FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_4_1 <= MUX1HOT_s_1_4_2(FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_4_mx0w0,
          FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_8_4_1, chn_inp_in_crt_sva_7_411_1, (inp_lookup_1_FpMul_6U_10U_xor_1_nl),
          {and_dcpl_785 , and_dcpl_787 , and_1270_rgt , and_1273_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_itm_2 <= 10'b0;
    end
    else if ( core_wen & (and_1277_rgt | and_1279_rgt | and_1280_rgt) & (~ mux_623_itm)
        ) begin
      FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_itm_2 <= MUX1HOT_v_10_3_2(FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_itm_mx0w0,
          FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_itm, FpMul_6U_10U_1_o_mant_1_lpi_1_dfm_11,
          {and_1277_rgt , and_1279_rgt , and_1280_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_10_5_1 <= 1'b0;
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_10_4_0_1 <= 5'b0;
    end
    else if ( FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_and_2_cse ) begin
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_10_5_1 <= FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_7_5_mx0w0;
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_10_4_0_1 <= FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_7_4_0_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_13_1_1 <= 1'b0;
      FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_5_1 <= 1'b0;
      FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_3_0_1 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_13_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_13_1_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_12_1_1,
          (inp_lookup_2_IsInf_6U_23U_1_IsInf_6U_23U_1_and_nl), and_dcpl_808);
      FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_5_1 <= MUX_s_1_2_2(FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_5_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_12_0_1, and_dcpl_807);
      FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_3_0_1 <= MUX_v_4_2_2(FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_3_0_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_21, and_dcpl_807);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_oelse_1_acc_1_itm_2 <= 7'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_630_nl) ) begin
      FpMul_6U_10U_oelse_1_acc_1_itm_2 <= z_out_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_6U_10U_lor_4_lpi_1_dfm_3_cse <= 1'b0;
      inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_13 <= 1'b0;
    end
    else if ( FpMul_6U_10U_oelse_and_2_cse ) begin
      reg_FpMul_6U_10U_lor_4_lpi_1_dfm_3_cse <= FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_2_tmp;
      inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_13 <= inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_12;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_4_1 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_808 | and_dcpl_810 | and_1293_rgt | and_1296_rgt)
        & (~ mux_632_itm) ) begin
      FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_4_1 <= MUX1HOT_s_1_4_2(FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_4_mx0w0,
          FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_8_4_1, chn_inp_in_crt_sva_7_427_1, (inp_lookup_2_FpMul_6U_10U_xor_1_nl),
          {and_dcpl_808 , and_dcpl_810 , and_1293_rgt , and_1296_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_1_itm_2 <= 10'b0;
    end
    else if ( core_wen & (nor_1733_rgt | and_1303_rgt | and_1304_rgt) & (~ mux_632_itm)
        ) begin
      FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_1_itm_2 <= MUX1HOT_v_10_3_2(FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_1_itm_mx0w0,
          FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_1_itm, FpMul_6U_10U_1_o_mant_2_lpi_1_dfm_11,
          {nor_1733_rgt , and_1303_rgt , and_1304_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_10_5_1 <= 1'b0;
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_10_4_0_1 <= 5'b0;
    end
    else if ( FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_and_4_cse ) begin
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_10_5_1 <= FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_7_5_mx0w0;
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_10_4_0_1 <= FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_7_4_0_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_13_1_1 <= 1'b0;
      FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_5_1 <= 1'b0;
      FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_3_0_1 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_14_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_13_1_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_12_1_1,
          (inp_lookup_3_IsInf_6U_23U_1_IsInf_6U_23U_1_and_nl), and_dcpl_832);
      FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_5_1 <= MUX_s_1_2_2(FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_5_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_12_0_1, and_dcpl_831);
      FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_3_0_1 <= MUX_v_4_2_2(FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_3_0_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_21, and_dcpl_831);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_oelse_1_acc_2_itm_2 <= 7'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_640_nl) ) begin
      FpMul_6U_10U_oelse_1_acc_2_itm_2 <= z_out_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_6U_10U_lor_5_lpi_1_dfm_3_cse <= 1'b0;
      inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_14 <= 1'b0;
    end
    else if ( FpMul_6U_10U_oelse_and_4_cse ) begin
      reg_FpMul_6U_10U_lor_5_lpi_1_dfm_3_cse <= FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_4_tmp;
      inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_14 <= inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_13;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_4_1 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_832 | and_dcpl_834 | and_1317_rgt | and_1320_rgt)
        & (~ mux_623_itm) ) begin
      FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_4_1 <= MUX1HOT_s_1_4_2(FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_4_mx0w0,
          FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_8_4_1, chn_inp_in_crt_sva_7_443_1, (inp_lookup_3_FpMul_6U_10U_xor_1_nl),
          {and_dcpl_832 , and_dcpl_834 , and_1317_rgt , and_1320_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_2_itm_2 <= 10'b0;
    end
    else if ( core_wen & (nor_1732_rgt | and_1327_rgt | and_dcpl_831 | and_1329_rgt)
        & not_tmp_546 ) begin
      FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_2_itm_2 <= MUX1HOT_v_10_4_2(FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_2_itm_mx0w0,
          FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_2_itm, FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_21,
          ({reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_8_itm_4_3 , reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_8_itm_2_0
          , reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_8_1_itm}), {nor_1732_rgt , and_1327_rgt
          , and_dcpl_831 , and_1329_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_10_5_1 <= 1'b0;
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_10_4_0_1 <= 5'b0;
    end
    else if ( FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_and_6_cse ) begin
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_10_5_1 <= FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_7_5_mx0w0;
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_10_4_0_1 <= FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_7_4_0_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_13_1_1 <= 1'b0;
      FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_5_1 <= 1'b0;
      FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_3_0_1 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_15_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_13_1_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_12_1_1,
          (inp_lookup_4_IsInf_6U_23U_1_IsInf_6U_23U_1_and_nl), and_dcpl_857);
      FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_5_1 <= MUX_s_1_2_2(FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_5_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_12_0_1, and_dcpl_856);
      FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_3_0_1 <= MUX_v_4_2_2(FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_3_0_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_21, and_dcpl_856);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_oelse_1_acc_3_itm_2 <= 7'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_650_nl) ) begin
      FpMul_6U_10U_oelse_1_acc_3_itm_2 <= z_out_11;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_6U_10U_lor_lpi_1_dfm_3_cse <= 1'b0;
      inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_14 <= 1'b0;
    end
    else if ( FpMul_6U_10U_oelse_and_6_cse ) begin
      reg_FpMul_6U_10U_lor_lpi_1_dfm_3_cse <= FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_6_tmp;
      inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_14 <= inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_13;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_4_1 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_857 | and_dcpl_859 | and_1342_rgt | and_1345_rgt)
        & (~ mux_623_itm) ) begin
      FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_4_1 <= MUX1HOT_s_1_4_2(FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_4_mx0w0,
          FpMul_6U_10U_1_o_expo_lpi_1_dfm_8_4_1, chn_inp_in_crt_sva_7_459_1, (inp_lookup_4_FpMul_6U_10U_xor_1_nl),
          {and_dcpl_857 , and_dcpl_859 , and_1342_rgt , and_1345_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_3_itm_2 <= 10'b0;
    end
    else if ( core_wen & (and_1349_rgt | and_1351_rgt | and_1352_rgt) & (~ mux_623_itm)
        ) begin
      FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_3_itm_2 <= MUX1HOT_v_10_3_2(FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_3_itm_mx0w0,
          FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_3_itm, FpMul_6U_10U_1_o_mant_lpi_1_dfm_10,
          {and_1349_rgt , and_1351_rgt , and_1352_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_9 <= 1'b0;
    end
    else if ( core_wen & ((or_11_cse & main_stage_v_8) | main_stage_v_9_mx0c1) )
        begin
      main_stage_v_9 <= ~ main_stage_v_9_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_else_2_else_ac_int_cctor_1_sva_2 <= 6'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_654_nl) ) begin
      FpMul_6U_10U_else_2_else_ac_int_cctor_1_sva_2 <= nl_FpMul_6U_10U_else_2_else_ac_int_cctor_1_sva_2[5:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpMul_6U_10U_else_2_else_slc_FpMul_6U_10U_p_mant_p1_21_itm_2 <=
          1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_656_nl) ) begin
      inp_lookup_1_FpMul_6U_10U_else_2_else_slc_FpMul_6U_10U_p_mant_p1_21_itm_2 <=
          inp_lookup_1_FpMul_6U_10U_p_mant_p1_mul_tmp[21];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_21 <= 1'b0;
      FpMul_6U_10U_lor_6_lpi_1_dfm_st_2 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_23 <= 10'b0;
      IsNaN_6U_10U_land_1_lpi_1_dfm_6 <= 1'b0;
      IsNaN_6U_10U_1_land_1_lpi_1_dfm_6 <= 1'b0;
      inp_lookup_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_4 <=
          1'b0;
    end
    else if ( IsNaN_6U_10U_2_aelse_and_cse ) begin
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_21 <= IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_20;
      FpMul_6U_10U_lor_6_lpi_1_dfm_st_2 <= or_5020_cse;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_23 <= FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_itm_2;
      IsNaN_6U_10U_land_1_lpi_1_dfm_6 <= IsNaN_6U_10U_land_1_lpi_1_dfm_5;
      IsNaN_6U_10U_1_land_1_lpi_1_dfm_6 <= IsNaN_6U_10U_1_land_1_lpi_1_dfm_5;
      inp_lookup_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_4 <=
          ~(chn_inp_in_crt_sva_8_283_1 ^ FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_4_1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_p_mant_p1_1_sva_2 <= 22'b0;
    end
    else if ( core_wen & (((~ inp_lookup_1_FpMul_6U_10U_oelse_1_acc_itm_7_1) & (~
        reg_FpMul_6U_10U_lor_3_lpi_1_dfm_3_cse) & or_11_cse & inp_lookup_1_FpMul_6U_10U_else_2_if_acc_itm_6_1)
        | and_1360_rgt) & (~ mux_659_itm) ) begin
      FpMul_6U_10U_p_mant_p1_1_sva_2 <= MUX_v_22_2_2(inp_lookup_1_FpMul_6U_10U_p_mant_p1_mul_tmp,
          FpMul_6U_10U_p_mant_p1_1_sva, and_1360_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_st_86 <= 2'b0;
      chn_inp_in_crt_sva_9_283_1 <= 1'b0;
    end
    else if ( cfg_precision_and_32_cse ) begin
      cfg_precision_1_sva_st_86 <= cfg_precision_1_sva_st_85;
      chn_inp_in_crt_sva_9_283_1 <= chn_inp_in_crt_sva_8_283_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_else_2_else_ac_int_cctor_2_sva_2 <= 6'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_662_nl) ) begin
      FpMul_6U_10U_else_2_else_ac_int_cctor_2_sva_2 <= nl_FpMul_6U_10U_else_2_else_ac_int_cctor_2_sva_2[5:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpMul_6U_10U_else_2_else_slc_FpMul_6U_10U_p_mant_p1_21_itm_2 <=
          1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_664_nl) ) begin
      inp_lookup_2_FpMul_6U_10U_else_2_else_slc_FpMul_6U_10U_p_mant_p1_21_itm_2 <=
          inp_lookup_2_FpMul_6U_10U_p_mant_p1_mul_tmp[21];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_21 <= 1'b0;
      FpMul_6U_10U_lor_7_lpi_1_dfm_st_2 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_23 <= 10'b0;
      IsNaN_6U_10U_land_2_lpi_1_dfm_6 <= 1'b0;
      IsNaN_6U_10U_1_land_2_lpi_1_dfm_6 <= 1'b0;
      inp_lookup_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_4 <=
          1'b0;
    end
    else if ( IsNaN_6U_10U_2_aelse_and_1_cse ) begin
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_21 <= IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_20;
      FpMul_6U_10U_lor_7_lpi_1_dfm_st_2 <= or_5021_cse;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_23 <= FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_1_itm_2;
      IsNaN_6U_10U_land_2_lpi_1_dfm_6 <= IsNaN_6U_10U_land_2_lpi_1_dfm_5;
      IsNaN_6U_10U_1_land_2_lpi_1_dfm_6 <= IsNaN_6U_10U_1_land_2_lpi_1_dfm_5;
      inp_lookup_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_4 <=
          ~(chn_inp_in_crt_sva_8_299_1 ^ FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_4_1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_p_mant_p1_2_sva_2 <= 22'b0;
    end
    else if ( core_wen & (((~ inp_lookup_2_FpMul_6U_10U_oelse_1_acc_itm_7_1) & (~
        reg_FpMul_6U_10U_lor_4_lpi_1_dfm_3_cse) & or_11_cse & inp_lookup_2_FpMul_6U_10U_else_2_if_acc_itm_6_1)
        | and_1364_rgt) & (~ mux_666_itm) ) begin
      FpMul_6U_10U_p_mant_p1_2_sva_2 <= MUX_v_22_2_2(inp_lookup_2_FpMul_6U_10U_p_mant_p1_mul_tmp,
          FpMul_6U_10U_p_mant_p1_2_sva, and_1364_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_st_100 <= 2'b0;
      chn_inp_in_crt_sva_9_299_1 <= 1'b0;
    end
    else if ( cfg_precision_and_33_cse ) begin
      cfg_precision_1_sva_st_100 <= cfg_precision_1_sva_st_85;
      chn_inp_in_crt_sva_9_299_1 <= chn_inp_in_crt_sva_8_299_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_else_2_else_ac_int_cctor_3_sva_2 <= 6'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_669_nl) ) begin
      FpMul_6U_10U_else_2_else_ac_int_cctor_3_sva_2 <= nl_FpMul_6U_10U_else_2_else_ac_int_cctor_3_sva_2[5:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpMul_6U_10U_else_2_else_slc_FpMul_6U_10U_p_mant_p1_21_itm_2 <=
          1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_671_nl) ) begin
      inp_lookup_3_FpMul_6U_10U_else_2_else_slc_FpMul_6U_10U_p_mant_p1_21_itm_2 <=
          inp_lookup_3_FpMul_6U_10U_p_mant_p1_mul_tmp[21];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_21 <= 1'b0;
      FpMul_6U_10U_lor_8_lpi_1_dfm_st_2 <= 1'b0;
      IsNaN_6U_10U_land_3_lpi_1_dfm_6 <= 1'b0;
      IsNaN_6U_10U_1_land_3_lpi_1_dfm_6 <= 1'b0;
      inp_lookup_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_4 <=
          1'b0;
    end
    else if ( IsNaN_6U_10U_2_aelse_and_2_cse ) begin
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_21 <= IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_20;
      FpMul_6U_10U_lor_8_lpi_1_dfm_st_2 <= or_5022_cse;
      IsNaN_6U_10U_land_3_lpi_1_dfm_6 <= IsNaN_6U_10U_land_3_lpi_1_dfm_5;
      IsNaN_6U_10U_1_land_3_lpi_1_dfm_6 <= IsNaN_6U_10U_1_land_3_lpi_1_dfm_5;
      inp_lookup_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_4 <=
          ~(chn_inp_in_crt_sva_8_315_1 ^ FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_4_1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_p_mant_p1_3_sva_2 <= 22'b0;
    end
    else if ( core_wen & (((~ inp_lookup_3_FpMul_6U_10U_oelse_1_acc_itm_7_1) & (~
        reg_FpMul_6U_10U_lor_5_lpi_1_dfm_3_cse) & or_11_cse & inp_lookup_3_FpMul_6U_10U_else_2_if_acc_itm_6_1)
        | and_1368_rgt) & (~ mux_673_itm) ) begin
      FpMul_6U_10U_p_mant_p1_3_sva_2 <= MUX_v_22_2_2(inp_lookup_3_FpMul_6U_10U_p_mant_p1_mul_tmp,
          FpMul_6U_10U_p_mant_p1_3_sva, and_1368_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_st_112 <= 2'b0;
      chn_inp_in_crt_sva_9_315_1 <= 1'b0;
    end
    else if ( cfg_precision_and_34_cse ) begin
      cfg_precision_1_sva_st_112 <= cfg_precision_1_sva_st_85;
      chn_inp_in_crt_sva_9_315_1 <= chn_inp_in_crt_sva_8_315_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_else_2_else_ac_int_cctor_sva_2 <= 6'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_676_nl) ) begin
      FpMul_6U_10U_else_2_else_ac_int_cctor_sva_2 <= nl_FpMul_6U_10U_else_2_else_ac_int_cctor_sva_2[5:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpMul_6U_10U_else_2_else_slc_FpMul_6U_10U_p_mant_p1_21_itm_2 <=
          1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_678_nl) ) begin
      inp_lookup_4_FpMul_6U_10U_else_2_else_slc_FpMul_6U_10U_p_mant_p1_21_itm_2 <=
          inp_lookup_4_FpMul_6U_10U_p_mant_p1_mul_tmp[21];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_20 <= 1'b0;
      FpMul_6U_10U_lor_1_lpi_1_dfm_st_2 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_23 <= 10'b0;
      IsNaN_6U_10U_land_lpi_1_dfm_6 <= 1'b0;
      IsNaN_6U_10U_1_land_lpi_1_dfm_6 <= 1'b0;
      inp_lookup_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_4 <=
          1'b0;
    end
    else if ( IsNaN_6U_10U_2_aelse_and_3_cse ) begin
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_20 <= IsNaN_6U_10U_2_land_lpi_1_dfm_st_19;
      FpMul_6U_10U_lor_1_lpi_1_dfm_st_2 <= or_5023_cse;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_23 <= FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_3_itm_2;
      IsNaN_6U_10U_land_lpi_1_dfm_6 <= IsNaN_6U_10U_land_lpi_1_dfm_5;
      IsNaN_6U_10U_1_land_lpi_1_dfm_6 <= IsNaN_6U_10U_1_land_lpi_1_dfm_5;
      inp_lookup_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_4 <=
          ~(chn_inp_in_crt_sva_8_331_1 ^ FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_4_1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_p_mant_p1_sva_2 <= 22'b0;
    end
    else if ( core_wen & (((~ inp_lookup_4_FpMul_6U_10U_oelse_1_acc_itm_7_1) & (~
        reg_FpMul_6U_10U_lor_lpi_1_dfm_3_cse) & or_11_cse & inp_lookup_4_FpMul_6U_10U_else_2_if_acc_itm_6_1)
        | and_1372_rgt) & (~ mux_680_itm) ) begin
      FpMul_6U_10U_p_mant_p1_sva_2 <= MUX_v_22_2_2(inp_lookup_4_FpMul_6U_10U_p_mant_p1_mul_tmp,
          FpMul_6U_10U_p_mant_p1_sva, and_1372_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_st_124 <= 2'b0;
      chn_inp_in_crt_sva_9_331_1 <= 1'b0;
    end
    else if ( cfg_precision_and_35_cse ) begin
      cfg_precision_1_sva_st_124 <= cfg_precision_1_sva_st_85;
      chn_inp_in_crt_sva_9_331_1 <= chn_inp_in_crt_sva_8_331_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_10 <= 1'b0;
    end
    else if ( core_wen & ((or_11_cse & main_stage_v_9) | main_stage_v_10_mx0c1) )
        begin
      main_stage_v_10 <= ~ main_stage_v_10_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpAdd_6U_10U_is_a_greater_oif_equal_svs <= 1'b0;
    end
    else if ( core_wen & (~(nand_653_cse | (cfg_precision_1_sva_st_87[0]) | reg_inp_lookup_1_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse
        | and_dcpl_78 | (~ (chn_inp_in_crt_sva_10_739_736_1[0])))) ) begin
      inp_lookup_1_FpAdd_6U_10U_is_a_greater_oif_equal_svs <= inp_lookup_1_FpAdd_6U_10U_is_a_greater_oif_equal_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_24 <= 10'b0;
      FpMul_6U_10U_o_mant_1_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_5_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_24 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_23;
      FpMul_6U_10U_o_mant_1_lpi_1_dfm_7 <= FpMul_6U_10U_o_mant_1_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_27 <= 4'b0;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_15_tmp <= 1'b0;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_15_tmp_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_27 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_26;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_15_tmp <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_14_1_1;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_15_tmp_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_14_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_3_0_1 <= 4'b0;
      reg_FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_5_4_tmp <= 1'b0;
      reg_FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_5_4_tmp_1 <= 1'b0;
    end
    else if ( FpMul_6U_10U_o_expo_and_8_cse ) begin
      FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_3_0_1 <= FpMul_6U_10U_o_expo_1_lpi_1_dfm_3_3_0_mx0w0;
      reg_FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_5_4_tmp <= FpMul_6U_10U_o_expo_1_lpi_1_dfm_3_5_mx0w0;
      reg_FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_5_4_tmp_1 <= FpMul_6U_10U_o_expo_1_lpi_1_dfm_3_4_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_inp_lookup_1_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse <= 1'b0;
      inp_lookup_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_5 <=
          1'b0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_22 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_is_a_greater_and_cse ) begin
      reg_inp_lookup_1_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse <= FpAdd_6U_10U_is_a_greater_acc_itm_6_1;
      inp_lookup_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_5 <=
          inp_lookup_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_4;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_22 <= IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_21;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_st_87 <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_700_nl) ) begin
      cfg_precision_1_sva_st_87 <= cfg_precision_1_sva_st_86;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpAdd_6U_10U_is_a_greater_oif_equal_svs <= 1'b0;
    end
    else if ( core_wen & (~(nand_652_cse | (cfg_precision_1_sva_st_101[0]) | (~ (chn_inp_in_crt_sva_10_739_736_1[1]))
        | and_dcpl_78 | reg_inp_lookup_2_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse))
        ) begin
      inp_lookup_2_FpAdd_6U_10U_is_a_greater_oif_equal_svs <= inp_lookup_2_FpAdd_6U_10U_is_a_greater_oif_equal_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_24 <= 10'b0;
      FpMul_6U_10U_o_mant_2_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_6_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_24 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_23;
      FpMul_6U_10U_o_mant_2_lpi_1_dfm_7 <= FpMul_6U_10U_o_mant_2_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_27 <= 4'b0;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_15_tmp <= 1'b0;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_15_tmp_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_13_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_27 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_26;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_15_tmp <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_14_1_1;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_15_tmp_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_14_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_3_0_1 <= 4'b0;
      reg_FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_5_4_tmp <= 1'b0;
      reg_FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_5_4_tmp_1 <= 1'b0;
    end
    else if ( FpMul_6U_10U_o_expo_and_10_cse ) begin
      FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_3_0_1 <= FpMul_6U_10U_o_expo_2_lpi_1_dfm_3_3_0_mx0w0;
      reg_FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_5_4_tmp <= FpMul_6U_10U_o_expo_2_lpi_1_dfm_3_5_mx0w0;
      reg_FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_5_4_tmp_1 <= FpMul_6U_10U_o_expo_2_lpi_1_dfm_3_4_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_inp_lookup_2_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse <= 1'b0;
      inp_lookup_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_5 <=
          1'b0;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_22 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_is_a_greater_and_2_cse ) begin
      reg_inp_lookup_2_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse <= FpAdd_6U_10U_is_a_greater_acc_1_itm_6_1;
      inp_lookup_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_5 <=
          inp_lookup_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_4;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_22 <= IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_21;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_st_101 <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_718_nl) ) begin
      cfg_precision_1_sva_st_101 <= cfg_precision_1_sva_st_100;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpAdd_6U_10U_is_a_greater_oif_equal_svs <= 1'b0;
    end
    else if ( core_wen & (~((~ main_stage_v_10) | (cfg_precision_1_sva_st_113!=2'b10)
        | (~ (chn_inp_in_crt_sva_10_739_736_1[2])) | and_dcpl_78 | reg_inp_lookup_3_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse))
        ) begin
      inp_lookup_3_FpAdd_6U_10U_is_a_greater_oif_equal_svs <= inp_lookup_3_FpAdd_6U_10U_is_a_greater_oif_equal_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_27 <= 10'b0;
      FpMul_6U_10U_o_mant_3_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_7_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_27 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_26;
      FpMul_6U_10U_o_mant_3_lpi_1_dfm_7 <= FpMul_6U_10U_o_mant_3_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_27 <= 4'b0;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_15_tmp <= 1'b0;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_15_tmp_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_15_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_27 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_26;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_15_tmp <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_14_1_1;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_15_tmp_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_14_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_3_0_1 <= 4'b0;
      reg_inp_lookup_3_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse <= 1'b0;
      inp_lookup_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_5 <=
          1'b0;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_22 <= 1'b0;
      reg_FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_5_4_tmp <= 1'b0;
      reg_FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_5_4_tmp_1 <= 1'b0;
    end
    else if ( FpMul_6U_10U_o_expo_and_12_cse ) begin
      FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_3_0_1 <= FpMul_6U_10U_o_expo_3_lpi_1_dfm_3_3_0_mx0w0;
      reg_inp_lookup_3_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse <= FpAdd_6U_10U_is_a_greater_acc_2_itm_6_1;
      inp_lookup_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_5 <=
          inp_lookup_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_4;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_22 <= IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_21;
      reg_FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_5_4_tmp <= FpMul_6U_10U_o_expo_3_lpi_1_dfm_3_5_mx0w0;
      reg_FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_5_4_tmp_1 <= FpMul_6U_10U_o_expo_3_lpi_1_dfm_3_4_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_st_113 <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_736_nl) ) begin
      cfg_precision_1_sva_st_113 <= cfg_precision_1_sva_st_112;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpAdd_6U_10U_is_a_greater_oif_equal_svs <= 1'b0;
    end
    else if ( core_wen & (~((~ main_stage_v_10) | reg_inp_lookup_4_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse
        | or_dcpl_257 | and_dcpl_78 | (~ (chn_inp_in_crt_sva_10_739_736_1[3]))))
        ) begin
      inp_lookup_4_FpAdd_6U_10U_is_a_greater_oif_equal_svs <= inp_lookup_4_FpAdd_6U_10U_is_a_greater_oif_equal_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_24 <= 10'b0;
      FpMul_6U_10U_o_mant_lpi_1_dfm_7 <= 10'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_8_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_24 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_23;
      FpMul_6U_10U_o_mant_lpi_1_dfm_7 <= FpMul_6U_10U_o_mant_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_27 <= 4'b0;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_15_tmp <= 1'b0;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_15_tmp_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_17_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_27 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_26;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_15_tmp <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_14_1_1;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_15_tmp_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_14_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_o_expo_lpi_1_dfm_6_3_0_1 <= 4'b0;
      reg_inp_lookup_4_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse <= 1'b0;
      inp_lookup_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_5 <=
          1'b0;
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_21 <= 1'b0;
      reg_FpMul_6U_10U_o_expo_lpi_1_dfm_6_5_4_tmp <= 1'b0;
      reg_FpMul_6U_10U_o_expo_lpi_1_dfm_6_5_4_tmp_1 <= 1'b0;
    end
    else if ( FpMul_6U_10U_o_expo_and_14_cse ) begin
      FpMul_6U_10U_o_expo_lpi_1_dfm_6_3_0_1 <= FpMul_6U_10U_o_expo_lpi_1_dfm_3_3_0_mx0w0;
      reg_inp_lookup_4_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse <= FpAdd_6U_10U_is_a_greater_acc_3_itm_6_1;
      inp_lookup_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_5 <=
          inp_lookup_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_4;
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_21 <= IsNaN_6U_10U_2_land_lpi_1_dfm_st_20;
      reg_FpMul_6U_10U_o_expo_lpi_1_dfm_6_5_4_tmp <= FpMul_6U_10U_o_expo_lpi_1_dfm_3_5_mx0w0;
      reg_FpMul_6U_10U_o_expo_lpi_1_dfm_6_5_4_tmp_1 <= FpMul_6U_10U_o_expo_lpi_1_dfm_3_4_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_st_125 <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_754_nl) ) begin
      cfg_precision_1_sva_st_125 <= cfg_precision_1_sva_st_124;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_11 <= 1'b0;
    end
    else if ( core_wen & ((or_11_cse & main_stage_v_10) | main_stage_v_11_mx0c1)
        ) begin
      main_stage_v_11 <= ~ main_stage_v_11_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_inp_lookup_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse
          <= 1'b0;
      FpAdd_6U_10U_a_int_mant_p1_1_sva_2 <= 23'b0;
      FpAdd_6U_10U_b_int_mant_p1_1_sva_2 <= 23'b0;
      FpAdd_6U_10U_is_a_greater_lor_1_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_25 <= 1'b0;
      IsNaN_6U_10U_3_land_1_lpi_1_dfm_7 <= 1'b0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_23 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_is_addition_and_cse ) begin
      reg_inp_lookup_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse
          <= inp_lookup_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_5;
      FpAdd_6U_10U_a_int_mant_p1_1_sva_2 <= inp_lookup_1_FpAdd_6U_10U_a_int_mant_p1_lshift_itm;
      FpAdd_6U_10U_b_int_mant_p1_1_sva_2 <= inp_lookup_1_FpAdd_6U_10U_b_int_mant_p1_lshift_itm;
      FpAdd_6U_10U_is_a_greater_lor_1_lpi_1_dfm_5 <= FpAdd_6U_10U_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_25 <= IsNaN_6U_10U_2_land_1_lpi_1_dfm_24;
      IsNaN_6U_10U_3_land_1_lpi_1_dfm_7 <= IsNaN_6U_10U_3_land_1_lpi_1_dfm_6;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_23 <= IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_22;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_st_88 <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_760_nl) ) begin
      cfg_precision_1_sva_st_88 <= cfg_precision_1_sva_st_87;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_inp_lookup_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse
          <= 1'b0;
      FpAdd_6U_10U_a_int_mant_p1_2_sva_2 <= 23'b0;
      FpAdd_6U_10U_b_int_mant_p1_2_sva_2 <= 23'b0;
      FpAdd_6U_10U_is_a_greater_lor_2_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_25 <= 1'b0;
      IsNaN_6U_10U_3_land_2_lpi_1_dfm_7 <= 1'b0;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_23 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_is_addition_and_2_cse ) begin
      reg_inp_lookup_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse
          <= inp_lookup_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_5;
      FpAdd_6U_10U_a_int_mant_p1_2_sva_2 <= inp_lookup_2_FpAdd_6U_10U_a_int_mant_p1_lshift_itm;
      FpAdd_6U_10U_b_int_mant_p1_2_sva_2 <= inp_lookup_2_FpAdd_6U_10U_b_int_mant_p1_lshift_itm;
      FpAdd_6U_10U_is_a_greater_lor_2_lpi_1_dfm_5 <= FpAdd_6U_10U_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_25 <= IsNaN_6U_10U_2_land_2_lpi_1_dfm_24;
      IsNaN_6U_10U_3_land_2_lpi_1_dfm_7 <= IsNaN_6U_10U_3_land_2_lpi_1_dfm_6;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_23 <= IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_22;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_st_102 <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_765_nl) ) begin
      cfg_precision_1_sva_st_102 <= cfg_precision_1_sva_st_101;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_inp_lookup_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse
          <= 1'b0;
      FpAdd_6U_10U_a_int_mant_p1_3_sva_2 <= 23'b0;
      FpAdd_6U_10U_b_int_mant_p1_3_sva_2 <= 23'b0;
      FpAdd_6U_10U_is_a_greater_lor_3_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_25 <= 1'b0;
      IsNaN_6U_10U_3_land_3_lpi_1_dfm_7 <= 1'b0;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_23 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_is_addition_and_4_cse ) begin
      reg_inp_lookup_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse
          <= inp_lookup_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_5;
      FpAdd_6U_10U_a_int_mant_p1_3_sva_2 <= inp_lookup_3_FpAdd_6U_10U_a_int_mant_p1_lshift_itm;
      FpAdd_6U_10U_b_int_mant_p1_3_sva_2 <= inp_lookup_3_FpAdd_6U_10U_b_int_mant_p1_lshift_itm;
      FpAdd_6U_10U_is_a_greater_lor_3_lpi_1_dfm_5 <= FpAdd_6U_10U_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_25 <= IsNaN_6U_10U_2_land_3_lpi_1_dfm_24;
      IsNaN_6U_10U_3_land_3_lpi_1_dfm_7 <= IsNaN_6U_10U_3_land_3_lpi_1_dfm_6;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_23 <= IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_22;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_st_114 <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_770_nl) ) begin
      cfg_precision_1_sva_st_114 <= cfg_precision_1_sva_st_113;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_inp_lookup_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse
          <= 1'b0;
      FpAdd_6U_10U_a_int_mant_p1_sva_2 <= 23'b0;
      FpAdd_6U_10U_b_int_mant_p1_sva_2 <= 23'b0;
      FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_2_land_lpi_1_dfm_25 <= 1'b0;
      IsNaN_6U_10U_3_land_lpi_1_dfm_7 <= 1'b0;
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_22 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_is_addition_and_6_cse ) begin
      reg_inp_lookup_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse
          <= inp_lookup_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_5;
      FpAdd_6U_10U_a_int_mant_p1_sva_2 <= inp_lookup_4_FpAdd_6U_10U_a_int_mant_p1_lshift_itm;
      FpAdd_6U_10U_b_int_mant_p1_sva_2 <= inp_lookup_4_FpAdd_6U_10U_b_int_mant_p1_lshift_itm;
      FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_5 <= FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_1_mx0w0;
      IsNaN_6U_10U_2_land_lpi_1_dfm_25 <= IsNaN_6U_10U_2_land_lpi_1_dfm_24;
      IsNaN_6U_10U_3_land_lpi_1_dfm_7 <= IsNaN_6U_10U_3_land_lpi_1_dfm_6;
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_22 <= IsNaN_6U_10U_2_land_lpi_1_dfm_st_21;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_st_126 <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_775_nl) ) begin
      cfg_precision_1_sva_st_126 <= cfg_precision_1_sva_st_125;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_12 <= 1'b0;
    end
    else if ( core_wen & ((or_11_cse & main_stage_v_11) | main_stage_v_12_mx0c1)
        ) begin
      main_stage_v_12 <= ~ main_stage_v_12_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsInf_6U_23U_land_1_lpi_1_dfm <= 1'b0;
      IsNaN_6U_23U_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( IsInf_6U_23U_aelse_and_cse ) begin
      IsInf_6U_23U_land_1_lpi_1_dfm <= IsInf_6U_23U_land_1_lpi_1_dfm_mx0w0;
      IsNaN_6U_23U_land_1_lpi_1_dfm <= IsNaN_6U_23U_IsNaN_6U_23U_nor_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_qr_2_lpi_1_dfm_4_3_0_1 <= 4'b0;
      reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_4_5_4_tmp <= 1'b0;
      reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_4_5_4_tmp_1 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_and_43_cse ) begin
      FpAdd_6U_10U_qr_2_lpi_1_dfm_4_3_0_1 <= FpAdd_6U_10U_qr_2_lpi_1_dfm_3_3_0_1;
      reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_4_5_4_tmp <= reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_3_5_4_tmp;
      reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_4_5_4_tmp_1 <= reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_3_5_4_tmp_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_1_sva_st_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_781_nl) ) begin
      FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_1_sva_st_2 <= inp_lookup_1_FpAdd_6U_10U_if_3_if_acc_1_itm_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_4 <= 24'b0;
    end
    else if ( core_wen & ((or_11_cse & reg_inp_lookup_1_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse)
        | and_1386_rgt) & (~ mux_782_itm) ) begin
      FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_4 <= MUX_v_24_2_2(FpAdd_6U_10U_int_mant_p1_1_sva,
          FpAdd_6U_10U_asn_23_mx0w1, and_1386_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_23U_leading_sign_23_0_rtn_1_sva_2 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_784_nl)) ) begin
      IntLeadZero_23U_leading_sign_23_0_rtn_1_sva_2 <= libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_12;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpNormalize_6U_23U_lor_1_lpi_1_dfm_4_cse <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_785_nl) ) begin
      reg_FpNormalize_6U_23U_lor_1_lpi_1_dfm_4_cse <= FpNormalize_6U_23U_if_FpNormalize_6U_23U_if_nand_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_3_land_1_lpi_1_dfm_8 <= 1'b0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_26 <= 1'b0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_24 <= 1'b0;
      FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_1_sva_2 <= 1'b0;
      inp_lookup_1_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_3_aelse_and_cse ) begin
      IsNaN_6U_10U_3_land_1_lpi_1_dfm_8 <= IsNaN_6U_10U_3_land_1_lpi_1_dfm_7;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_26 <= IsNaN_6U_10U_2_land_1_lpi_1_dfm_25;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_24 <= IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_23;
      FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_1_sva_2 <= inp_lookup_1_FpAdd_6U_10U_if_3_if_acc_1_itm_5;
      inp_lookup_1_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2 <= FpAdd_6U_10U_int_mant_p1_1_lpi_1_dfm_mx0[23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_26 <= 10'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_788_nl)) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_26 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_25;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_29 <= 4'b0;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_17_tmp <= 1'b0;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_17_tmp_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_19_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_29 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_28;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_17_tmp <= reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_16_tmp;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_17_tmp_1 <= reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_16_tmp_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_st_89 <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_791_nl) ) begin
      cfg_precision_1_sva_st_89 <= cfg_precision_1_sva_st_88;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsInf_6U_23U_land_2_lpi_1_dfm <= 1'b0;
      IsNaN_6U_23U_land_2_lpi_1_dfm <= 1'b0;
    end
    else if ( IsInf_6U_23U_aelse_and_1_cse ) begin
      IsInf_6U_23U_land_2_lpi_1_dfm <= IsInf_6U_23U_land_2_lpi_1_dfm_mx0w0;
      IsNaN_6U_23U_land_2_lpi_1_dfm <= IsNaN_6U_23U_IsNaN_6U_23U_nor_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_qr_3_lpi_1_dfm_4_3_0_1 <= 4'b0;
      reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_4_5_4_tmp <= 1'b0;
      reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_4_5_4_tmp_1 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_and_45_cse ) begin
      FpAdd_6U_10U_qr_3_lpi_1_dfm_4_3_0_1 <= FpAdd_6U_10U_qr_3_lpi_1_dfm_3_3_0_1;
      reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_4_5_4_tmp <= reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_3_5_4_tmp;
      reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_4_5_4_tmp_1 <= reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_3_5_4_tmp_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_2_sva_st_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_798_nl)) ) begin
      FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_2_sva_st_2 <= inp_lookup_2_FpAdd_6U_10U_if_3_if_acc_1_itm_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_4 <= 24'b0;
    end
    else if ( core_wen & ((or_11_cse & reg_inp_lookup_2_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse)
        | and_1388_rgt) & (~ mux_799_itm) ) begin
      FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_4 <= MUX_v_24_2_2(FpAdd_6U_10U_int_mant_p1_2_sva,
          FpAdd_6U_10U_asn_20_mx0w1, and_1388_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_23U_leading_sign_23_0_rtn_2_sva_2 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_800_nl)) ) begin
      IntLeadZero_23U_leading_sign_23_0_rtn_2_sva_2 <= libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_13;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpNormalize_6U_23U_lor_2_lpi_1_dfm_4_cse <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_801_nl) ) begin
      reg_FpNormalize_6U_23U_lor_2_lpi_1_dfm_4_cse <= FpNormalize_6U_23U_if_FpNormalize_6U_23U_if_nand_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_3_land_2_lpi_1_dfm_8 <= 1'b0;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_26 <= 1'b0;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_24 <= 1'b0;
      FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_2_sva_2 <= 1'b0;
      inp_lookup_2_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_3_aelse_and_1_cse ) begin
      IsNaN_6U_10U_3_land_2_lpi_1_dfm_8 <= IsNaN_6U_10U_3_land_2_lpi_1_dfm_7;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_26 <= IsNaN_6U_10U_2_land_2_lpi_1_dfm_25;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_24 <= IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_23;
      FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_2_sva_2 <= inp_lookup_2_FpAdd_6U_10U_if_3_if_acc_1_itm_5;
      inp_lookup_2_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2 <= FpAdd_6U_10U_int_mant_p1_2_lpi_1_dfm_mx0[23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_26 <= 10'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_802_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_26 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_25;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_29 <= 4'b0;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_17_tmp <= 1'b0;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_17_tmp_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_21_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_29 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_28;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_17_tmp <= reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_16_tmp;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_17_tmp_1 <= reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_16_tmp_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_st_103 <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_805_nl) ) begin
      cfg_precision_1_sva_st_103 <= cfg_precision_1_sva_st_102;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsInf_6U_23U_land_3_lpi_1_dfm <= 1'b0;
      IsNaN_6U_23U_land_3_lpi_1_dfm <= 1'b0;
    end
    else if ( IsInf_6U_23U_aelse_and_2_cse ) begin
      IsInf_6U_23U_land_3_lpi_1_dfm <= IsInf_6U_23U_land_3_lpi_1_dfm_mx0w0;
      IsNaN_6U_23U_land_3_lpi_1_dfm <= IsNaN_6U_23U_IsNaN_6U_23U_nor_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_qr_4_lpi_1_dfm_4_3_0_1 <= 4'b0;
      reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_4_5_4_tmp <= 1'b0;
      reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_4_5_4_tmp_1 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_and_47_cse ) begin
      FpAdd_6U_10U_qr_4_lpi_1_dfm_4_3_0_1 <= FpAdd_6U_10U_qr_4_lpi_1_dfm_3_3_0_1;
      reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_4_5_4_tmp <= reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_3_5_4_tmp;
      reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_4_5_4_tmp_1 <= reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_3_5_4_tmp_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_3_sva_st_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_815_nl) ) begin
      FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_3_sva_st_2 <= inp_lookup_3_FpAdd_6U_10U_if_3_if_acc_1_itm_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_4 <= 24'b0;
    end
    else if ( core_wen & ((or_11_cse & reg_inp_lookup_3_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse)
        | and_1390_rgt) & (~ mux_816_itm) ) begin
      FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_4 <= MUX_v_24_2_2(FpAdd_6U_10U_int_mant_p1_3_sva,
          FpAdd_6U_10U_asn_17_mx0w1, and_1390_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_23U_leading_sign_23_0_rtn_3_sva_2 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_818_nl) ) begin
      IntLeadZero_23U_leading_sign_23_0_rtn_3_sva_2 <= libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_14;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpNormalize_6U_23U_lor_3_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_819_nl)) ) begin
      FpNormalize_6U_23U_lor_3_lpi_1_dfm_5 <= FpNormalize_6U_23U_if_FpNormalize_6U_23U_if_nand_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_3_land_3_lpi_1_dfm_8 <= 1'b0;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_26 <= 1'b0;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_24 <= 1'b0;
      FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_3_sva_2 <= 1'b0;
      inp_lookup_3_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_3_aelse_and_2_cse ) begin
      IsNaN_6U_10U_3_land_3_lpi_1_dfm_8 <= IsNaN_6U_10U_3_land_3_lpi_1_dfm_7;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_26 <= IsNaN_6U_10U_2_land_3_lpi_1_dfm_25;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_24 <= IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_23;
      FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_3_sva_2 <= inp_lookup_3_FpAdd_6U_10U_if_3_if_acc_1_itm_5;
      inp_lookup_3_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2 <= FpAdd_6U_10U_int_mant_p1_3_lpi_1_dfm_mx0[23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_29 <= 10'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_820_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_29 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_28;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_29 <= 4'b0;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_17_tmp <= 1'b0;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_17_tmp_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_23_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_29 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_28;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_17_tmp <= reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_16_tmp;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_17_tmp_1 <= reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_16_tmp_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_st_115 <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_823_nl) ) begin
      cfg_precision_1_sva_st_115 <= cfg_precision_1_sva_st_114;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsInf_6U_23U_land_lpi_1_dfm <= 1'b0;
      IsNaN_6U_23U_land_lpi_1_dfm <= 1'b0;
    end
    else if ( IsInf_6U_23U_aelse_and_3_cse ) begin
      IsInf_6U_23U_land_lpi_1_dfm <= IsInf_6U_23U_land_lpi_1_dfm_mx0w0;
      IsNaN_6U_23U_land_lpi_1_dfm <= IsNaN_6U_23U_IsNaN_6U_23U_nor_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_qr_lpi_1_dfm_4_3_0_1 <= 4'b0;
      reg_FpAdd_6U_10U_qr_lpi_1_dfm_4_5_4_tmp <= 1'b0;
      reg_FpAdd_6U_10U_qr_lpi_1_dfm_4_5_4_tmp_1 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_and_49_cse ) begin
      FpAdd_6U_10U_qr_lpi_1_dfm_4_3_0_1 <= FpAdd_6U_10U_qr_lpi_1_dfm_3_3_0_1;
      reg_FpAdd_6U_10U_qr_lpi_1_dfm_4_5_4_tmp <= reg_FpAdd_6U_10U_qr_lpi_1_dfm_3_5_4_tmp;
      reg_FpAdd_6U_10U_qr_lpi_1_dfm_4_5_4_tmp_1 <= reg_FpAdd_6U_10U_qr_lpi_1_dfm_3_5_4_tmp_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_sva_st_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_828_nl) ) begin
      FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_sva_st_2 <= inp_lookup_4_FpAdd_6U_10U_if_3_if_acc_1_itm_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_4 <= 24'b0;
    end
    else if ( core_wen & ((or_11_cse & reg_inp_lookup_4_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_3_cse)
        | and_1392_rgt) & (~ mux_829_itm) ) begin
      FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_4 <= MUX_v_24_2_2(FpAdd_6U_10U_int_mant_p1_sva,
          FpAdd_6U_10U_asn_mx0w1, and_1392_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_23U_leading_sign_23_0_rtn_sva_2 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_830_nl)) ) begin
      IntLeadZero_23U_leading_sign_23_0_rtn_sva_2 <= libraries_leading_sign_23_0_aebf38bbf639c970da88b55f070b6a2d5444_15;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpNormalize_6U_23U_lor_lpi_1_dfm_4_cse <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_831_nl) ) begin
      reg_FpNormalize_6U_23U_lor_lpi_1_dfm_4_cse <= FpNormalize_6U_23U_if_FpNormalize_6U_23U_if_nand_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_3_land_lpi_1_dfm_8 <= 1'b0;
      IsNaN_6U_10U_2_land_lpi_1_dfm_26 <= 1'b0;
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_23 <= 1'b0;
      FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_sva_2 <= 1'b0;
      inp_lookup_4_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_3_aelse_and_3_cse ) begin
      IsNaN_6U_10U_3_land_lpi_1_dfm_8 <= IsNaN_6U_10U_3_land_lpi_1_dfm_7;
      IsNaN_6U_10U_2_land_lpi_1_dfm_26 <= IsNaN_6U_10U_2_land_lpi_1_dfm_25;
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_23 <= IsNaN_6U_10U_2_land_lpi_1_dfm_st_22;
      FpAdd_6U_10U_if_3_if_slc_FpAdd_6U_10U_if_3_if_acc_1_5_mdf_sva_2 <= inp_lookup_4_FpAdd_6U_10U_if_3_if_acc_1_itm_5;
      inp_lookup_4_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2 <= FpAdd_6U_10U_int_mant_p1_lpi_1_dfm_mx0[23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_26 <= 10'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_833_nl)) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_26 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_25;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_29 <= 4'b0;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_17_tmp <= 1'b0;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_17_tmp_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_25_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_29 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_28;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_17_tmp <= reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_16_tmp;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_17_tmp_1 <= reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_16_tmp_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_st_127 <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_835_nl) ) begin
      cfg_precision_1_sva_st_127 <= cfg_precision_1_sva_st_126;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_mux_1057_itm_4 <= 1'b0;
      inp_lookup_if_unequal_tmp_19 <= 1'b0;
      chn_inp_in_crt_sva_12_739_736_1 <= 4'b0;
      IsNaN_6U_23U_3_land_lpi_1_dfm_10 <= 1'b0;
      IsNaN_6U_23U_3_land_1_lpi_1_dfm_10 <= 1'b0;
      inp_lookup_else_unequal_tmp_38 <= 1'b0;
      inp_lookup_mux_259_itm_4 <= 1'b0;
      inp_lookup_mux_791_itm_4 <= 1'b0;
      IsNaN_6U_23U_3_land_3_lpi_1_dfm_10 <= 1'b0;
      IsNaN_6U_23U_3_land_2_lpi_1_dfm_10 <= 1'b0;
      inp_lookup_mux_525_itm_4 <= 1'b0;
    end
    else if ( inp_lookup_and_cse ) begin
      inp_lookup_mux_1057_itm_4 <= inp_lookup_mux_1057_itm_3;
      inp_lookup_if_unequal_tmp_19 <= inp_lookup_if_unequal_tmp_12;
      chn_inp_in_crt_sva_12_739_736_1 <= chn_inp_in_crt_sva_11_739_736_1;
      IsNaN_6U_23U_3_land_lpi_1_dfm_10 <= IsNaN_6U_23U_3_land_lpi_1_dfm_9;
      IsNaN_6U_23U_3_land_1_lpi_1_dfm_10 <= IsNaN_6U_23U_3_land_1_lpi_1_dfm_9;
      inp_lookup_else_unequal_tmp_38 <= inp_lookup_else_unequal_tmp_37;
      inp_lookup_mux_259_itm_4 <= inp_lookup_mux_259_itm_3;
      inp_lookup_mux_791_itm_4 <= inp_lookup_mux_791_itm_3;
      IsNaN_6U_23U_3_land_3_lpi_1_dfm_10 <= IsNaN_6U_23U_3_land_3_lpi_1_dfm_9;
      IsNaN_6U_23U_3_land_2_lpi_1_dfm_10 <= IsNaN_6U_23U_3_land_2_lpi_1_dfm_9;
      inp_lookup_mux_525_itm_4 <= inp_lookup_mux_525_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_122_itm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_837_nl)) ) begin
      inp_lookup_else_mux_122_itm_8 <= inp_lookup_else_mux_122_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_1_lpi_1_dfm_12_30_0_1 <= 31'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_839_nl) ) begin
      IntSaturation_51U_32U_o_1_lpi_1_dfm_12_30_0_1 <= IntSaturation_51U_32U_o_1_lpi_1_dfm_11_30_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_lpi_1_dfm_12 <= 3'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_8_4_1 <= 1'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_8_3_0_1 <= 4'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_lpi_1_dfm_12 <= 10'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_19_itm_8
          <= 1'b0;
    end
    else if ( FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_and_cse ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_lpi_1_dfm_12 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_lpi_1_dfm_11;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_8_4_1 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_7_4_1;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_8_3_0_1 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_7_3_0_1;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_lpi_1_dfm_12 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_lpi_1_dfm_11;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_19_itm_8
          <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_19_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_10_17_1_itm <= 8'b0;
    end
    else if ( or_11_cse & core_wen & main_stage_v_11 & (~ (chn_inp_in_crt_sva_11_739_736_1[3]))
        & inp_lookup_else_unequal_tmp_37 ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_10_17_1_itm <= reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_9_17_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_10_17_1_1_itm <= 9'b0;
    end
    else if ( and_dcpl_2279 & (~ (chn_inp_in_crt_sva_11_739_736_1[3])) & or_11_cse
        ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_10_17_1_1_itm <= reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_9_17_1_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_lpi_1_dfm_12_30_0_1 <= 31'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_844_nl) ) begin
      IntSaturation_51U_32U_o_lpi_1_dfm_12_30_0_1 <= IntSaturation_51U_32U_o_lpi_1_dfm_11_30_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_10_17_1_itm <= 8'b0;
    end
    else if ( or_11_cse & core_wen & main_stage_v_11 & (~ (chn_inp_in_crt_sva_11_739_736_1[0]))
        & inp_lookup_else_unequal_tmp_37 ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_10_17_1_itm <= reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_9_17_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_10_17_1_1_itm <= 9'b0;
    end
    else if ( and_dcpl_2279 & (~ (chn_inp_in_crt_sva_11_739_736_1[0])) & or_11_cse
        ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_10_17_1_1_itm <= reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_9_17_1_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_4_itm_8
          <= 1'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_1_lpi_1_dfm_12 <= 10'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_8_4_1 <= 1'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_8_3_0_1 <= 4'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_1_lpi_1_dfm_12 <= 3'b0;
    end
    else if ( FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_cse ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_4_itm_8
          <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_4_itm_7;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_1_lpi_1_dfm_12 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_1_lpi_1_dfm_11;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_8_4_1 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_7_4_1;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_8_3_0_1 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_7_3_0_1;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_1_lpi_1_dfm_12 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_1_lpi_1_dfm_11;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_491_itm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_842_nl)) ) begin
      inp_lookup_else_mux_491_itm_8 <= inp_lookup_else_mux_491_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_245_itm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_847_nl)) ) begin
      inp_lookup_else_mux_245_itm_8 <= inp_lookup_else_mux_245_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_2_lpi_1_dfm_12_30_0_1 <= 31'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_848_nl) ) begin
      IntSaturation_51U_32U_o_2_lpi_1_dfm_12_30_0_1 <= IntSaturation_51U_32U_o_2_lpi_1_dfm_11_30_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_3_lpi_1_dfm_12 <= 3'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_8_4_1 <= 1'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_8_3_0_1 <= 4'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_3_lpi_1_dfm_12 <= 10'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_14_itm_8
          <= 1'b0;
    end
    else if ( FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_and_6_cse ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_3_lpi_1_dfm_12 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_3_lpi_1_dfm_11;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_8_4_1 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_7_4_1;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_8_3_0_1 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_7_3_0_1;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_3_lpi_1_dfm_12 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_3_lpi_1_dfm_11;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_14_itm_8
          <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_14_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_10_17_1_itm <= 8'b0;
    end
    else if ( or_11_cse & core_wen & main_stage_v_11 & (~ (chn_inp_in_crt_sva_11_739_736_1[2]))
        & inp_lookup_else_unequal_tmp_37 ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_10_17_1_itm <= reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_9_17_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_10_17_1_1_itm <= 9'b0;
    end
    else if ( and_dcpl_2279 & (~ (chn_inp_in_crt_sva_11_739_736_1[2])) & or_11_cse
        ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_10_17_1_1_itm <= reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_9_17_1_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_3_lpi_1_dfm_12_30_0_1 <= 31'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_852_nl) ) begin
      IntSaturation_51U_32U_o_3_lpi_1_dfm_12_30_0_1 <= IntSaturation_51U_32U_o_3_lpi_1_dfm_11_30_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_10_17_1_itm <= 8'b0;
    end
    else if ( or_11_cse & core_wen & main_stage_v_11 & (~ (chn_inp_in_crt_sva_11_739_736_1[1]))
        & inp_lookup_else_unequal_tmp_37 ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_10_17_1_itm <= reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_9_17_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_10_17_1_1_itm <= 9'b0;
    end
    else if ( and_dcpl_2279 & (~ (chn_inp_in_crt_sva_11_739_736_1[1])) & or_11_cse
        ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_10_17_1_1_itm <= reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_9_17_1_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_9_itm_8
          <= 1'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_2_lpi_1_dfm_12 <= 10'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_8_4_1 <= 1'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_8_3_0_1 <= 4'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_2_lpi_1_dfm_12 <= 3'b0;
    end
    else if ( FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_2_cse ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_9_itm_8
          <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_9_itm_7;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_2_lpi_1_dfm_12 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_2_lpi_1_dfm_11;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_8_4_1 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_7_4_1;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_8_3_0_1 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_7_3_0_1;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_2_lpi_1_dfm_12 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_2_lpi_1_dfm_11;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_368_itm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_850_nl)) ) begin
      inp_lookup_else_mux_368_itm_8 <= inp_lookup_else_mux_368_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_qr_2_lpi_1_dfm_3_3_0_1 <= 4'b0;
      reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_3_5_4_tmp <= 1'b0;
      reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_3_5_4_tmp_1 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_and_51_cse ) begin
      FpAdd_6U_10U_qr_2_lpi_1_dfm_3_3_0_1 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_27,
          FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_3_0_1, FpAdd_6U_10U_qr_2_lpi_1_dfm_3_0,
          {and_dcpl_930 , and_dcpl_935 , and_dcpl_936});
      reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_3_5_4_tmp <= MUX1HOT_s_1_3_2(reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_15_tmp,
          reg_FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_5_4_tmp, reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_5_4_tmp,
          {and_dcpl_930 , and_dcpl_935 , and_dcpl_936});
      reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_3_5_4_tmp_1 <= MUX1HOT_s_1_3_2(reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_15_tmp_1,
          reg_FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_5_4_tmp_1, reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_5_4_tmp_1,
          {and_dcpl_930 , and_dcpl_935 , and_dcpl_936});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_qr_3_lpi_1_dfm_3_3_0_1 <= 4'b0;
      reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_3_5_4_tmp <= 1'b0;
      reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_3_5_4_tmp_1 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_and_53_cse ) begin
      FpAdd_6U_10U_qr_3_lpi_1_dfm_3_3_0_1 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_27,
          FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_3_0_1, FpAdd_6U_10U_qr_3_lpi_1_dfm_3_0,
          {and_dcpl_940 , and_dcpl_944 , and_dcpl_945});
      reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_3_5_4_tmp <= MUX1HOT_s_1_3_2(reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_15_tmp,
          reg_FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_5_4_tmp, reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_5_4_tmp,
          {and_dcpl_940 , and_dcpl_944 , and_dcpl_945});
      reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_3_5_4_tmp_1 <= MUX1HOT_s_1_3_2(reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_15_tmp_1,
          reg_FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_5_4_tmp_1, reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_5_4_tmp_1,
          {and_dcpl_940 , and_dcpl_944 , and_dcpl_945});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_qr_4_lpi_1_dfm_3_3_0_1 <= 4'b0;
      reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_3_5_4_tmp <= 1'b0;
      reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_3_5_4_tmp_1 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_and_55_cse ) begin
      FpAdd_6U_10U_qr_4_lpi_1_dfm_3_3_0_1 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_27,
          FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_3_0_1, FpAdd_6U_10U_qr_4_lpi_1_dfm_3_0,
          {and_dcpl_949 , and_dcpl_954 , and_dcpl_955});
      reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_3_5_4_tmp <= MUX1HOT_s_1_3_2(reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_15_tmp,
          reg_FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_5_4_tmp, reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_5_4_tmp,
          {and_dcpl_949 , and_dcpl_954 , and_dcpl_955});
      reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_3_5_4_tmp_1 <= MUX1HOT_s_1_3_2(reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_15_tmp_1,
          reg_FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_5_4_tmp_1, reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_5_4_tmp_1,
          {and_dcpl_949 , and_dcpl_954 , and_dcpl_955});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_qr_lpi_1_dfm_3_3_0_1 <= 4'b0;
      reg_FpAdd_6U_10U_qr_lpi_1_dfm_3_5_4_tmp <= 1'b0;
      reg_FpAdd_6U_10U_qr_lpi_1_dfm_3_5_4_tmp_1 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_and_57_cse ) begin
      FpAdd_6U_10U_qr_lpi_1_dfm_3_3_0_1 <= MUX1HOT_v_4_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_27,
          FpMul_6U_10U_o_expo_lpi_1_dfm_6_3_0_1, FpAdd_6U_10U_qr_lpi_1_dfm_3_0, {and_dcpl_959
          , and_dcpl_961 , and_dcpl_962});
      reg_FpAdd_6U_10U_qr_lpi_1_dfm_3_5_4_tmp <= MUX1HOT_s_1_3_2(reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_15_tmp,
          reg_FpMul_6U_10U_o_expo_lpi_1_dfm_6_5_4_tmp, reg_FpAdd_6U_10U_qr_lpi_1_dfm_5_4_tmp,
          {and_dcpl_959 , and_dcpl_961 , and_dcpl_962});
      reg_FpAdd_6U_10U_qr_lpi_1_dfm_3_5_4_tmp_1 <= MUX1HOT_s_1_3_2(reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_15_tmp_1,
          reg_FpMul_6U_10U_o_expo_lpi_1_dfm_6_5_4_tmp_1, reg_FpAdd_6U_10U_qr_lpi_1_dfm_5_4_tmp_1,
          {and_dcpl_959 , and_dcpl_961 , and_dcpl_962});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_14_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_14_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_26 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_14_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_14_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_26 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_26 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_14_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_14_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_26 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_14_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_14_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_26 <= 4'b0;
      FpMul_6U_10U_o_sign_lpi_1_dfm_5 <= 1'b0;
      FpMul_6U_10U_o_sign_3_lpi_1_dfm_5 <= 1'b0;
      FpMul_6U_10U_o_sign_2_lpi_1_dfm_5 <= 1'b0;
      FpMul_6U_10U_o_sign_1_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_23U_3_land_lpi_1_dfm_7 <= 1'b0;
      IsNaN_6U_23U_3_land_3_lpi_1_dfm_7 <= 1'b0;
      IsNaN_6U_23U_3_land_2_lpi_1_dfm_7 <= 1'b0;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_23 <= 1'b0;
      IsNaN_6U_23U_3_land_1_lpi_1_dfm_7 <= 1'b0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_23 <= 1'b0;
      inp_lookup_else_unequal_tmp_35 <= 1'b0;
      chn_inp_in_crt_sva_9_739_736_1 <= 4'b0;
    end
    else if ( chn_inp_in_flow_and_32_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_14_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_13_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_14_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_13_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_26 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_25;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_14_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_13_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_14_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_13_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_26 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_25;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_26 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_25;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_14_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_13_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_14_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_13_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_26 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_25;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_14_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_13_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_14_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_13_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_26 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_25;
      FpMul_6U_10U_o_sign_lpi_1_dfm_5 <= FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_4_1;
      FpMul_6U_10U_o_sign_3_lpi_1_dfm_5 <= FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_4_1;
      FpMul_6U_10U_o_sign_2_lpi_1_dfm_5 <= FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_4_1;
      FpMul_6U_10U_o_sign_1_lpi_1_dfm_5 <= FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_4_1;
      IsNaN_6U_23U_3_land_lpi_1_dfm_7 <= and_3588_cse;
      IsNaN_6U_23U_3_land_3_lpi_1_dfm_7 <= and_3587_cse;
      IsNaN_6U_23U_3_land_2_lpi_1_dfm_7 <= and_3586_cse;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_23 <= IsNaN_6U_10U_2_land_2_lpi_1_dfm_22;
      IsNaN_6U_23U_3_land_1_lpi_1_dfm_7 <= and_3585_cse;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_23 <= IsNaN_6U_10U_2_land_1_lpi_1_dfm_22;
      inp_lookup_else_unequal_tmp_35 <= inp_lookup_else_unequal_tmp_55;
      chn_inp_in_crt_sva_9_739_736_1 <= chn_inp_in_crt_sva_8_739_736_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_p_mant_p1_1_sva <= 22'b0;
    end
    else if ( core_wen & (~(or_dcpl_295 | inp_lookup_1_FpMul_6U_10U_oelse_1_acc_itm_7_1
        | (~ (chn_inp_in_crt_sva_8_739_736_1[0])) | reg_FpMul_6U_10U_lor_3_lpi_1_dfm_3_cse
        | (~ inp_lookup_1_FpMul_6U_10U_else_2_if_acc_itm_6_1) | and_dcpl_78)) ) begin
      FpMul_6U_10U_p_mant_p1_1_sva <= inp_lookup_1_FpMul_6U_10U_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_p_mant_p1_2_sva <= 22'b0;
    end
    else if ( core_wen & (~(nand_544_cse | (~ (chn_inp_in_crt_sva_8_739_736_1[1]))
        | inp_lookup_2_FpMul_6U_10U_oelse_1_acc_itm_7_1 | (cfg_precision_1_sva_st_85[0])
        | reg_FpMul_6U_10U_lor_4_lpi_1_dfm_3_cse | (~ inp_lookup_2_FpMul_6U_10U_else_2_if_acc_itm_6_1)
        | and_dcpl_78)) ) begin
      FpMul_6U_10U_p_mant_p1_2_sva <= inp_lookup_2_FpMul_6U_10U_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_p_mant_p1_3_sva <= 22'b0;
    end
    else if ( core_wen & (~(or_dcpl_295 | inp_lookup_3_FpMul_6U_10U_oelse_1_acc_itm_7_1
        | (~ (chn_inp_in_crt_sva_8_739_736_1[2])) | reg_FpMul_6U_10U_lor_5_lpi_1_dfm_3_cse
        | (~ inp_lookup_3_FpMul_6U_10U_else_2_if_acc_itm_6_1) | and_dcpl_78)) ) begin
      FpMul_6U_10U_p_mant_p1_3_sva <= inp_lookup_3_FpMul_6U_10U_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_p_mant_p1_sva <= 22'b0;
    end
    else if ( core_wen & (~(or_dcpl_295 | inp_lookup_4_FpMul_6U_10U_oelse_1_acc_itm_7_1
        | (~ (chn_inp_in_crt_sva_8_739_736_1[3])) | reg_FpMul_6U_10U_lor_lpi_1_dfm_3_cse
        | (~ inp_lookup_4_FpMul_6U_10U_else_2_if_acc_itm_6_1) | and_dcpl_78)) ) begin
      FpMul_6U_10U_p_mant_p1_sva <= inp_lookup_4_FpMul_6U_10U_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_itm <= 10'b0;
    end
    else if ( core_wen & (~(IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_19 | (~ main_stage_v_7)
        | (cfg_precision_1_sva_st_84!=2'b10) | and_dcpl_78 | (chn_inp_in_crt_sva_7_739_736_1[0])))
        ) begin
      FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_itm <= FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_8_land_1_lpi_1_dfm_7 <= 1'b0;
      IsNaN_6U_10U_9_land_1_lpi_1_dfm_8 <= 1'b0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_19 <= 1'b0;
      chn_inp_in_crt_sva_7_411_1 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_8_aelse_and_3_cse ) begin
      IsNaN_6U_10U_8_land_1_lpi_1_dfm_7 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_18,
          IsNaN_8U_23U_4_IsNaN_8U_23U_4_nand_tmp, and_dcpl_741);
      IsNaN_6U_10U_9_land_1_lpi_1_dfm_8 <= MUX_s_1_2_2(IsNaN_6U_10U_9_land_1_lpi_1_dfm_7,
          IsNaN_8U_23U_4_nor_tmp, and_dcpl_741);
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_19 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_18,
          IsNaN_6U_10U_8_land_1_lpi_1_dfm_st_3, and_dcpl_740);
      chn_inp_in_crt_sva_7_411_1 <= MUX_s_1_2_2(chn_inp_in_crt_sva_6_411_1, (FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_mx0[23]),
          and_dcpl_740);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_1_itm <= 10'b0;
    end
    else if ( core_wen & (~(nand_557_cse | (cfg_precision_1_sva_st_84[0]) | (chn_inp_in_crt_sva_7_739_736_1[1])
        | and_dcpl_78 | IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_5)) ) begin
      FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_1_itm <= FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_1_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_2_itm <= 10'b0;
    end
    else if ( core_wen & (~((~ main_stage_v_7) | IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_5
        | (cfg_precision_1_sva_st_84!=2'b10) | and_dcpl_78 | (chn_inp_in_crt_sva_7_739_736_1[2])))
        ) begin
      FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_2_itm <= FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_2_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_3_itm <= 10'b0;
    end
    else if ( core_wen & (~(or_dcpl_336 | (~ (cfg_precision_1_sva_st_84[1])) | (chn_inp_in_crt_sva_7_739_736_1[3])
        | and_dcpl_78 | IsNaN_6U_10U_8_land_lpi_1_dfm_st_5)) ) begin
      FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_3_itm <= FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_3_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpMantRNE_24U_11U_else_and_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_342 | (~ (chn_inp_in_crt_sva_6_739_736_1[0]))
        | (~ (cfg_precision_1_sva_st_83[1])) | (~ inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8)
        | inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7 | (~ inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8)
        | and_dcpl_78)) ) begin
      inp_lookup_1_FpMantRNE_24U_11U_else_and_svs <= inp_lookup_1_FpMantRNE_24U_11U_else_and_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_342 | (~ (chn_inp_in_crt_sva_6_739_736_1[0]))
        | (~ (cfg_precision_1_sva_st_83[1])) | and_dcpl_78 | (~ inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8)))
        ) begin
      inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
          <= inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpMantRNE_24U_11U_else_and_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_357 | (cfg_precision_1_sva_st_83!=2'b10) | (~
        inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8) | inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7
        | (~ inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8) | and_dcpl_78))
        ) begin
      inp_lookup_2_FpMantRNE_24U_11U_else_and_svs <= inp_lookup_2_FpMantRNE_24U_11U_else_and_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_357 | (cfg_precision_1_sva_st_83!=2'b10) | and_dcpl_78
        | (~ inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8))) ) begin
      inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
          <= inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpMantRNE_24U_11U_else_and_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_342 | (~ (cfg_precision_1_sva_st_83[1])) | (~
        (chn_inp_in_crt_sva_6_739_736_1[2])) | (~ inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8)
        | inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7 | (~ inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8)
        | and_dcpl_78)) ) begin
      inp_lookup_3_FpMantRNE_24U_11U_else_and_svs <= inp_lookup_3_FpMantRNE_24U_11U_else_and_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_342 | (~ (cfg_precision_1_sva_st_83[1])) | (~
        (chn_inp_in_crt_sva_6_739_736_1[2])) | and_dcpl_78 | (~ inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8)))
        ) begin
      inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
          <= inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2 <= 23'b0;
    end
    else if ( core_wen & (FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx0c0 | FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx0c1
        | FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx0c2) ) begin
      FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2 <= MUX1HOT_v_23_3_2(reg_chn_inp_in_crt_sva_6_94_64_1_reg,
          FpAdd_8U_23U_1_asn_40_mx0w1, reg_chn_inp_in_crt_sva_5_94_64_1_itm, {FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx0c0
          , FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx0c1 , FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_2_mx0c2});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpMantRNE_24U_11U_else_and_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_342 | (~ (cfg_precision_1_sva_st_83[1])) | (~
        (chn_inp_in_crt_sva_6_739_736_1[3])) | (~ inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8)
        | inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7 | (~ inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8)
        | and_dcpl_78)) ) begin
      inp_lookup_4_FpMantRNE_24U_11U_else_and_svs <= inp_lookup_4_FpMantRNE_24U_11U_else_and_svs_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_342 | (~ (cfg_precision_1_sva_st_83[1])) | (~
        (chn_inp_in_crt_sva_6_739_736_1[3])) | and_dcpl_78 | (~ inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8)))
        ) begin
      inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
          <= inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpAdd_6U_10U_1_is_a_greater_oif_equal_svs <= 1'b0;
    end
    else if ( core_wen & (~((cfg_precision_1_sva_st_81!=2'b10) | FpAdd_6U_10U_1_is_a_greater_acc_itm_6
        | (chn_inp_in_crt_sva_4_739_736_1[0]) | or_dcpl_409)) ) begin
      inp_lookup_1_FpAdd_6U_10U_1_is_a_greater_oif_equal_svs <= inp_lookup_1_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpAdd_6U_10U_1_is_a_greater_oif_equal_svs <= 1'b0;
    end
    else if ( core_wen & (~((cfg_precision_1_sva_st_81!=2'b10) | FpAdd_6U_10U_1_is_a_greater_acc_1_itm_6
        | (chn_inp_in_crt_sva_4_739_736_1[1]) | or_dcpl_409)) ) begin
      inp_lookup_2_FpAdd_6U_10U_1_is_a_greater_oif_equal_svs <= inp_lookup_2_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpAdd_6U_10U_1_is_a_greater_oif_equal_svs <= 1'b0;
    end
    else if ( core_wen & (~((cfg_precision_1_sva_st_81!=2'b10) | FpAdd_6U_10U_1_is_a_greater_acc_2_itm_6
        | (chn_inp_in_crt_sva_4_739_736_1[2]) | or_dcpl_409)) ) begin
      inp_lookup_3_FpAdd_6U_10U_1_is_a_greater_oif_equal_svs <= inp_lookup_3_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpAdd_6U_10U_1_is_a_greater_oif_equal_svs <= 1'b0;
    end
    else if ( core_wen & (~((cfg_precision_1_sva_st_81!=2'b10) | FpAdd_6U_10U_1_is_a_greater_acc_3_itm_6_1
        | (chn_inp_in_crt_sva_4_739_736_1[3]) | or_dcpl_409)) ) begin
      inp_lookup_4_FpAdd_6U_10U_1_is_a_greater_oif_equal_svs <= inp_lookup_4_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpMantWidthDec_6U_21U_10U_0U_0U_1_overflow_slc_FpMantRNE_22U_11U_i_data_1_20_1_19_10_itm
          <= 10'b0;
    end
    else if ( core_wen & ((~((mux_1919_nl) | (fsm_output[0]))) | and_dcpl_458 | and_dcpl_453)
        ) begin
      inp_lookup_1_FpMantWidthDec_6U_21U_10U_0U_0U_1_overflow_slc_FpMantRNE_22U_11U_i_data_1_20_1_19_10_itm
          <= MUX_v_10_2_2((FpMul_6U_10U_1_p_mant_20_1_1_lpi_1_dfm_3_mx0[19:10]),
          (FpMul_6U_10U_2_p_mant_20_1_1_lpi_1_dfm_3_mx0[19:10]), and_dcpl_453);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_22U_11U_1_else_carry_1_sva_1 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_458 | and_1468_rgt | and_1471_rgt) & (~ (mux_865_nl))
        ) begin
      FpMantRNE_22U_11U_1_else_carry_1_sva_1 <= MUX1HOT_s_1_3_2(FpMantRNE_22U_11U_1_else_carry_1_sva,
          FpMantRNE_22U_11U_2_else_carry_1_sva_mx1w1, FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_7_1_1,
          {and_dcpl_458 , and_1468_rgt , and_1471_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_8_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_10 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_31_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_8_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_7_1_1,
          FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_3_4_mx0w0, and_dcpl_458);
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_10 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_9,
          FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_3_3_0_mx0w0, and_dcpl_458);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_8_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_10 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_33_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_8_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_7_1_1,
          FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_3_4_mx0w0, and_dcpl_495);
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_10 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_9,
          FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_3_3_0_mx0w0, and_dcpl_495);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_22U_11U_1_else_carry_3_sva_1 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_530 | and_1474_rgt | and_1477_rgt) & (~ (mux_899_nl))
        ) begin
      FpMantRNE_22U_11U_1_else_carry_3_sva_1 <= MUX1HOT_s_1_3_2(FpMantRNE_22U_11U_1_else_carry_3_sva,
          FpMantRNE_22U_11U_2_else_carry_3_sva_mx1w1, FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_7_1_1,
          {and_dcpl_530 , and_1474_rgt , and_1477_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpMantWidthDec_6U_21U_10U_0U_0U_1_overflow_slc_FpMantRNE_22U_11U_i_data_1_20_1_19_10_itm
          <= 10'b0;
    end
    else if ( core_wen & ((~ or_tmp_4457) | and_dcpl_1007 | and_dcpl_1009) ) begin
      inp_lookup_4_FpMantWidthDec_6U_21U_10U_0U_0U_1_overflow_slc_FpMantRNE_22U_11U_i_data_1_20_1_19_10_itm
          <= MUX_v_10_2_2((FpMul_6U_10U_1_p_mant_20_1_lpi_1_dfm_3_mx0[19:10]), (FpMul_6U_10U_2_p_mant_20_1_lpi_1_dfm_3_mx0[19:10]),
          and_dcpl_1009);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_8_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_8_0 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_10 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_and_37_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_8_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_7_1_1,
          FpMul_6U_10U_2_o_expo_lpi_1_dfm_3_5_mx0w0, and_dcpl_1007);
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_8_0 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_7_0_1,
          FpMul_6U_10U_2_o_expo_lpi_1_dfm_3_4_mx0w0, and_dcpl_1007);
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_10 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_9,
          FpMul_6U_10U_2_o_expo_lpi_1_dfm_3_3_0_mx0w0, and_dcpl_1007);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_7_itm <= 2'b0;
    end
    else if ( core_wen & (cfg_precision_1_sva_st_90[1]) & or_11_cse & (~ (cfg_precision_1_sva_st_90[0]))
        & main_stage_v_1 & (~ (chn_inp_in_crt_sva_1_739_395_1[343])) ) begin
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_7_itm <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_mux1h_4_itm[9:8];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_7_1_itm <= 8'b0;
    end
    else if ( core_wen & (cfg_precision_1_sva_st_90==2'b10) & or_11_cse & main_stage_v_1
        ) begin
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_7_1_itm <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_mux1h_4_itm[7:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_8 <= 10'b0;
    end
    else if ( core_wen & (and_1537_rgt | and_1538_rgt | and_dcpl_145) & mux_tmp_6
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_8 <= MUX1HOT_v_10_3_2((chn_inp_in_rsci_d_mxwt[341:332]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_or_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_3, {and_1537_rgt ,
          and_1538_rgt , and_dcpl_145});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_8 <= 10'b0;
    end
    else if ( core_wen & (and_1588_rgt | and_1589_rgt | and_dcpl_215) & mux_tmp_6
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_8 <= MUX1HOT_v_10_3_2((chn_inp_in_rsci_d_mxwt[357:348]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_or_4_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_3, {and_1588_rgt ,
          and_1589_rgt , and_dcpl_215});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_3_lpi_1_dfm_8 <= 10'b0;
    end
    else if ( core_wen & (and_1639_rgt | and_1640_rgt | and_dcpl_285) & mux_tmp_6
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_3_lpi_1_dfm_8 <= MUX1HOT_v_10_3_2((chn_inp_in_rsci_d_mxwt[373:364]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_or_8_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_3_lpi_1_dfm_3, {and_1639_rgt ,
          and_1640_rgt , and_dcpl_285});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_8 <= 10'b0;
    end
    else if ( core_wen & (and_1690_rgt | and_1691_rgt | and_dcpl_355) & mux_tmp_6
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_8 <= MUX1HOT_v_10_3_2((chn_inp_in_rsci_d_mxwt[389:380]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_or_12_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_3, {and_1690_rgt , and_1691_rgt
          , and_dcpl_355});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_35U_1_leading_sign_35_0_rtn_1_sva <= 6'b0;
      inp_lookup_1_FpMantRNE_36U_11U_1_else_and_svs <= 1'b0;
    end
    else if ( IntLeadZero_35U_1_leading_sign_35_0_rtn_and_cse ) begin
      IntLeadZero_35U_1_leading_sign_35_0_rtn_1_sva <= libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_12;
      inp_lookup_1_FpMantRNE_36U_11U_1_else_and_svs <= inp_lookup_1_FpMantRNE_36U_11U_1_else_and_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_35U_1_leading_sign_35_0_rtn_2_sva <= 6'b0;
      inp_lookup_2_FpMantRNE_36U_11U_1_else_and_svs <= 1'b0;
    end
    else if ( IntLeadZero_35U_1_leading_sign_35_0_rtn_and_1_cse ) begin
      IntLeadZero_35U_1_leading_sign_35_0_rtn_2_sva <= libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_13;
      inp_lookup_2_FpMantRNE_36U_11U_1_else_and_svs <= inp_lookup_2_FpMantRNE_36U_11U_1_else_and_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_35U_1_leading_sign_35_0_rtn_3_sva <= 6'b0;
      inp_lookup_3_FpMantRNE_36U_11U_1_else_and_svs <= 1'b0;
    end
    else if ( IntLeadZero_35U_1_leading_sign_35_0_rtn_and_2_cse ) begin
      IntLeadZero_35U_1_leading_sign_35_0_rtn_3_sva <= libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_14;
      inp_lookup_3_FpMantRNE_36U_11U_1_else_and_svs <= inp_lookup_3_FpMantRNE_36U_11U_1_else_and_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntLeadZero_35U_1_leading_sign_35_0_rtn_sva <= 6'b0;
      inp_lookup_4_FpMantRNE_36U_11U_1_else_and_svs <= 1'b0;
    end
    else if ( IntLeadZero_35U_1_leading_sign_35_0_rtn_and_3_cse ) begin
      IntLeadZero_35U_1_leading_sign_35_0_rtn_sva <= libraries_leading_sign_35_0_ac2f757814855ba106465f8cb39af0da6a26_15;
      inp_lookup_4_FpMantRNE_36U_11U_1_else_and_svs <= inp_lookup_4_FpMantRNE_36U_11U_1_else_and_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3 <=
          1'b0;
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_land_2_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_2_land_2_lpi_1_dfm_st_6 <= 1'b0;
      inp_lookup_2_IsZero_6U_10U_1_aif_IsZero_6U_10U_1_aelse_nor_itm_2 <= 1'b0;
      inp_lookup_2_IsZero_6U_10U_2_aif_IsZero_6U_10U_2_aelse_nor_itm_2 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_is_addition_and_9_cse ) begin
      inp_lookup_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3 <=
          ~((chn_inp_in_rsci_d_mxwt[543]) ^ (chn_inp_in_rsci_d_mxwt[671]));
      IsNaN_8U_23U_1_land_2_lpi_1_dfm_4 <= ~((~((chn_inp_in_rsci_d_mxwt[662:640]!=23'b00000000000000000000000)))
          | (chn_inp_in_rsci_d_mxwt[670:663]!=8'b11111111));
      IsNaN_8U_23U_land_2_lpi_1_dfm_4 <= ~((~((chn_inp_in_rsci_d_mxwt[534:512]!=23'b00000000000000000000000)))
          | (chn_inp_in_rsci_d_mxwt[542:535]!=8'b11111111));
      IsNaN_8U_23U_2_land_2_lpi_1_dfm_st_6 <= ~((~((chn_inp_in_rsci_d_mxwt[54:32]!=23'b00000000000000000000000)))
          | (chn_inp_in_rsci_d_mxwt[62:55]!=8'b11111111));
      inp_lookup_2_IsZero_6U_10U_1_aif_IsZero_6U_10U_1_aelse_nor_itm_2 <= ~((FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_3_mx1!=10'b0000000000));
      inp_lookup_2_IsZero_6U_10U_2_aif_IsZero_6U_10U_2_aelse_nor_itm_2 <= inp_lookup_2_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3 <=
          1'b0;
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_land_3_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_2_land_3_lpi_1_dfm_st_6 <= 1'b0;
      inp_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_5 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_is_addition_and_10_cse ) begin
      inp_lookup_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3 <=
          ~((chn_inp_in_rsci_d_mxwt[575]) ^ (chn_inp_in_rsci_d_mxwt[703]));
      IsNaN_8U_23U_1_land_3_lpi_1_dfm_4 <= ~((~((chn_inp_in_rsci_d_mxwt[694:672]!=23'b00000000000000000000000)))
          | (chn_inp_in_rsci_d_mxwt[702:695]!=8'b11111111));
      IsNaN_8U_23U_land_3_lpi_1_dfm_4 <= ~((~((chn_inp_in_rsci_d_mxwt[566:544]!=23'b00000000000000000000000)))
          | (chn_inp_in_rsci_d_mxwt[574:567]!=8'b11111111));
      IsNaN_8U_23U_2_land_3_lpi_1_dfm_st_6 <= ~((~((chn_inp_in_rsci_d_mxwt[86:64]!=23'b00000000000000000000000)))
          | (chn_inp_in_rsci_d_mxwt[94:87]!=8'b11111111));
      inp_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_5 <= (chn_inp_in_rsci_d_mxwt[94:64]!=31'b0000000000000000000000000000000);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3 <=
          1'b0;
      IsNaN_8U_23U_1_land_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_land_lpi_1_dfm_4 <= 1'b0;
      IsNaN_8U_23U_2_land_lpi_1_dfm_st_6 <= 1'b0;
      inp_lookup_4_IsZero_6U_10U_1_aif_IsZero_6U_10U_1_aelse_nor_itm_2 <= 1'b0;
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_13 <= 1'b0;
      inp_lookup_4_IsZero_6U_10U_2_aif_IsZero_6U_10U_2_aelse_nor_itm_2 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_is_addition_and_11_cse ) begin
      inp_lookup_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_3 <=
          ~((chn_inp_in_rsci_d_mxwt[607]) ^ (chn_inp_in_rsci_d_mxwt[735]));
      IsNaN_8U_23U_1_land_lpi_1_dfm_4 <= ~((~((chn_inp_in_rsci_d_mxwt[726:704]!=23'b00000000000000000000000)))
          | (chn_inp_in_rsci_d_mxwt[734:727]!=8'b11111111));
      IsNaN_8U_23U_land_lpi_1_dfm_4 <= ~((~((chn_inp_in_rsci_d_mxwt[598:576]!=23'b00000000000000000000000)))
          | (chn_inp_in_rsci_d_mxwt[606:599]!=8'b11111111));
      IsNaN_8U_23U_2_land_lpi_1_dfm_st_6 <= ~((~((chn_inp_in_rsci_d_mxwt[118:96]!=23'b00000000000000000000000)))
          | (chn_inp_in_rsci_d_mxwt[126:119]!=8'b11111111));
      inp_lookup_4_IsZero_6U_10U_1_aif_IsZero_6U_10U_1_aelse_nor_itm_2 <= ~((FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_3_mx1!=10'b0000000000));
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_13 <= IsNaN_6U_10U_2_land_lpi_1_dfm_mx0w0;
      inp_lookup_4_IsZero_6U_10U_2_aif_IsZero_6U_10U_2_aelse_nor_itm_2 <= inp_lookup_4_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2 <= 1'b0;
      inp_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_2 <= 1'b0;
    end
    else if ( IsZero_8U_23U_1_and_cse ) begin
      inp_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2 <= (chn_inp_in_rsci_d_mxwt[638:608]!=31'b0000000000000000000000000000000);
      inp_lookup_1_FpAdd_8U_23U_IsZero_8U_23U_or_itm_2 <= (chn_inp_in_rsci_d_mxwt[510:480]!=31'b0000000000000000000000000000000);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_922_nl)) ) begin
      inp_lookup_2_FpAdd_8U_23U_IsZero_8U_23U_or_itm_2 <= (chn_inp_in_rsci_d_mxwt[542:512]!=31'b0000000000000000000000000000000);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2 <= 1'b0;
      inp_lookup_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_2 <= 1'b0;
    end
    else if ( IsZero_8U_23U_1_and_1_cse ) begin
      inp_lookup_3_FpAdd_8U_23U_IsZero_8U_23U_1_or_itm_2 <= (chn_inp_in_rsci_d_mxwt[702:672]!=31'b0000000000000000000000000000000);
      inp_lookup_3_FpAdd_8U_23U_IsZero_8U_23U_or_itm_2 <= (chn_inp_in_rsci_d_mxwt[574:544]!=31'b0000000000000000000000000000000);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_924_nl)) ) begin
      inp_lookup_4_FpAdd_8U_23U_IsZero_8U_23U_or_itm_2 <= (chn_inp_in_rsci_d_mxwt[606:576]!=31'b0000000000000000000000000000000);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_2_606_576_itm <= 12'b0;
    end
    else if ( or_5695_itm & core_wen & main_stage_v_1 & (cfg_precision_1_sva_st_90==2'b10)
        & (chn_inp_in_crt_sva_1_739_395_1[344]) & or_11_cse ) begin
      reg_chn_inp_in_crt_sva_2_606_576_itm <= mux1h_34_itm[30:19];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_2_606_576_1_itm <= 19'b0;
    end
    else if ( (~ (mux_2106_nl)) & and_dcpl_2318 & or_11_cse ) begin
      reg_chn_inp_in_crt_sva_2_606_576_1_itm <= mux1h_34_itm[18:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_2_574_544_itm <= 12'b0;
    end
    else if ( or_5694_itm & core_wen & main_stage_v_1 & (chn_inp_in_crt_sva_1_739_395_1[343])
        & (cfg_precision_1_sva_st_90==2'b10) & or_11_cse ) begin
      reg_chn_inp_in_crt_sva_2_574_544_itm <= mux1h_36_itm[30:19];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_2_574_544_1_itm <= 19'b0;
    end
    else if ( (~ (mux_2109_nl)) & and_dcpl_2318 & or_11_cse ) begin
      reg_chn_inp_in_crt_sva_2_574_544_1_itm <= mux1h_36_itm[18:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_2_510_480_itm <= 12'b0;
    end
    else if ( or_6042_cse & core_wen & (chn_inp_in_crt_sva_1_739_395_1[341]) & main_stage_v_1
        & (cfg_precision_1_sva_st_90==2'b10) & or_11_cse ) begin
      reg_chn_inp_in_crt_sva_2_510_480_itm <= mux1h_38_itm[30:19];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_2_510_480_1_itm <= 19'b0;
    end
    else if ( (~ (mux_2113_nl)) & and_dcpl_2318 & or_11_cse ) begin
      reg_chn_inp_in_crt_sva_2_510_480_1_itm <= mux1h_38_itm[18:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_2_542_512_itm <= 12'b0;
    end
    else if ( or_5693_itm & core_wen & main_stage_v_1 & (cfg_precision_1_sva_st_90==2'b10)
        & (chn_inp_in_crt_sva_1_739_395_1[342]) & or_11_cse ) begin
      reg_chn_inp_in_crt_sva_2_542_512_itm <= mux1h_40_itm[30:19];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_2_542_512_1_itm <= 19'b0;
    end
    else if ( (~ (mux_2116_nl)) & and_dcpl_2318 & or_11_cse ) begin
      reg_chn_inp_in_crt_sva_2_542_512_1_itm <= mux1h_40_itm[18:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSignedShiftRight_50U_5U_32U_mbits_fixed_1_sva_1_80_14_1 <= 67'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_939_nl) ) begin
      IntSignedShiftRight_50U_5U_32U_mbits_fixed_1_sva_1_80_14_1 <= IntSignedShiftRight_50U_5U_32U_mbits_fixed_1_sva[80:14];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_p_mant_p1_1_sva <= 22'b0;
    end
    else if ( FpAdd_8U_23U_o_expo_and_cse & inp_lookup_1_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs
        & (~(or_dcpl_159 | and_dcpl_78 | FpMul_6U_10U_2_lor_6_lpi_1_dfm_st_3)) &
        (mux_118_nl) ) begin
      FpMul_6U_10U_2_p_mant_p1_1_sva <= inp_lookup_1_FpMul_6U_10U_2_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_7_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_10 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_24_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_7_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_6_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_10 <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_7_0_1 <= 1'b0;
    end
    else if ( core_wen & FpFractionToFloat_35U_6U_10U_is_zero_FpFractionToFloat_35U_6U_10U_is_zero_or_3_cse
        & (mux_123_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_7_0_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_6_0_1,
          inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_mx0w1,
          and_dcpl_394);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSignedShiftRight_50U_5U_32U_mbits_fixed_2_sva_1_80_14_1 <= 67'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_941_nl) ) begin
      IntSignedShiftRight_50U_5U_32U_mbits_fixed_2_sva_1_80_14_1 <= IntSignedShiftRight_50U_5U_32U_mbits_fixed_2_sva[80:14];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_p_mant_p1_2_sva <= 22'b0;
    end
    else if ( FpAdd_8U_23U_o_expo_and_cse & inp_lookup_2_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs
        & (~(or_tmp_439 | FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_3 | (chn_inp_in_crt_sva_2_739_736_1[1])
        | or_dcpl_660)) & (mux_140_nl) ) begin
      FpMul_6U_10U_2_p_mant_p1_2_sva <= inp_lookup_2_FpMul_6U_10U_2_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_7_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_10 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_27_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_7_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_6_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_10 <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_7_0_1 <= 1'b0;
    end
    else if ( core_wen & FpFractionToFloat_35U_6U_10U_is_zero_FpFractionToFloat_35U_6U_10U_is_zero_or_2_cse
        & (mux_146_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_7_0_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_6_0_1,
          inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_mx0w1,
          and_dcpl_402);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSignedShiftRight_50U_5U_32U_mbits_fixed_3_sva_1_80_14_1 <= 67'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_943_nl) ) begin
      IntSignedShiftRight_50U_5U_32U_mbits_fixed_3_sva_1_80_14_1 <= IntSignedShiftRight_50U_5U_32U_mbits_fixed_3_sva[80:14];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_p_mant_p1_3_sva <= 22'b0;
    end
    else if ( FpAdd_8U_23U_o_expo_and_cse & inp_lookup_3_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs
        & (~(or_dcpl_167 | and_dcpl_78 | FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_3)) &
        (mux_163_nl) ) begin
      FpMul_6U_10U_2_p_mant_p1_3_sva <= inp_lookup_3_FpMul_6U_10U_2_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_7_0_1 <= 1'b0;
    end
    else if ( core_wen & FpFractionToFloat_35U_6U_10U_is_zero_FpFractionToFloat_35U_6U_10U_is_zero_or_1_cse
        & (mux_946_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_7_0_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_6_0_1,
          inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_mx0w1,
          and_dcpl_410);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSignedShiftRight_50U_5U_32U_mbits_fixed_sva_1_80_14_1 <= 67'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_947_nl) ) begin
      IntSignedShiftRight_50U_5U_32U_mbits_fixed_sva_1_80_14_1 <= IntSignedShiftRight_50U_5U_32U_mbits_fixed_sva[80:14];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_p_mant_p1_sva <= 22'b0;
    end
    else if ( FpAdd_8U_23U_o_expo_and_cse & inp_lookup_4_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs
        & (~(or_5809_cse | and_dcpl_78 | FpMul_6U_10U_2_lor_1_lpi_1_dfm_st_3)) &
        (mux_180_nl) ) begin
      FpMul_6U_10U_2_p_mant_p1_sva <= inp_lookup_4_FpMul_6U_10U_2_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_7_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_7_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_10 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_33_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_7_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_6_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_7_0_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_6_0_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_10 <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_lor_6_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & FpMul_6U_10U_2_oelse_1_FpMul_6U_10U_2_oelse_1_or_11_cse
        & (mux_951_nl) ) begin
      FpMul_6U_10U_1_lor_6_lpi_1_dfm_5 <= MUX_s_1_2_2(or_457_cse, FpNormalize_8U_49U_if_FpNormalize_8U_49U_if_nand_tmp,
          and_dcpl_427);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_5_land_1_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & (and_1717_rgt | and_1725_rgt | and_dcpl_427) & (~ mux_197_itm)
        ) begin
      IsNaN_6U_10U_5_land_1_lpi_1_dfm_5 <= MUX1HOT_s_1_3_2(and_3246_cse, IsNaN_6U_10U_5_land_1_lpi_1_dfm,
          FpFractionToFloat_35U_6U_10U_is_zero_1_lpi_1_dfm_5, {and_1717_rgt , and_1725_rgt
          , and_dcpl_427});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_lor_7_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_2_cse
        & (mux_954_nl) ) begin
      FpMul_6U_10U_1_lor_7_lpi_1_dfm_5 <= MUX_s_1_2_2(or_519_cse, FpNormalize_8U_49U_if_FpNormalize_8U_49U_if_nand_1_tmp,
          and_dcpl_464);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_5_land_2_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & (and_1726_rgt | and_1734_rgt | and_dcpl_464) & (~ mux_197_itm)
        ) begin
      IsNaN_6U_10U_5_land_2_lpi_1_dfm_5 <= MUX1HOT_s_1_3_2(and_3244_cse, IsNaN_6U_10U_5_land_2_lpi_1_dfm,
          FpFractionToFloat_35U_6U_10U_is_zero_2_lpi_1_dfm_5, {and_1726_rgt , and_1734_rgt
          , and_dcpl_464});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_lor_8_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_1_cse
        & (mux_957_nl) ) begin
      FpMul_6U_10U_1_lor_8_lpi_1_dfm_5 <= MUX_s_1_2_2(or_593_cse, FpNormalize_8U_49U_if_FpNormalize_8U_49U_if_nand_2_tmp,
          and_dcpl_496);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_5_land_3_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & (and_1735_rgt | and_1743_rgt | and_dcpl_496) & (~ mux_197_itm)
        ) begin
      IsNaN_6U_10U_5_land_3_lpi_1_dfm_5 <= MUX1HOT_s_1_3_2(and_3242_cse, IsNaN_6U_10U_5_land_3_lpi_1_dfm,
          FpFractionToFloat_35U_6U_10U_is_zero_3_lpi_1_dfm_5, {and_1735_rgt , and_1743_rgt
          , and_dcpl_496});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_lor_1_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_cse
        & (mux_960_nl) ) begin
      FpMul_6U_10U_1_lor_1_lpi_1_dfm_5 <= MUX_s_1_2_2(or_648_cse, FpNormalize_8U_49U_if_FpNormalize_8U_49U_if_nand_3_tmp,
          and_dcpl_535);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_5_land_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & (and_1744_rgt | and_1752_rgt | and_dcpl_535) & (~ mux_197_itm)
        ) begin
      IsNaN_6U_10U_5_land_lpi_1_dfm_5 <= MUX1HOT_s_1_3_2(and_3240_cse, IsNaN_6U_10U_5_land_lpi_1_dfm,
          FpFractionToFloat_35U_6U_10U_is_zero_lpi_1_dfm_5, {and_1744_rgt , and_1752_rgt
          , and_dcpl_535});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_427 | and_1754_rgt | and_1755_rgt) & (mux_962_nl)
        ) begin
      inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4
          <= MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_7_0_1,
          inp_lookup_1_FpMul_6U_10U_1_else_2_if_acc_itm_6_1, inp_lookup_1_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs,
          {and_dcpl_427 , and_1754_rgt , and_1755_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_464 | and_1757_rgt | and_1758_rgt) & (mux_964_nl)
        ) begin
      inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4
          <= MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_7_0_1,
          inp_lookup_2_FpMul_6U_10U_1_else_2_if_acc_itm_6_1, inp_lookup_2_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs,
          {and_dcpl_464 , and_1757_rgt , and_1758_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4
          <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_496 | and_1760_rgt | and_1761_rgt) & (mux_966_nl)
        ) begin
      inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4
          <= MUX1HOT_s_1_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_7_0_1,
          inp_lookup_3_FpMul_6U_10U_1_else_2_if_acc_itm_6_1, inp_lookup_3_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs,
          {and_dcpl_496 , and_1760_rgt , and_1761_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_p_mant_p1_1_sva <= 22'b0;
    end
    else if ( FpAdd_8U_23U_o_expo_and_cse & inp_lookup_1_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs
        & (~(FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_3 | (cfg_precision_1_sva_st_80!=2'b10)
        | (chn_inp_in_crt_sva_3_739_736_1[0]) | or_dcpl_699)) & (mux_210_nl) ) begin
      FpMul_6U_10U_1_p_mant_p1_1_sva <= inp_lookup_1_FpMul_6U_10U_1_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_else_2_else_and_itm_2 <= 1'b0;
    end
    else if ( core_wen & FpMul_6U_10U_2_oelse_1_FpMul_6U_10U_2_oelse_1_or_11_cse
        & (~ (mux_970_nl)) ) begin
      FpMul_6U_10U_2_else_2_else_and_itm_2 <= MUX_s_1_2_2((FpMul_6U_10U_2_else_2_else_and_nl),
          IsZero_6U_10U_1_IsZero_6U_10U_1_and_itm_8, and_dcpl_427);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_7_4_0_1 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_971_nl) ) begin
      FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_7_4_0_1 <= FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_6_4_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_972_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_11 <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_7_land_1_lpi_1_dfm_6 <= 1'b0;
      IsNaN_6U_10U_7_land_2_lpi_1_dfm_6 <= 1'b0;
      IsNaN_6U_10U_7_land_3_lpi_1_dfm_6 <= 1'b0;
      IsNaN_6U_10U_7_land_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_7_aelse_and_4_cse ) begin
      IsNaN_6U_10U_7_land_1_lpi_1_dfm_6 <= IsNaN_6U_10U_7_land_1_lpi_1_dfm_5;
      IsNaN_6U_10U_7_land_2_lpi_1_dfm_6 <= IsNaN_6U_10U_7_land_2_lpi_1_dfm_5;
      IsNaN_6U_10U_7_land_3_lpi_1_dfm_6 <= IsNaN_6U_10U_7_land_3_lpi_1_dfm_5;
      IsNaN_6U_10U_7_land_lpi_1_dfm_6 <= IsNaN_6U_10U_7_land_lpi_1_dfm_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_lor_6_lpi_1_dfm_6 <= 1'b0;
      FpMul_6U_10U_2_FpMul_6U_10U_2_and_itm_2 <= 1'b0;
    end
    else if ( FpMul_6U_10U_2_oelse_1_and_8_cse ) begin
      FpMul_6U_10U_2_lor_6_lpi_1_dfm_6 <= MUX_s_1_2_2(FpMul_6U_10U_2_lor_6_lpi_1_dfm_5,
          chn_inp_in_crt_sva_2_347_1, and_dcpl_427);
      FpMul_6U_10U_2_FpMul_6U_10U_2_and_itm_2 <= MUX_s_1_2_2((FpMul_6U_10U_2_FpMul_6U_10U_2_and_nl),
          IsNaN_8U_23U_land_1_lpi_1_dfm_st_4, and_dcpl_427);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_p_mant_p1_2_sva <= 22'b0;
    end
    else if ( FpAdd_8U_23U_o_expo_and_cse & inp_lookup_2_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs
        & (~(or_tmp_440 | FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_3 | (chn_inp_in_crt_sva_3_739_736_1[1])
        | or_dcpl_699)) & (mux_248_nl) ) begin
      FpMul_6U_10U_1_p_mant_p1_2_sva <= inp_lookup_2_FpMul_6U_10U_1_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_else_2_else_ac_int_cctor_2_sva_2 <= 6'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_976_nl) ) begin
      FpMul_6U_10U_2_else_2_else_ac_int_cctor_2_sva_2 <= FpMul_6U_10U_2_else_2_else_ac_int_cctor_2_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_else_2_else_and_1_itm_2 <= 1'b0;
    end
    else if ( core_wen & IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_2_cse
        & (~ (mux_980_nl)) ) begin
      FpMul_6U_10U_2_else_2_else_and_1_itm_2 <= MUX_s_1_2_2((FpMul_6U_10U_2_else_2_else_and_1_nl),
          IsZero_6U_10U_1_IsZero_6U_10U_1_and_1_itm_6, and_dcpl_464);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_7_4_0_1 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_981_nl) ) begin
      FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_7_4_0_1 <= FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_6_4_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_982_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_11 <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_lor_7_lpi_1_dfm_6 <= 1'b0;
      FpMul_6U_10U_2_FpMul_6U_10U_2_and_16_itm_2 <= 1'b0;
    end
    else if ( FpMul_6U_10U_2_oelse_1_and_9_cse ) begin
      FpMul_6U_10U_2_lor_7_lpi_1_dfm_6 <= MUX_s_1_2_2(FpMul_6U_10U_2_lor_7_lpi_1_dfm_5,
          chn_inp_in_crt_sva_2_363_1, and_dcpl_464);
      FpMul_6U_10U_2_FpMul_6U_10U_2_and_16_itm_2 <= MUX_s_1_2_2((FpMul_6U_10U_2_FpMul_6U_10U_2_and_16_nl),
          IsNaN_8U_23U_land_2_lpi_1_dfm_st_4, and_dcpl_464);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_p_mant_p1_3_sva <= 22'b0;
    end
    else if ( FpAdd_8U_23U_o_expo_and_cse & inp_lookup_3_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs
        & (~(or_tmp_440 | FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_3 | (chn_inp_in_crt_sva_3_739_736_1[2])
        | or_dcpl_699)) & (mux_286_nl) ) begin
      FpMul_6U_10U_1_p_mant_p1_3_sva <= inp_lookup_3_FpMul_6U_10U_1_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_else_2_else_ac_int_cctor_3_sva_2 <= 6'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_986_nl) ) begin
      FpMul_6U_10U_2_else_2_else_ac_int_cctor_3_sva_2 <= FpMul_6U_10U_2_else_2_else_ac_int_cctor_3_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_else_2_else_and_2_itm_2 <= 1'b0;
    end
    else if ( core_wen & IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_1_cse
        & (~ (mux_990_nl)) ) begin
      FpMul_6U_10U_2_else_2_else_and_2_itm_2 <= MUX_s_1_2_2((FpMul_6U_10U_2_else_2_else_and_2_nl),
          IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_itm_8, and_dcpl_496);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_7_4_0_1 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_991_nl) ) begin
      FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_7_4_0_1 <= FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_6_4_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_3_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_992_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_3_lpi_1_dfm_11 <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_3_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_lor_8_lpi_1_dfm_6 <= 1'b0;
      FpMul_6U_10U_2_FpMul_6U_10U_2_and_17_itm_2 <= 1'b0;
    end
    else if ( FpMul_6U_10U_2_oelse_1_and_10_cse ) begin
      FpMul_6U_10U_2_lor_8_lpi_1_dfm_6 <= MUX_s_1_2_2(FpMul_6U_10U_2_lor_8_lpi_1_dfm_5,
          chn_inp_in_crt_sva_2_379_1, and_dcpl_496);
      FpMul_6U_10U_2_FpMul_6U_10U_2_and_17_itm_2 <= MUX_s_1_2_2((FpMul_6U_10U_2_FpMul_6U_10U_2_and_17_nl),
          IsNaN_8U_23U_land_3_lpi_1_dfm_st_4, and_dcpl_496);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_p_mant_p1_sva <= 22'b0;
    end
    else if ( FpAdd_8U_23U_o_expo_and_cse & inp_lookup_4_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs
        & (~(or_dcpl_186 | and_dcpl_78 | FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_3)) &
        (mux_336_nl) ) begin
      FpMul_6U_10U_1_p_mant_p1_sva <= inp_lookup_4_FpMul_6U_10U_1_p_mant_p1_mul_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_else_2_else_and_3_itm_2 <= 1'b0;
    end
    else if ( core_wen & IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_cse
        & (~ (mux_1001_nl)) ) begin
      FpMul_6U_10U_2_else_2_else_and_3_itm_2 <= MUX_s_1_2_2((FpMul_6U_10U_2_else_2_else_and_3_nl),
          IsZero_6U_10U_1_IsZero_6U_10U_1_and_3_itm_6, and_dcpl_535);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_7_4_0_1 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1002_nl) ) begin
      FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_7_4_0_1 <= FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_6_4_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_11 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1003_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_11 <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_lor_1_lpi_1_dfm_6 <= 1'b0;
      FpMul_6U_10U_2_FpMul_6U_10U_2_and_18_itm_2 <= 1'b0;
    end
    else if ( FpMul_6U_10U_2_oelse_1_and_11_cse ) begin
      FpMul_6U_10U_2_lor_1_lpi_1_dfm_6 <= MUX_s_1_2_2(FpMul_6U_10U_2_lor_1_lpi_1_dfm_5,
          chn_inp_in_crt_sva_2_395_1, and_dcpl_535);
      FpMul_6U_10U_2_FpMul_6U_10U_2_and_18_itm_2 <= MUX_s_1_2_2((FpMul_6U_10U_2_FpMul_6U_10U_2_and_18_nl),
          IsNaN_8U_23U_land_lpi_1_dfm_st_4, and_dcpl_535);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs_2
          <= 1'b0;
    end
    else if ( core_wen & ((or_11_cse & (~(FpMul_6U_10U_1_if_2_FpMul_6U_10U_1_if_2_or_6_tmp
        | inp_lookup_4_FpMul_6U_10U_1_oelse_1_acc_itm_7_1))) | and_1764_rgt) & (mux_1006_nl)
        ) begin
      inp_lookup_4_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs_2
          <= MUX_s_1_2_2(inp_lookup_4_FpMul_6U_10U_1_else_2_if_acc_itm_6_1, inp_lookup_4_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs,
          and_1764_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_8U_23U_o_expo_1_lpi_1_dfm_11_reg <= 2'b0;
    end
    else if ( or_11_cse & core_wen & (chn_inp_in_crt_sva_3_739_736_1[0]) ) begin
      reg_FpAdd_8U_23U_o_expo_1_lpi_1_dfm_11_reg <= FpAdd_8U_23U_o_expo_FpAdd_8U_23U_o_expo_mux_rgt[7:6];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_or_6_cse
        & (mux_1011_nl) ) begin
      FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_1_mx0w0,
          (FpMul_6U_10U_1_else_2_else_and_nl), and_dcpl_565);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1014_nl) ) begin
      inp_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2 <= (FpAdd_8U_23U_o_mant_1_lpi_1_dfm_2_mx2!=23'b00000000000000000000000)
          | (FpAdd_8U_23U_o_expo_1_lpi_1_dfm_7_mx1w1!=8'b00000000);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_o_mant_1_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((or_11_cse & IsNaN_6U_10U_6_land_1_lpi_1_dfm_5) | and_1768_rgt)
        & (mux_1017_nl) ) begin
      FpAdd_8U_23U_o_mant_1_lpi_1_dfm_6 <= MUX_v_23_2_2(reg_chn_inp_in_crt_sva_3_510_480_1_reg,
          FpAdd_8U_23U_FpAdd_8U_23U_or_4_itm, and_4218_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_7 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_or_6_cse
        & (mux_1022_nl) ) begin
      inp_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_7 <= MUX_s_1_2_2(inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4,
          (inp_lookup_1_FpMul_6U_10U_1_p_mant_p1_mul_tmp[21]), and_dcpl_565);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_8U_23U_o_expo_2_lpi_1_dfm_11_reg <= 2'b0;
    end
    else if ( or_11_cse & core_wen & (chn_inp_in_crt_sva_3_739_736_1[1]) ) begin
      reg_FpAdd_8U_23U_o_expo_2_lpi_1_dfm_11_reg <= FpAdd_8U_23U_o_expo_FpAdd_8U_23U_o_expo_mux_1_rgt[7:6];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_or_5_cse
        & (mux_1027_nl) ) begin
      FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_1_mx0w0,
          (FpMul_6U_10U_1_else_2_else_and_1_nl), and_dcpl_583);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1030_nl) ) begin
      inp_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2 <= (FpAdd_8U_23U_o_mant_2_lpi_1_dfm_2_mx2!=23'b00000000000000000000000)
          | (FpAdd_8U_23U_o_expo_2_lpi_1_dfm_7_mx1w1!=8'b00000000);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_o_mant_2_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((or_11_cse & IsNaN_6U_10U_6_land_2_lpi_1_dfm_5) | and_1772_rgt)
        & (mux_1033_nl) ) begin
      FpAdd_8U_23U_o_mant_2_lpi_1_dfm_6 <= MUX_v_23_2_2(reg_chn_inp_in_crt_sva_3_542_512_1_reg,
          FpAdd_8U_23U_FpAdd_8U_23U_or_5_itm, and_4217_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_6 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_or_5_cse
        & (mux_1038_nl) ) begin
      inp_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_6 <= MUX_s_1_2_2(inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4,
          (inp_lookup_2_FpMul_6U_10U_1_p_mant_p1_mul_tmp[21]), and_dcpl_583);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_8U_23U_o_expo_3_lpi_1_dfm_11_reg <= 2'b0;
    end
    else if ( or_11_cse & core_wen & (chn_inp_in_crt_sva_3_739_736_1[2]) ) begin
      reg_FpAdd_8U_23U_o_expo_3_lpi_1_dfm_11_reg <= FpAdd_8U_23U_o_expo_FpAdd_8U_23U_o_expo_mux_2_rgt[7:6];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_or_4_cse
        & (mux_1043_nl) ) begin
      FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_1_mx0w0,
          (FpMul_6U_10U_1_else_2_else_and_2_nl), and_dcpl_601);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1046_nl) ) begin
      inp_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2 <= (FpAdd_8U_23U_o_mant_3_lpi_1_dfm_2_mx2!=23'b00000000000000000000000)
          | (FpAdd_8U_23U_o_expo_3_lpi_1_dfm_7_mx1w1!=8'b00000000);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_o_mant_3_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((or_11_cse & IsNaN_6U_10U_6_land_3_lpi_1_dfm_5) | and_1776_rgt)
        & (mux_1049_nl) ) begin
      FpAdd_8U_23U_o_mant_3_lpi_1_dfm_6 <= MUX_v_23_2_2(reg_chn_inp_in_crt_sva_3_574_544_1_reg,
          FpAdd_8U_23U_FpAdd_8U_23U_or_6_itm, and_4216_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_7 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_or_4_cse
        & (mux_1052_nl) ) begin
      inp_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_7 <= MUX_s_1_2_2(inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4,
          (inp_lookup_3_FpMul_6U_10U_1_p_mant_p1_mul_tmp[21]), and_dcpl_601);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_8U_23U_o_expo_lpi_1_dfm_11_reg <= 2'b0;
    end
    else if ( or_11_cse & core_wen & (chn_inp_in_crt_sva_3_739_736_1[3]) ) begin
      reg_FpAdd_8U_23U_o_expo_lpi_1_dfm_11_reg <= FpAdd_8U_23U_o_expo_FpAdd_8U_23U_o_expo_mux_3_rgt[7:6];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_4_cse & (~
        (mux_1056_nl)) ) begin
      FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5 <= MUX_s_1_2_2(FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_1_mx0w0,
          (FpMul_6U_10U_1_else_2_else_and_3_nl), and_dcpl_631);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2 <= 1'b0;
      inp_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_6 <= 1'b0;
    end
    else if ( IsZero_8U_23U_3_and_3_cse ) begin
      inp_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_3_or_itm_2 <= (FpAdd_8U_23U_o_mant_lpi_1_dfm_2_mx2!=23'b00000000000000000000000)
          | (FpAdd_8U_23U_o_expo_lpi_1_dfm_7_mx1w1!=8'b00000000);
      inp_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_6 <= inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_o_mant_lpi_1_dfm_6 <= 23'b0;
    end
    else if ( core_wen & ((or_11_cse & IsNaN_6U_10U_6_land_lpi_1_dfm_5) | and_1780_rgt)
        & (mux_1063_nl) ) begin
      FpAdd_8U_23U_o_mant_lpi_1_dfm_6 <= MUX_v_23_2_2(reg_chn_inp_in_crt_sva_3_606_576_1_reg,
          FpAdd_8U_23U_FpAdd_8U_23U_or_7_itm, and_4117_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_3_land_lpi_1_dfm_5 <= 1'b0;
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_16 <= 1'b0;
      chn_inp_in_crt_sva_5_459_1 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_3_aelse_and_4_cse ) begin
      IsNaN_8U_23U_3_land_lpi_1_dfm_5 <= MUX_s_1_2_2(IsNaN_8U_23U_3_land_lpi_1_dfm_mx0w0,
          FpAdd_6U_10U_1_is_a_greater_acc_3_itm_6_1, and_dcpl_679);
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_16 <= MUX_s_1_2_2(FpMul_6U_10U_1_lor_1_lpi_1_dfm_6,
          IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_3_tmp, and_dcpl_679);
      chn_inp_in_crt_sva_5_459_1 <= MUX_s_1_2_2(chn_inp_in_crt_sva_4_459_1, FpAdd_6U_10U_1_is_a_greater_acc_3_itm_6_1,
          and_dcpl_679);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_3_land_3_lpi_1_dfm_6 <= 1'b0;
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_17 <= 1'b0;
      chn_inp_in_crt_sva_5_443_1 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_3_aelse_and_5_cse ) begin
      IsNaN_8U_23U_3_land_3_lpi_1_dfm_6 <= MUX_s_1_2_2(FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_4,
          FpAdd_6U_10U_1_is_a_greater_acc_2_itm_6, and_dcpl_671);
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_17 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_16,
          IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_2_tmp, and_dcpl_671);
      chn_inp_in_crt_sva_5_443_1 <= MUX_s_1_2_2(chn_inp_in_crt_sva_4_443_1, FpAdd_6U_10U_1_is_a_greater_acc_2_itm_6,
          and_dcpl_671);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_3_land_2_lpi_1_dfm_6 <= 1'b0;
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_17 <= 1'b0;
      chn_inp_in_crt_sva_5_427_1 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_3_aelse_and_6_cse ) begin
      IsNaN_8U_23U_3_land_2_lpi_1_dfm_6 <= MUX_s_1_2_2(FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_4,
          FpAdd_6U_10U_1_is_a_greater_acc_1_itm_6, and_dcpl_663);
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_17 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_16,
          IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_1_tmp, and_dcpl_663);
      chn_inp_in_crt_sva_5_427_1 <= MUX_s_1_2_2(chn_inp_in_crt_sva_4_427_1, FpAdd_6U_10U_1_is_a_greater_acc_1_itm_6,
          and_dcpl_663);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_3_land_1_lpi_1_dfm_6 <= 1'b0;
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_17 <= 1'b0;
      chn_inp_in_crt_sva_5_411_1 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_3_aelse_and_7_cse ) begin
      IsNaN_8U_23U_3_land_1_lpi_1_dfm_6 <= MUX_s_1_2_2(FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_4,
          FpAdd_6U_10U_1_is_a_greater_acc_itm_6, and_dcpl_655);
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_17 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_16,
          IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_tmp, and_dcpl_655);
      chn_inp_in_crt_sva_5_411_1 <= MUX_s_1_2_2(chn_inp_in_crt_sva_4_411_1, FpAdd_6U_10U_1_is_a_greater_acc_itm_6,
          and_dcpl_655);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_5_30_0_itm <= 8'b0;
    end
    else if ( core_wen & (cfg_precision_1_sva_st_81==2'b10) & (chn_inp_in_crt_sva_4_739_736_1[0])
        & main_stage_v_4 & IsNaN_6U_10U_5_land_1_lpi_1_dfm_6 & or_11_cse ) begin
      reg_chn_inp_in_crt_sva_5_30_0_itm <= mux1h_47_itm[30:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_5_30_0_1_itm <= 23'b0;
    end
    else if ( ((FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_4 & (~ FpMul_6U_10U_1_lor_6_lpi_1_dfm_6))
        | IsNaN_6U_10U_5_land_1_lpi_1_dfm_6) & core_wen & (cfg_precision_1_sva_st_81==2'b10)
        & (chn_inp_in_crt_sva_4_739_736_1[0]) & main_stage_v_4 & or_11_cse ) begin
      reg_chn_inp_in_crt_sva_5_30_0_1_itm <= mux1h_47_itm[22:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_5_62_32_itm <= 8'b0;
    end
    else if ( core_wen & (cfg_precision_1_sva_st_81==2'b10) & (chn_inp_in_crt_sva_4_739_736_1[1])
        & main_stage_v_4 & IsNaN_6U_10U_5_land_2_lpi_1_dfm_6 & or_11_cse ) begin
      reg_chn_inp_in_crt_sva_5_62_32_itm <= mux1h_49_itm[30:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_5_62_32_1_itm <= 23'b0;
    end
    else if ( ((FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_4 & (~ FpMul_6U_10U_1_lor_7_lpi_1_dfm_6))
        | IsNaN_6U_10U_5_land_2_lpi_1_dfm_6) & core_wen & (cfg_precision_1_sva_st_81==2'b10)
        & (chn_inp_in_crt_sva_4_739_736_1[1]) & main_stage_v_4 & or_11_cse ) begin
      reg_chn_inp_in_crt_sva_5_62_32_1_itm <= mux1h_49_itm[22:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_5_94_64_itm <= 8'b0;
    end
    else if ( core_wen & (cfg_precision_1_sva_st_81==2'b10) & (chn_inp_in_crt_sva_4_739_736_1[2])
        & main_stage_v_4 & IsNaN_6U_10U_5_land_3_lpi_1_dfm_6 & or_11_cse ) begin
      reg_chn_inp_in_crt_sva_5_94_64_itm <= mux1h_51_itm[30:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_5_94_64_1_itm <= 23'b0;
    end
    else if ( ((FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_4 & (~ FpMul_6U_10U_1_lor_8_lpi_1_dfm_6))
        | IsNaN_6U_10U_5_land_3_lpi_1_dfm_6) & core_wen & (cfg_precision_1_sva_st_81==2'b10)
        & (chn_inp_in_crt_sva_4_739_736_1[2]) & main_stage_v_4 & or_11_cse ) begin
      reg_chn_inp_in_crt_sva_5_94_64_1_itm <= mux1h_51_itm[22:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_5_126_96_itm <= 8'b0;
    end
    else if ( core_wen & (cfg_precision_1_sva_st_81==2'b10) & (chn_inp_in_crt_sva_4_739_736_1[3])
        & main_stage_v_4 & FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_4 & or_11_cse ) begin
      reg_chn_inp_in_crt_sva_5_126_96_itm <= mux1h_53_itm[30:23];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_inp_in_crt_sva_5_126_96_1_itm <= 23'b0;
    end
    else if ( ((~(IsNaN_8U_23U_2_land_lpi_1_dfm_st_7 | IsNaN_6U_10U_5_land_lpi_1_dfm_6
        | IsNaN_6U_10U_4_land_lpi_1_dfm_5)) | FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_4)
        & core_wen & (cfg_precision_1_sva_st_81==2'b10) & (chn_inp_in_crt_sva_4_739_736_1[3])
        & main_stage_v_4 & or_11_cse ) begin
      reg_chn_inp_in_crt_sva_5_126_96_1_itm <= mux1h_53_itm[22:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_2_land_1_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_654 | and_1794_rgt | and_1796_rgt) & (~ mux_1066_itm)
        ) begin
      IsNaN_8U_23U_2_land_1_lpi_1_dfm_9 <= MUX1HOT_s_1_3_2(IsNaN_6U_10U_5_land_1_lpi_1_dfm_6,
          inp_lookup_1_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp, inp_lookup_1_FpAdd_6U_10U_1_is_a_greater_oif_equal_svs,
          {and_dcpl_654 , and_1794_rgt , and_1796_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
          <= 1'b0;
      inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6
          <= 1'b0;
    end
    else if ( FpAdd_6U_10U_1_is_addition_and_cse ) begin
      inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
          <= chn_inp_in_crt_sva_4_411_1;
      inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6
          <= inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_2_land_2_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_662 | and_1798_rgt | and_1800_rgt) & (~ mux_1067_itm)
        ) begin
      IsNaN_8U_23U_2_land_2_lpi_1_dfm_9 <= MUX1HOT_s_1_3_2(IsNaN_6U_10U_5_land_2_lpi_1_dfm_6,
          inp_lookup_2_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp, inp_lookup_2_FpAdd_6U_10U_1_is_a_greater_oif_equal_svs,
          {and_dcpl_662 , and_1798_rgt , and_1800_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
          <= 1'b0;
      inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6
          <= 1'b0;
    end
    else if ( FpAdd_6U_10U_1_is_addition_and_1_cse ) begin
      inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
          <= chn_inp_in_crt_sva_4_427_1;
      inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6
          <= inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_2_land_3_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_670 | and_1802_rgt | and_1804_rgt) & (~ mux_1067_itm)
        ) begin
      IsNaN_8U_23U_2_land_3_lpi_1_dfm_9 <= MUX1HOT_s_1_3_2(IsNaN_6U_10U_5_land_3_lpi_1_dfm_6,
          inp_lookup_3_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp, inp_lookup_3_FpAdd_6U_10U_1_is_a_greater_oif_equal_svs,
          {and_dcpl_670 , and_1802_rgt , and_1804_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
          <= 1'b0;
      inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6
          <= 1'b0;
    end
    else if ( FpAdd_6U_10U_1_is_addition_and_2_cse ) begin
      inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
          <= chn_inp_in_crt_sva_4_443_1;
      inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6
          <= inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_2_land_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_678 | and_1806_rgt | and_1808_rgt) & (~ mux_1066_itm)
        ) begin
      IsNaN_8U_23U_2_land_lpi_1_dfm_9 <= MUX1HOT_s_1_3_2(FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_4,
          inp_lookup_4_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp, inp_lookup_4_FpAdd_6U_10U_1_is_a_greater_oif_equal_svs,
          {and_dcpl_678 , and_1806_rgt , and_1808_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
          <= 1'b0;
      inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5
          <= 1'b0;
    end
    else if ( FpAdd_6U_10U_1_is_addition_and_3_cse ) begin
      inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
          <= IsNaN_8U_23U_2_land_lpi_1_dfm_st_7;
      inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5
          <= chn_inp_in_crt_sva_4_459_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_6_5_1 <= 1'b0;
    end
    else if ( core_wen & FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_3_cse & not_tmp_1029
        ) begin
      FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_6_5_1 <= MUX_s_1_2_2(FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_3_5_mx1w1,
          inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5,
          and_dcpl_654);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_6_3_0_1 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1091_nl) ) begin
      FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_6_3_0_1 <= FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_3_3_0_mx1w1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_7_5_1 <= 1'b0;
      FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_7_4_1 <= 1'b0;
      FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_7_3_0_1 <= 4'b0;
    end
    else if ( FpMul_6U_10U_2_o_expo_and_12_cse ) begin
      FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_7_5_1 <= FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_5_1;
      FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_7_4_1 <= FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_4_1;
      FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_7_3_0_1 <= FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_3_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_itm_3 <= 1'b0;
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_itm_10 <= 1'b0;
    end
    else if ( IsZero_6U_10U_9_and_cse ) begin
      inp_lookup_1_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_itm_3 <= MUX_s_1_2_2(IsZero_6U_10U_1_IsZero_6U_10U_1_and_itm_9,
          inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5,
          and_dcpl_654);
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_itm_10 <= MUX_s_1_2_2(IsZero_6U_10U_1_IsZero_6U_10U_1_and_itm_9,
          (inp_lookup_1_FpAdd_6U_10U_1_IsZero_6U_10U_8_or_nl), and_dcpl_655);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_6_5_1 <= 1'b0;
    end
    else if ( core_wen & FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_2_cse & not_tmp_1046
        ) begin
      FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_6_5_1 <= MUX_s_1_2_2(FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_3_5_mx1w1,
          inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5,
          and_dcpl_662);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_6_3_0_1 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1108_nl) ) begin
      FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_6_3_0_1 <= FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_3_3_0_mx1w1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_7_5_1 <= 1'b0;
      FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_7_4_1 <= 1'b0;
      FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_7_3_0_1 <= 4'b0;
    end
    else if ( FpMul_6U_10U_2_o_expo_and_15_cse ) begin
      FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_7_5_1 <= FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_5_1;
      FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_7_4_1 <= FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_4_1;
      FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_7_3_0_1 <= FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_3_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_itm_3 <= 1'b0;
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_1_itm_8 <= 1'b0;
    end
    else if ( IsZero_6U_10U_9_and_1_cse ) begin
      inp_lookup_2_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_itm_3 <= MUX_s_1_2_2(IsZero_6U_10U_1_IsZero_6U_10U_1_and_1_itm_7,
          inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5,
          and_dcpl_662);
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_1_itm_8 <= MUX_s_1_2_2(IsZero_6U_10U_1_IsZero_6U_10U_1_and_1_itm_7,
          (inp_lookup_2_FpAdd_6U_10U_1_IsZero_6U_10U_8_or_nl), and_dcpl_663);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_6_5_1 <= 1'b0;
    end
    else if ( core_wen & FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_1_cse & not_tmp_1063
        ) begin
      FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_6_5_1 <= MUX_s_1_2_2(FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_5_mx1w1,
          inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5,
          and_dcpl_670);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_6_3_0_1 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1125_nl) ) begin
      FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_6_3_0_1 <= FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_3_0_mx1w1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_7_5_1 <= 1'b0;
      FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_7_4_1 <= 1'b0;
      FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_7_3_0_1 <= 4'b0;
    end
    else if ( FpMul_6U_10U_2_o_expo_and_18_cse ) begin
      FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_7_5_1 <= FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_5_1;
      FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_7_4_1 <= FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_4_1;
      FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_7_3_0_1 <= FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_3_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_itm_3 <= 1'b0;
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_itm_10 <= 1'b0;
    end
    else if ( IsZero_6U_10U_9_and_2_cse ) begin
      inp_lookup_3_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_itm_3 <= MUX_s_1_2_2(IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_itm_9,
          inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5,
          and_dcpl_670);
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_itm_10 <= MUX_s_1_2_2(IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_itm_9,
          (inp_lookup_3_FpAdd_6U_10U_1_IsZero_6U_10U_8_or_nl), and_dcpl_671);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_lpi_1_dfm_6_5_1 <= 1'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_2_aelse_IsNaN_8U_23U_2_aelse_or_cse & not_tmp_1080
        ) begin
      FpMul_6U_10U_1_o_expo_lpi_1_dfm_6_5_1 <= MUX_s_1_2_2(FpMul_6U_10U_1_o_expo_lpi_1_dfm_3_5_mx0w1,
          inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4,
          and_dcpl_678);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_lpi_1_dfm_6_3_0_1 <= 4'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1143_nl) ) begin
      FpMul_6U_10U_1_o_expo_lpi_1_dfm_6_3_0_1 <= FpMul_6U_10U_1_o_expo_lpi_1_dfm_3_3_0_mx0w1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_o_expo_lpi_1_dfm_7_5_1 <= 1'b0;
      FpMul_6U_10U_2_o_expo_lpi_1_dfm_7_4_1 <= 1'b0;
      FpMul_6U_10U_2_o_expo_lpi_1_dfm_7_3_0_1 <= 4'b0;
    end
    else if ( FpMul_6U_10U_2_o_expo_and_21_cse ) begin
      FpMul_6U_10U_2_o_expo_lpi_1_dfm_7_5_1 <= FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_5_1;
      FpMul_6U_10U_2_o_expo_lpi_1_dfm_7_4_1 <= FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_4_1;
      FpMul_6U_10U_2_o_expo_lpi_1_dfm_7_3_0_1 <= FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_3_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_itm_3 <= 1'b0;
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_3_itm_8 <= 1'b0;
    end
    else if ( IsZero_6U_10U_9_and_3_cse ) begin
      inp_lookup_4_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_itm_3 <= MUX_s_1_2_2(IsZero_6U_10U_1_IsZero_6U_10U_1_and_3_itm_7,
          inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_11, and_dcpl_678);
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_3_itm_8 <= MUX_s_1_2_2(IsZero_6U_10U_1_IsZero_6U_10U_1_and_3_itm_7,
          (inp_lookup_4_FpAdd_6U_10U_1_IsZero_6U_10U_8_or_nl), and_dcpl_679);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_2_lpi_1_dfm_3_5_1 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_1335 | and_dcpl_1338 | and_1816_rgt) & (mux_1156_nl)
        ) begin
      FpAdd_6U_10U_1_qr_2_lpi_1_dfm_3_5_1 <= MUX1HOT_s_1_3_2(FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_6_5_1,
          FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_7_5_1, FpMantRNE_49U_24U_1_else_carry_1_sva_mx0w2,
          {and_dcpl_1335 , and_dcpl_1338 , and_1816_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_2_lpi_1_dfm_3_4_1 <= 1'b0;
    end
    else if ( core_wen & (((FpAdd_6U_10U_1_is_a_greater_oelse_FpAdd_6U_10U_1_is_a_greater_oelse_and_cse
        | IsNaN_8U_23U_3_land_1_lpi_1_dfm_6 | (chn_inp_in_crt_sva_5_739_736_1[0]))
        & or_11_cse) | and_dcpl_1338) & (~ mux_516_itm) ) begin
      FpAdd_6U_10U_1_qr_2_lpi_1_dfm_3_4_1 <= MUX_s_1_2_2(FpAdd_8U_23U_1_o_sign_1_lpi_1_dfm_5,
          FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_7_4_1, and_dcpl_1338);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_2_lpi_1_dfm_3_3_0_1 <= 4'b0;
    end
    else if ( core_wen & (and_dcpl_1335 | and_1821_rgt) & (~ (mux_1157_nl)) ) begin
      FpAdd_6U_10U_1_qr_2_lpi_1_dfm_3_3_0_1 <= MUX_v_4_2_2(FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_6_3_0_1,
          FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_7_3_0_1, and_1821_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_3_lpi_1_dfm_3_5_1 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_1348 | and_dcpl_1351 | and_1829_rgt) & (mux_1160_nl)
        ) begin
      FpAdd_6U_10U_1_qr_3_lpi_1_dfm_3_5_1 <= MUX1HOT_s_1_3_2(FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_6_5_1,
          FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_7_5_1, FpMantRNE_49U_24U_1_else_carry_2_sva_mx0w2,
          {and_dcpl_1348 , and_dcpl_1351 , and_1829_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_3_lpi_1_dfm_3_4_1 <= 1'b0;
    end
    else if ( core_wen & (((FpAdd_6U_10U_1_is_a_greater_oelse_FpAdd_6U_10U_1_is_a_greater_oelse_and_1_cse
        | IsNaN_8U_23U_3_land_2_lpi_1_dfm_6 | (chn_inp_in_crt_sva_5_739_736_1[1]))
        & or_11_cse) | and_dcpl_1351) & (~ mux_530_itm) ) begin
      FpAdd_6U_10U_1_qr_3_lpi_1_dfm_3_4_1 <= MUX_s_1_2_2(FpAdd_8U_23U_1_o_sign_2_lpi_1_dfm_5,
          FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_7_4_1, and_dcpl_1351);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_3_lpi_1_dfm_3_3_0_1 <= 4'b0;
    end
    else if ( core_wen & (and_dcpl_1348 | and_1834_rgt) & (~ (mux_1161_nl)) ) begin
      FpAdd_6U_10U_1_qr_3_lpi_1_dfm_3_3_0_1 <= MUX_v_4_2_2(FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_6_3_0_1,
          FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_7_3_0_1, and_1834_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_4_lpi_1_dfm_3_5_1 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_1361 | and_dcpl_1364 | and_1842_rgt) & (mux_1164_nl)
        ) begin
      FpAdd_6U_10U_1_qr_4_lpi_1_dfm_3_5_1 <= MUX1HOT_s_1_3_2(FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_6_5_1,
          FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_7_5_1, FpMantRNE_49U_24U_1_else_carry_3_sva_mx0w2,
          {and_dcpl_1361 , and_dcpl_1364 , and_1842_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_4_lpi_1_dfm_3_4_1 <= 1'b0;
    end
    else if ( core_wen & (((FpAdd_6U_10U_1_is_a_greater_oelse_FpAdd_6U_10U_1_is_a_greater_oelse_and_2_cse
        | IsNaN_8U_23U_3_land_3_lpi_1_dfm_6 | (chn_inp_in_crt_sva_5_739_736_1[2]))
        & or_11_cse) | and_dcpl_1364) & (~ mux_540_itm) ) begin
      FpAdd_6U_10U_1_qr_4_lpi_1_dfm_3_4_1 <= MUX_s_1_2_2(FpAdd_8U_23U_1_o_sign_3_lpi_1_dfm_5,
          FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_7_4_1, and_dcpl_1364);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_4_lpi_1_dfm_3_3_0_1 <= 4'b0;
    end
    else if ( core_wen & (and_dcpl_1361 | and_1847_rgt) & (~ (mux_1165_nl)) ) begin
      FpAdd_6U_10U_1_qr_4_lpi_1_dfm_3_3_0_1 <= MUX_v_4_2_2(FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_6_3_0_1,
          FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_7_3_0_1, and_1847_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_lpi_1_dfm_3_5_1 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_1374 | and_dcpl_1377 | and_1855_rgt) & (mux_1168_nl)
        ) begin
      FpAdd_6U_10U_1_qr_lpi_1_dfm_3_5_1 <= MUX1HOT_s_1_3_2(FpMul_6U_10U_1_o_expo_lpi_1_dfm_6_5_1,
          FpMul_6U_10U_2_o_expo_lpi_1_dfm_7_5_1, FpMantRNE_49U_24U_1_else_carry_sva_mx0w2,
          {and_dcpl_1374 , and_dcpl_1377 , and_1855_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_lpi_1_dfm_3_4_1 <= 1'b0;
    end
    else if ( core_wen & (((and_dcpl_1373 | IsNaN_8U_23U_3_land_lpi_1_dfm_5 | (chn_inp_in_crt_sva_5_739_736_1[3]))
        & or_11_cse) | and_dcpl_1377) & (~ mux_516_itm) ) begin
      FpAdd_6U_10U_1_qr_lpi_1_dfm_3_4_1 <= MUX_s_1_2_2(FpAdd_8U_23U_1_o_sign_lpi_1_dfm_5,
          FpMul_6U_10U_2_o_expo_lpi_1_dfm_7_4_1, and_dcpl_1377);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_1_qr_lpi_1_dfm_3_3_0_1 <= 4'b0;
    end
    else if ( core_wen & (and_dcpl_1374 | and_1860_rgt) & (~ (mux_1169_nl)) ) begin
      FpAdd_6U_10U_1_qr_lpi_1_dfm_3_3_0_1 <= MUX_v_4_2_2(FpMul_6U_10U_1_o_expo_lpi_1_dfm_6_3_0_1,
          FpMul_6U_10U_2_o_expo_lpi_1_dfm_7_3_0_1, and_1860_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_mant_lpi_1_dfm_10 <= 10'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ mux_1172_itm) ) begin
      FpMul_6U_10U_1_o_mant_lpi_1_dfm_10 <= FpMul_6U_10U_1_o_mant_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_8_itm_4_3 <= 2'b0;
      reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_8_itm_2_0 <= 3'b0;
      reg_FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_8_3_0_itm <= 1'b0;
    end
    else if ( and_3875_ssc ) begin
      reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_8_itm_4_3 <= reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_7_itm;
      reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_8_itm_2_0 <= reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_7_1_itm[7:5];
      reg_FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_8_3_0_itm <= FpMul_6U_10U_1_o_expo_mux1h_35_itm[3];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_8_1_itm <= 5'b0;
      reg_FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_8_3_0_1_itm <= 3'b0;
    end
    else if ( and_3880_cse ) begin
      reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_8_1_itm <= MUX_v_5_2_2((reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_7_1_itm[4:0]),
          (inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_nl), mux_tmp_1862);
      reg_FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_8_3_0_1_itm <= FpMul_6U_10U_1_o_expo_mux1h_35_itm[2:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_mant_2_lpi_1_dfm_11 <= 10'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ mux_1179_itm) ) begin
      FpMul_6U_10U_1_o_mant_2_lpi_1_dfm_11 <= FpMul_6U_10U_1_o_mant_2_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_mant_1_lpi_1_dfm_11 <= 10'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ mux_1182_itm) ) begin
      FpMul_6U_10U_1_o_mant_1_lpi_1_dfm_11 <= FpMul_6U_10U_1_o_mant_1_lpi_1_dfm_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_8_5_1 <= 1'b0;
    end
    else if ( core_wen & FpNormalize_6U_23U_1_if_FpNormalize_6U_23U_1_if_or_3_cse
        & (mux_1184_nl) ) begin
      FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_8_5_1 <= MUX_s_1_2_2(FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_7_5_1,
          FpMantRNE_24U_11U_else_carry_1_sva, and_dcpl_741);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_8_3_0_itm <= 1'b0;
    end
    else if ( core_wen & (cfg_precision_1_sva_st_83==2'b10) & or_tmp_2723 & main_stage_v_6
        & (~ (chn_inp_in_crt_sva_6_739_736_1[0])) & or_11_cse ) begin
      reg_FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_8_3_0_itm <= FpMul_6U_10U_1_o_expo_mux1h_23_itm[3];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_8_3_0_1_itm <= 3'b0;
    end
    else if ( (~ (mux_2120_nl)) & core_wen & (cfg_precision_1_sva_st_83==2'b10) &
        or_11_cse & main_stage_v_6 ) begin
      reg_FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_8_3_0_1_itm <= FpMul_6U_10U_1_o_expo_mux1h_23_itm[2:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_8_4_1 <= 1'b0;
    end
    else if ( core_wen & FpNormalize_6U_23U_1_if_FpNormalize_6U_23U_1_if_or_3_cse
        & (~ mux_1182_itm) ) begin
      FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_8_4_1 <= MUX_s_1_2_2(FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_7_4_1,
          FpAdd_6U_10U_1_qr_2_lpi_1_dfm_3_4_1, and_dcpl_741);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_8_5_1 <= 1'b0;
    end
    else if ( core_wen & FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_14_cse & (mux_1190_nl)
        ) begin
      FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_8_5_1 <= MUX_s_1_2_2(FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_7_5_1,
          FpMantRNE_24U_11U_else_carry_2_sva_mx0w1, and_dcpl_753);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_8_3_0_itm <= 1'b0;
    end
    else if ( core_wen & (cfg_precision_1_sva_st_83==2'b10) & or_tmp_2738 & main_stage_v_6
        & (~ (chn_inp_in_crt_sva_6_739_736_1[1])) & or_11_cse ) begin
      reg_FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_8_3_0_itm <= FpMul_6U_10U_1_o_expo_mux1h_29_itm[3];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_8_3_0_1_itm <= 3'b0;
    end
    else if ( (~ (mux_2122_nl)) & core_wen & (cfg_precision_1_sva_st_83==2'b10) &
        or_11_cse & main_stage_v_6 ) begin
      reg_FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_8_3_0_1_itm <= FpMul_6U_10U_1_o_expo_mux1h_29_itm[2:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_8_4_1 <= 1'b0;
    end
    else if ( core_wen & FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_14_cse & (~ mux_1179_itm)
        ) begin
      FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_8_4_1 <= MUX_s_1_2_2(FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_7_4_1,
          FpAdd_6U_10U_1_qr_3_lpi_1_dfm_3_4_1, and_dcpl_753);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_8_5_1 <= 1'b0;
    end
    else if ( core_wen & FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_13_cse & (mux_1196_nl)
        ) begin
      FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_8_5_1 <= MUX_s_1_2_2(FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_7_5_1,
          FpMantRNE_24U_11U_else_carry_3_sva_mx0w1, and_dcpl_765);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_8_4_1 <= 1'b0;
    end
    else if ( core_wen & FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_13_cse & (~ (mux_1198_nl))
        ) begin
      FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_8_4_1 <= MUX_s_1_2_2(FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_7_4_1,
          FpAdd_6U_10U_1_qr_4_lpi_1_dfm_3_4_1, and_dcpl_765);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_lpi_1_dfm_8_5_1 <= 1'b0;
    end
    else if ( core_wen & FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_12_cse & (mux_1201_nl)
        ) begin
      FpMul_6U_10U_1_o_expo_lpi_1_dfm_8_5_1 <= MUX_s_1_2_2(FpMul_6U_10U_1_o_expo_lpi_1_dfm_7_5_1,
          FpMantRNE_24U_11U_else_carry_sva_mx0w1, and_dcpl_777);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_6U_10U_1_o_expo_lpi_1_dfm_8_3_0_itm <= 1'b0;
    end
    else if ( core_wen & (cfg_precision_1_sva_st_83==2'b10) & or_tmp_2695 & main_stage_v_6
        & (~ (chn_inp_in_crt_sva_6_739_736_1[3])) & or_11_cse ) begin
      reg_FpMul_6U_10U_1_o_expo_lpi_1_dfm_8_3_0_itm <= FpMul_6U_10U_1_o_expo_mux1h_41_itm[3];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_6U_10U_1_o_expo_lpi_1_dfm_8_3_0_1_itm <= 3'b0;
    end
    else if ( (~ (mux_2126_nl)) & core_wen & (cfg_precision_1_sva_st_83==2'b10) &
        or_11_cse & main_stage_v_6 ) begin
      reg_FpMul_6U_10U_1_o_expo_lpi_1_dfm_8_3_0_1_itm <= FpMul_6U_10U_1_o_expo_mux1h_41_itm[2:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_lpi_1_dfm_8_4_1 <= 1'b0;
    end
    else if ( core_wen & FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_12_cse & (~ mux_1172_itm)
        ) begin
      FpMul_6U_10U_1_o_expo_lpi_1_dfm_8_4_1 <= MUX_s_1_2_2(FpMul_6U_10U_1_o_expo_lpi_1_dfm_7_4_1,
          FpAdd_6U_10U_1_qr_lpi_1_dfm_3_4_1, and_dcpl_777);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_20 <= 1'b0;
      IsNaN_6U_10U_land_1_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_2_aelse_and_12_cse ) begin
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_20 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_19,
          IsNaN_6U_10U_9_land_1_lpi_1_dfm_8, and_dcpl_785);
      IsNaN_6U_10U_land_1_lpi_1_dfm_5 <= MUX_s_1_2_2(IsNaN_6U_10U_IsNaN_6U_10U_nor_tmp,
          (IsNaN_6U_23U_2_IsNaN_6U_23U_2_nand_nl), and_dcpl_785);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_20 <= 1'b0;
      IsNaN_6U_10U_land_2_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_2_aelse_and_13_cse ) begin
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_20 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_19,
          IsNaN_6U_10U_9_land_2_lpi_1_dfm_8, and_dcpl_808);
      IsNaN_6U_10U_land_2_lpi_1_dfm_5 <= MUX_s_1_2_2(IsNaN_6U_10U_IsNaN_6U_10U_nor_1_tmp,
          (IsNaN_6U_23U_2_IsNaN_6U_23U_2_nand_1_nl), and_dcpl_808);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_20 <= 1'b0;
      IsNaN_6U_10U_land_3_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_2_aelse_and_14_cse ) begin
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_20 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_19,
          IsNaN_6U_10U_9_land_3_lpi_1_dfm_8, and_dcpl_832);
      IsNaN_6U_10U_land_3_lpi_1_dfm_5 <= MUX_s_1_2_2(IsNaN_6U_10U_IsNaN_6U_10U_nor_2_tmp,
          (IsNaN_6U_23U_2_IsNaN_6U_23U_2_nand_2_nl), and_dcpl_832);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_19 <= 1'b0;
      IsNaN_6U_10U_land_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_2_aelse_and_15_cse ) begin
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_19 <= MUX_s_1_2_2(IsNaN_6U_10U_2_land_lpi_1_dfm_st_18,
          IsNaN_6U_10U_9_land_lpi_1_dfm_8, and_dcpl_857);
      IsNaN_6U_10U_land_lpi_1_dfm_5 <= MUX_s_1_2_2(IsNaN_6U_10U_IsNaN_6U_10U_nor_3_tmp,
          (IsNaN_6U_23U_2_IsNaN_6U_23U_2_nand_3_nl), and_dcpl_857);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_1_lpi_1_dfm_9 <= 10'b0;
    end
    else if ( core_wen & ((or_11_cse & nor_1727_cse) | and_1871_rgt) & (~ mux_615_cse)
        ) begin
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_1_lpi_1_dfm_9 <= MUX_v_10_2_2((FpAdd_8U_23U_1_o_mant_1_lpi_1_dfm_6[9:0]),
          FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_mx0w1,
          and_1871_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_22 <= 10'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1208_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_22 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_21;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_2_lpi_1_dfm_9 <= 10'b0;
    end
    else if ( core_wen & ((or_11_cse & IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_5) | and_1873_rgt)
        & (~ (mux_1211_nl)) ) begin
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_2_lpi_1_dfm_9 <= MUX_v_10_2_2((FpAdd_8U_23U_1_o_mant_2_lpi_1_dfm_6[9:0]),
          FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_1_mx0w1,
          and_1873_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_22 <= 10'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1213_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_22 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_21;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_3_lpi_1_dfm_9 <= 10'b0;
    end
    else if ( core_wen & ((or_11_cse & IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_5) | and_1875_rgt)
        & (~ mux_635_cse) ) begin
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_3_lpi_1_dfm_9 <= MUX_v_10_2_2((FpAdd_8U_23U_1_o_mant_3_lpi_1_dfm_6[9:0]),
          FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_2_mx0w1,
          and_1875_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_lpi_1_dfm_9 <= 10'b0;
    end
    else if ( core_wen & ((or_11_cse & IsNaN_6U_10U_8_land_lpi_1_dfm_st_5) | and_1877_rgt)
        & (~ mux_645_cse) ) begin
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_lpi_1_dfm_9 <= MUX_v_10_2_2((FpAdd_8U_23U_1_o_mant_lpi_1_dfm_6[9:0]),
          FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_2_nor_3_mx0w1,
          and_1877_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_22 <= 10'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1219_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_22 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_21;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_23 <= 10'b0;
    end
    else if ( core_wen & ((or_11_cse & (~ IsNaN_6U_10U_land_1_lpi_1_dfm_5)) | and_dcpl_1404)
        & (mux_1220_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_23 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_22,
          FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_1_lpi_1_dfm_9, and_dcpl_1404);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_14_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_22 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_28_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_14_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_13_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_22 <= FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_3_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_11_4_0_1 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1222_nl)) ) begin
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_11_4_0_1 <= FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_10_4_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_14_0_1 <= 1'b0;
    end
    else if ( core_wen & (and_1881_rgt | and_dcpl_1404 | nor_1765_rgt | and_1888_rgt)
        & (~ mux_659_itm) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_14_0_1 <= MUX1HOT_s_1_4_2(FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_5_1,
          FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_10_5_1, inp_lookup_1_FpMul_6U_10U_else_2_if_acc_itm_6_1,
          inp_lookup_1_FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs,
          {and_1881_rgt , and_dcpl_1404 , nor_1765_rgt , and_1888_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_lor_6_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1223_nl) ) begin
      FpMul_6U_10U_lor_6_lpi_1_dfm_4 <= or_5020_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_23 <= 10'b0;
    end
    else if ( core_wen & ((or_11_cse & (~ IsNaN_6U_10U_land_2_lpi_1_dfm_5)) | and_dcpl_1415)
        & (mux_1224_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_23 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_22,
          FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_2_lpi_1_dfm_9, and_dcpl_1415);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_14_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_22 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_31_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_14_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_13_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_22 <= FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_3_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_11_4_0_1 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1226_nl)) ) begin
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_11_4_0_1 <= FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_10_4_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_14_0_1 <= 1'b0;
    end
    else if ( core_wen & (and_1892_rgt | and_dcpl_1415 | nor_1764_rgt | and_1899_rgt)
        & (~ mux_666_itm) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_14_0_1 <= MUX1HOT_s_1_4_2(FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_5_1,
          FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_10_5_1, inp_lookup_2_FpMul_6U_10U_else_2_if_acc_itm_6_1,
          inp_lookup_2_FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs,
          {and_1892_rgt , and_dcpl_1415 , nor_1764_rgt , and_1899_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_lor_7_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1227_nl) ) begin
      FpMul_6U_10U_lor_7_lpi_1_dfm_4 <= or_5021_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_22 <= 10'b0;
    end
    else if ( core_wen & ((or_11_cse & (~ IsNaN_6U_10U_land_3_lpi_1_dfm_5)) | and_dcpl_1426)
        & (mux_1228_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_22 <= MUX_v_10_2_2(FpAdd_6U_10U_1_FpAdd_6U_10U_1_or_2_itm_2,
          FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_3_lpi_1_dfm_9, and_dcpl_1426);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_14_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_22 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_34_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_14_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_13_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_22 <= FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_3_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_11_4_0_1 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1230_nl)) ) begin
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_11_4_0_1 <= FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_10_4_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_14_0_1 <= 1'b0;
    end
    else if ( core_wen & (and_1903_rgt | and_dcpl_1426 | nor_1763_rgt | and_1910_rgt)
        & (~ mux_673_itm) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_14_0_1 <= MUX1HOT_s_1_4_2(FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_5_1,
          FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_10_5_1, inp_lookup_3_FpMul_6U_10U_else_2_if_acc_itm_6_1,
          inp_lookup_3_FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs,
          {and_1903_rgt , and_dcpl_1426 , nor_1763_rgt , and_1910_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_lor_8_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1231_nl) ) begin
      FpMul_6U_10U_lor_8_lpi_1_dfm_4 <= or_5022_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_23 <= 10'b0;
    end
    else if ( core_wen & ((or_11_cse & (~ IsNaN_6U_10U_land_lpi_1_dfm_5)) | and_dcpl_1437)
        & (mux_1232_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_23 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_22,
          FpWidthDec_8U_23U_6U_10U_0U_1U_o_mant_lpi_1_dfm_9, and_dcpl_1437);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_14_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_22 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_37_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_14_1_1 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_13_1_1;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_22 <= FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_3_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_11_4_0_1 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1234_nl)) ) begin
      FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_11_4_0_1 <= FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_10_4_0_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_14_0_1 <= 1'b0;
    end
    else if ( core_wen & (and_1914_rgt | and_dcpl_1437 | nor_1762_rgt | and_1921_rgt)
        & (~ mux_680_itm) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_14_0_1 <= MUX1HOT_s_1_4_2(FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_5_1,
          FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_10_5_1, inp_lookup_4_FpMul_6U_10U_else_2_if_acc_itm_6_1,
          inp_lookup_4_FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs,
          {and_1914_rgt , and_dcpl_1437 , nor_1762_rgt , and_1921_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_lor_1_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1235_nl) ) begin
      FpMul_6U_10U_lor_1_lpi_1_dfm_4 <= or_5023_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_3_or_itm_2 <= 1'b0;
      inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_16 <= 1'b0;
    end
    else if ( IsZero_6U_10U_3_and_cse ) begin
      inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_3_or_itm_2 <= (FpMul_6U_10U_o_mant_1_lpi_1_dfm_3_mx0w0!=10'b0000000000)
          | FpMul_6U_10U_o_expo_1_lpi_1_dfm_3_5_mx0w0 | FpMul_6U_10U_o_expo_1_lpi_1_dfm_3_4_mx0w0
          | (FpMul_6U_10U_o_expo_1_lpi_1_dfm_3_3_0_mx0w0!=4'b0000);
      inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_16 <= inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_15;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_3_or_itm_2 <= 1'b0;
      inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_15 <= 1'b0;
    end
    else if ( IsZero_6U_10U_3_and_1_cse ) begin
      inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_3_or_itm_2 <= (FpMul_6U_10U_o_mant_2_lpi_1_dfm_3_mx0w0!=10'b0000000000)
          | FpMul_6U_10U_o_expo_2_lpi_1_dfm_3_5_mx0w0 | FpMul_6U_10U_o_expo_2_lpi_1_dfm_3_4_mx0w0
          | (FpMul_6U_10U_o_expo_2_lpi_1_dfm_3_3_0_mx0w0!=4'b0000);
      inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_15 <= inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_14;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_3_or_itm_2 <= 1'b0;
      inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_16 <= 1'b0;
    end
    else if ( IsZero_6U_10U_3_and_2_cse ) begin
      inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_3_or_itm_2 <= (FpMul_6U_10U_o_mant_3_lpi_1_dfm_3_mx0w0!=10'b0000000000)
          | FpMul_6U_10U_o_expo_3_lpi_1_dfm_3_5_mx0w0 | FpMul_6U_10U_o_expo_3_lpi_1_dfm_3_4_mx0w0
          | (FpMul_6U_10U_o_expo_3_lpi_1_dfm_3_3_0_mx0w0!=4'b0000);
      inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_16 <= inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_15;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_3_or_itm_2 <= 1'b0;
      inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_16 <= 1'b0;
    end
    else if ( IsZero_6U_10U_3_and_3_cse ) begin
      inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_3_or_itm_2 <= (FpMul_6U_10U_o_mant_lpi_1_dfm_3_mx0w0!=10'b0000000000)
          | FpMul_6U_10U_o_expo_lpi_1_dfm_3_5_mx0w0 | FpMul_6U_10U_o_expo_lpi_1_dfm_3_4_mx0w0
          | (FpMul_6U_10U_o_expo_lpi_1_dfm_3_3_0_mx0w0!=4'b0000);
      inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_16 <= inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_15;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_lpi_1_dfm_11 <= 10'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_7_4_1 <= 1'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_7_3_0_1 <= 4'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_lpi_1_dfm_11 <= 3'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_19_itm_7
          <= 1'b0;
    end
    else if ( FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_4_cse ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_lpi_1_dfm_11 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_lpi_1_dfm_10;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_7_4_1 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_6_4_1;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_7_3_0_1 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_6_3_0_1;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_lpi_1_dfm_11 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_lpi_1_dfm_10;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_19_itm_7
          <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_19_itm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_23U_3_land_lpi_1_dfm_9 <= 1'b0;
      IsNaN_6U_23U_3_land_3_lpi_1_dfm_9 <= 1'b0;
      IsNaN_6U_23U_3_land_2_lpi_1_dfm_9 <= 1'b0;
      IsNaN_6U_23U_3_land_1_lpi_1_dfm_9 <= 1'b0;
      inp_lookup_if_unequal_tmp_12 <= 1'b0;
      inp_lookup_else_unequal_tmp_37 <= 1'b0;
      chn_inp_in_crt_sva_11_739_736_1 <= 4'b0;
    end
    else if ( chn_inp_in_flow_and_40_cse ) begin
      IsNaN_6U_23U_3_land_lpi_1_dfm_9 <= IsNaN_6U_23U_3_land_lpi_1_dfm_8;
      IsNaN_6U_23U_3_land_3_lpi_1_dfm_9 <= IsNaN_6U_23U_3_land_3_lpi_1_dfm_8;
      IsNaN_6U_23U_3_land_2_lpi_1_dfm_9 <= IsNaN_6U_23U_3_land_2_lpi_1_dfm_8;
      IsNaN_6U_23U_3_land_1_lpi_1_dfm_9 <= IsNaN_6U_23U_3_land_1_lpi_1_dfm_8;
      inp_lookup_if_unequal_tmp_12 <= inp_lookup_if_unequal_tmp_1_mx0w0;
      inp_lookup_else_unequal_tmp_37 <= inp_lookup_else_unequal_tmp_36;
      chn_inp_in_crt_sva_11_739_736_1 <= chn_inp_in_crt_sva_10_739_736_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_25 <= 10'b0;
    end
    else if ( core_wen & FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_9_cse
        & (~ (mux_1246_nl)) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_25 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_24,
          FpMul_6U_10U_o_mant_lpi_1_dfm_7, and_dcpl_1448);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_28 <= 4'b0;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_16_tmp <= 1'b0;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_16_tmp_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_39_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_28 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_27,
          FpMul_6U_10U_o_expo_lpi_1_dfm_6_3_0_1, and_dcpl_1448);
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_16_tmp <= MUX_s_1_2_2(reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_15_tmp,
          reg_FpMul_6U_10U_o_expo_lpi_1_dfm_6_5_4_tmp, and_dcpl_1448);
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_16_tmp_1 <= MUX_s_1_2_2(reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_15_tmp_1,
          reg_FpMul_6U_10U_o_expo_lpi_1_dfm_6_5_4_tmp_1, and_dcpl_1448);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_3_lpi_1_dfm_11 <= 10'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_7_4_1 <= 1'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_7_3_0_1 <= 4'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_3_lpi_1_dfm_11 <= 3'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_14_itm_7
          <= 1'b0;
    end
    else if ( FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_5_cse ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_3_lpi_1_dfm_11 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_3_lpi_1_dfm_10;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_7_4_1 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_6_4_1;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_7_3_0_1 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_6_3_0_1;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_3_lpi_1_dfm_11 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_3_lpi_1_dfm_10;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_14_itm_7
          <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_14_itm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_28 <= 10'b0;
    end
    else if ( core_wen & FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_8_cse
        & (mux_1249_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_28 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_27,
          FpMul_6U_10U_o_mant_3_lpi_1_dfm_7, and_dcpl_1450);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_28 <= 4'b0;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_16_tmp <= 1'b0;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_16_tmp_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_41_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_28 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_27,
          FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_3_0_1, and_dcpl_1450);
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_16_tmp <= MUX_s_1_2_2(reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_15_tmp,
          reg_FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_5_4_tmp, and_dcpl_1450);
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_16_tmp_1 <= MUX_s_1_2_2(reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_15_tmp_1,
          reg_FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_5_4_tmp_1, and_dcpl_1450);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_2_lpi_1_dfm_11 <= 10'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_7_4_1 <= 1'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_7_3_0_1 <= 4'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_2_lpi_1_dfm_11 <= 3'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_9_itm_7
          <= 1'b0;
    end
    else if ( FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_6_cse ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_2_lpi_1_dfm_11 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_2_lpi_1_dfm_10;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_7_4_1 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_6_4_1;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_7_3_0_1 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_6_3_0_1;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_2_lpi_1_dfm_11 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_2_lpi_1_dfm_10;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_9_itm_7
          <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_9_itm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_25 <= 10'b0;
    end
    else if ( core_wen & FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_7_cse
        & (mux_1253_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_25 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_24,
          FpMul_6U_10U_o_mant_2_lpi_1_dfm_7, and_dcpl_1452);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_28 <= 4'b0;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_16_tmp <= 1'b0;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_16_tmp_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_43_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_28 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_27,
          FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_3_0_1, and_dcpl_1452);
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_16_tmp <= MUX_s_1_2_2(reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_15_tmp,
          reg_FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_5_4_tmp, and_dcpl_1452);
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_16_tmp_1 <= MUX_s_1_2_2(reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_15_tmp_1,
          reg_FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_5_4_tmp_1, and_dcpl_1452);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_1_lpi_1_dfm_11 <= 10'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_7_4_1 <= 1'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_7_3_0_1 <= 4'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_1_lpi_1_dfm_11 <= 3'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_4_itm_7
          <= 1'b0;
    end
    else if ( FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_7_cse ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_1_lpi_1_dfm_11 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_1_lpi_1_dfm_10;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_7_4_1 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_6_4_1;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_7_3_0_1 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_6_3_0_1;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_1_lpi_1_dfm_11 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_1_lpi_1_dfm_10;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_4_itm_7
          <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_4_itm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_25 <= 10'b0;
    end
    else if ( core_wen & FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_or_6_cse
        & (~ (mux_1259_nl)) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_25 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_24,
          FpMul_6U_10U_o_mant_1_lpi_1_dfm_7, and_dcpl_1454);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_28 <= 4'b0;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_16_tmp <= 1'b0;
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_16_tmp_1 <= 1'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_and_45_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_28 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_27,
          FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_3_0_1, and_dcpl_1454);
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_16_tmp <= MUX_s_1_2_2(reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_15_tmp,
          reg_FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_5_4_tmp, and_dcpl_1454);
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_16_tmp_1 <= MUX_s_1_2_2(reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_15_tmp_1,
          reg_FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_5_4_tmp_1, and_dcpl_1454);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_lpi_1_dfm_11_30_0_1 <= 31'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1263_nl) ) begin
      IntSaturation_51U_32U_o_lpi_1_dfm_11_30_0_1 <= IntSaturation_51U_32U_o_lpi_1_dfm_17[30:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_9_17_1_itm <= 8'b0;
    end
    else if ( or_11_cse & core_wen & main_stage_v_10 & (~ (chn_inp_in_crt_sva_10_739_736_1[3]))
        & inp_lookup_else_unequal_tmp_36 ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_9_17_1_itm <= reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_8_17_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_9_17_1_1_itm <= 9'b0;
    end
    else if ( and_dcpl_2461 & (~ (chn_inp_in_crt_sva_10_739_736_1[3])) & or_11_cse
        ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_9_17_1_1_itm <= reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_8_17_1_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_3_lpi_1_dfm_11_30_0_1 <= 31'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1267_nl) ) begin
      IntSaturation_51U_32U_o_3_lpi_1_dfm_11_30_0_1 <= IntSaturation_51U_32U_o_3_lpi_1_dfm_17[30:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_9_17_1_itm <= 8'b0;
    end
    else if ( or_11_cse & core_wen & main_stage_v_10 & (~ (chn_inp_in_crt_sva_10_739_736_1[2]))
        & inp_lookup_else_unequal_tmp_36 ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_9_17_1_itm <= reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_8_17_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_9_17_1_1_itm <= 9'b0;
    end
    else if ( and_dcpl_2461 & (~ (chn_inp_in_crt_sva_10_739_736_1[2])) & or_11_cse
        ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_9_17_1_1_itm <= reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_8_17_1_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_2_lpi_1_dfm_11_30_0_1 <= 31'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1271_nl) ) begin
      IntSaturation_51U_32U_o_2_lpi_1_dfm_11_30_0_1 <= IntSaturation_51U_32U_o_2_lpi_1_dfm_17[30:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_9_17_1_itm <= 8'b0;
    end
    else if ( or_11_cse & core_wen & main_stage_v_10 & (~ (chn_inp_in_crt_sva_10_739_736_1[1]))
        & inp_lookup_else_unequal_tmp_36 ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_9_17_1_itm <= reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_8_17_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_9_17_1_1_itm <= 9'b0;
    end
    else if ( and_dcpl_2461 & (~ (chn_inp_in_crt_sva_10_739_736_1[1])) & or_11_cse
        ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_9_17_1_1_itm <= reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_8_17_1_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_1_lpi_1_dfm_11_30_0_1 <= 31'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1275_nl) ) begin
      IntSaturation_51U_32U_o_1_lpi_1_dfm_11_30_0_1 <= IntSaturation_51U_32U_o_1_lpi_1_dfm_17[30:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_9_17_1_itm <= 8'b0;
    end
    else if ( or_11_cse & core_wen & main_stage_v_10 & (~ (chn_inp_in_crt_sva_10_739_736_1[0]))
        & inp_lookup_else_unequal_tmp_36 ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_9_17_1_itm <= reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_8_17_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_9_17_1_1_itm <= 9'b0;
    end
    else if ( and_dcpl_2461 & (~ (chn_inp_in_crt_sva_10_739_736_1[0])) & or_11_cse
        ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_9_17_1_1_itm <= reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_8_17_1_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_491_itm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1264_nl)) ) begin
      inp_lookup_else_mux_491_itm_7 <= inp_lookup_else_mux_491_itm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_368_itm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1268_nl)) ) begin
      inp_lookup_else_mux_368_itm_7 <= inp_lookup_else_mux_368_itm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_245_itm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1272_nl)) ) begin
      inp_lookup_else_mux_245_itm_7 <= inp_lookup_else_mux_245_itm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_122_itm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1276_nl)) ) begin
      inp_lookup_else_mux_122_itm_7 <= inp_lookup_else_mux_122_itm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_mux_1057_itm_3 <= 1'b0;
    end
    else if ( core_wen & (inp_lookup_if_or_6_rgt | inp_lookup_if_or_7_rgt | inp_lookup_if_and_31_rgt
        | and_1941_rgt) & mux_tmp_698 ) begin
      inp_lookup_mux_1057_itm_3 <= MUX1HOT_s_1_4_2(FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_19_itm_6,
          chn_inp_in_crt_sva_10_331_1, (IntSaturation_51U_32U_o_lpi_1_dfm_17[31]),
          inp_lookup_else_mux_485_itm_10, {inp_lookup_if_or_6_rgt , inp_lookup_if_or_7_rgt
          , inp_lookup_if_and_31_rgt , and_1941_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_mux_791_itm_3 <= 1'b0;
    end
    else if ( core_wen & (inp_lookup_if_or_4_rgt | inp_lookup_if_or_5_rgt | inp_lookup_if_and_23_rgt
        | and_1943_rgt) & mux_tmp_698 ) begin
      inp_lookup_mux_791_itm_3 <= MUX1HOT_s_1_4_2(FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_14_itm_6,
          chn_inp_in_crt_sva_10_315_1, (IntSaturation_51U_32U_o_3_lpi_1_dfm_17[31]),
          inp_lookup_else_mux_362_itm_10, {inp_lookup_if_or_4_rgt , inp_lookup_if_or_5_rgt
          , inp_lookup_if_and_23_rgt , and_1943_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_mux_525_itm_3 <= 1'b0;
    end
    else if ( core_wen & (inp_lookup_if_or_2_rgt | inp_lookup_if_or_3_rgt | inp_lookup_if_and_15_rgt
        | and_1945_rgt) & mux_tmp_698 ) begin
      inp_lookup_mux_525_itm_3 <= MUX1HOT_s_1_4_2(FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_9_itm_6,
          chn_inp_in_crt_sva_10_299_1, (IntSaturation_51U_32U_o_2_lpi_1_dfm_17[31]),
          inp_lookup_else_mux_239_itm_10, {inp_lookup_if_or_2_rgt , inp_lookup_if_or_3_rgt
          , inp_lookup_if_and_15_rgt , and_1945_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_mux_259_itm_3 <= 1'b0;
    end
    else if ( core_wen & (inp_lookup_if_or_rgt | inp_lookup_if_or_1_rgt | inp_lookup_if_and_7_rgt
        | and_1947_rgt) & mux_tmp_698 ) begin
      inp_lookup_mux_259_itm_3 <= MUX1HOT_s_1_4_2(FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_4_itm_6,
          chn_inp_in_crt_sva_10_283_1, (IntSaturation_51U_32U_o_1_lpi_1_dfm_17[31]),
          inp_lookup_else_mux_116_itm_10, {inp_lookup_if_or_rgt , inp_lookup_if_or_1_rgt
          , inp_lookup_if_and_7_rgt , and_1947_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_qr_2_lpi_1_dfm_3_0 <= 4'b0;
      reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_5_4_tmp <= 1'b0;
      reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_5_4_tmp_1 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_and_35_cse ) begin
      FpAdd_6U_10U_qr_2_lpi_1_dfm_3_0 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_27,
          FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_3_0_1, and_dcpl_1481);
      reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_5_4_tmp <= MUX_s_1_2_2(reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_15_tmp,
          reg_FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_5_4_tmp, and_dcpl_1481);
      reg_FpAdd_6U_10U_qr_2_lpi_1_dfm_5_4_tmp_1 <= MUX_s_1_2_2(reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_15_tmp_1,
          reg_FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_5_4_tmp_1, and_dcpl_1481);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_3_land_1_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1281_nl) ) begin
      IsNaN_6U_10U_3_land_1_lpi_1_dfm_6 <= IsNaN_6U_10U_3_IsNaN_6U_10U_3_nor_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_24 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1286_nl) ) begin
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_24 <= IsNaN_6U_10U_2_land_1_lpi_1_dfm_23;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_1_lpi_1_dfm_17 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1288_nl) ) begin
      IntSaturation_51U_32U_o_1_lpi_1_dfm_17 <= IntSaturation_51U_32U_o_1_lpi_1_dfm_16;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_qr_3_lpi_1_dfm_3_0 <= 4'b0;
      reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_5_4_tmp <= 1'b0;
      reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_5_4_tmp_1 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_and_37_cse ) begin
      FpAdd_6U_10U_qr_3_lpi_1_dfm_3_0 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_27,
          FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_3_0_1, and_dcpl_1488);
      reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_5_4_tmp <= MUX_s_1_2_2(reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_15_tmp,
          reg_FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_5_4_tmp, and_dcpl_1488);
      reg_FpAdd_6U_10U_qr_3_lpi_1_dfm_5_4_tmp_1 <= MUX_s_1_2_2(reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_15_tmp_1,
          reg_FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_5_4_tmp_1, and_dcpl_1488);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_3_land_2_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1293_nl) ) begin
      IsNaN_6U_10U_3_land_2_lpi_1_dfm_6 <= IsNaN_6U_10U_3_IsNaN_6U_10U_3_nor_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_24 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1298_nl) ) begin
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_24 <= IsNaN_6U_10U_2_land_2_lpi_1_dfm_23;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_2_lpi_1_dfm_17 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1300_nl) ) begin
      IntSaturation_51U_32U_o_2_lpi_1_dfm_17 <= IntSaturation_51U_32U_o_2_lpi_1_dfm_16;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_qr_4_lpi_1_dfm_3_0 <= 4'b0;
      reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_5_4_tmp <= 1'b0;
      reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_5_4_tmp_1 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_and_39_cse ) begin
      FpAdd_6U_10U_qr_4_lpi_1_dfm_3_0 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_27,
          FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_3_0_1, and_dcpl_1497);
      reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_5_4_tmp <= MUX_s_1_2_2(reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_15_tmp,
          reg_FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_5_4_tmp, and_dcpl_1497);
      reg_FpAdd_6U_10U_qr_4_lpi_1_dfm_5_4_tmp_1 <= MUX_s_1_2_2(reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_15_tmp_1,
          reg_FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_5_4_tmp_1, and_dcpl_1497);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_3_land_3_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1305_nl) ) begin
      IsNaN_6U_10U_3_land_3_lpi_1_dfm_6 <= IsNaN_6U_10U_3_IsNaN_6U_10U_3_nor_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_24 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1310_nl) ) begin
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_24 <= IsNaN_6U_10U_2_land_3_lpi_1_dfm_23;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_3_lpi_1_dfm_17 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1312_nl) ) begin
      IntSaturation_51U_32U_o_3_lpi_1_dfm_17 <= IntSaturation_51U_32U_o_3_lpi_1_dfm_16;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_3_land_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1317_nl) ) begin
      IsNaN_6U_10U_3_land_lpi_1_dfm_6 <= IsNaN_6U_10U_3_IsNaN_6U_10U_3_nor_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_2_land_lpi_1_dfm_24 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1322_nl) ) begin
      IsNaN_6U_10U_2_land_lpi_1_dfm_24 <= IsNaN_6U_10U_2_land_lpi_1_dfm_23;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_lpi_1_dfm_17 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1324_nl) ) begin
      IntSaturation_51U_32U_o_lpi_1_dfm_17 <= IntSaturation_51U_32U_o_lpi_1_dfm_16;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_10_739_736_1 <= 4'b0;
      IsNaN_6U_23U_3_land_lpi_1_dfm_8 <= 1'b0;
      IsNaN_6U_23U_3_land_3_lpi_1_dfm_8 <= 1'b0;
      IsNaN_6U_23U_3_land_2_lpi_1_dfm_8 <= 1'b0;
      IsNaN_6U_23U_3_land_1_lpi_1_dfm_8 <= 1'b0;
      inp_lookup_else_unequal_tmp_36 <= 1'b0;
    end
    else if ( chn_inp_in_flow_and_36_cse ) begin
      chn_inp_in_crt_sva_10_739_736_1 <= chn_inp_in_crt_sva_9_739_736_1;
      IsNaN_6U_23U_3_land_lpi_1_dfm_8 <= IsNaN_6U_23U_3_land_lpi_1_dfm_7;
      IsNaN_6U_23U_3_land_3_lpi_1_dfm_8 <= IsNaN_6U_23U_3_land_3_lpi_1_dfm_7;
      IsNaN_6U_23U_3_land_2_lpi_1_dfm_8 <= IsNaN_6U_23U_3_land_2_lpi_1_dfm_7;
      IsNaN_6U_23U_3_land_1_lpi_1_dfm_8 <= IsNaN_6U_23U_3_land_1_lpi_1_dfm_7;
      inp_lookup_else_unequal_tmp_36 <= inp_lookup_else_unequal_tmp_35;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs <=
          1'b0;
    end
    else if ( core_wen & (~(inp_lookup_1_FpMul_6U_10U_oelse_1_acc_itm_7_1 | or_dcpl_294
        | (~ (cfg_precision_1_sva_st_85[1])) | (~ (chn_inp_in_crt_sva_8_739_736_1[0]))
        | reg_FpMul_6U_10U_lor_3_lpi_1_dfm_3_cse | and_dcpl_78)) ) begin
      inp_lookup_1_FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs <=
          inp_lookup_1_FpMul_6U_10U_else_2_if_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs <=
          1'b0;
    end
    else if ( core_wen & (~(inp_lookup_2_FpMul_6U_10U_oelse_1_acc_itm_7_1 | nand_544_cse
        | (~ (chn_inp_in_crt_sva_8_739_736_1[1])) | (cfg_precision_1_sva_st_85[0])
        | reg_FpMul_6U_10U_lor_4_lpi_1_dfm_3_cse | and_dcpl_78)) ) begin
      inp_lookup_2_FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs <=
          inp_lookup_2_FpMul_6U_10U_else_2_if_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs <=
          1'b0;
    end
    else if ( core_wen & (~(inp_lookup_3_FpMul_6U_10U_oelse_1_acc_itm_7_1 | or_dcpl_294
        | (~ (cfg_precision_1_sva_st_85[1])) | (~ (chn_inp_in_crt_sva_8_739_736_1[2]))
        | reg_FpMul_6U_10U_lor_5_lpi_1_dfm_3_cse | and_dcpl_78)) ) begin
      inp_lookup_3_FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs <=
          inp_lookup_3_FpMul_6U_10U_else_2_if_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs <=
          1'b0;
    end
    else if ( core_wen & (~(inp_lookup_4_FpMul_6U_10U_oelse_1_acc_itm_7_1 | or_dcpl_294
        | (~ (cfg_precision_1_sva_st_85[1])) | (~ (chn_inp_in_crt_sva_8_739_736_1[3]))
        | reg_FpMul_6U_10U_lor_lpi_1_dfm_3_cse | and_dcpl_78)) ) begin
      inp_lookup_4_FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs <=
          inp_lookup_4_FpMul_6U_10U_else_2_if_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_22U_11U_1_else_carry_2_sva_1 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_495 | and_1975_rgt | and_1978_rgt) & (~ (mux_882_nl))
        ) begin
      FpMantRNE_22U_11U_1_else_carry_2_sva_1 <= MUX1HOT_s_1_3_2(FpMantRNE_22U_11U_1_else_carry_2_sva,
          FpMantRNE_22U_11U_2_else_carry_2_sva_mx1w1, FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_7_1_1,
          {and_dcpl_495 , and_1975_rgt , and_1978_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_22U_11U_1_else_carry_sva <= 1'b0;
    end
    else if ( core_wen & ((~ or_tmp_4457) | and_dcpl_1007 | and_1982_rgt | and_1985_rgt)
        ) begin
      FpMantRNE_22U_11U_1_else_carry_sva <= MUX1HOT_s_1_3_2(FpMantRNE_22U_11U_1_else_carry_sva_mx0w1,
          FpMantRNE_22U_11U_2_else_carry_sva_mx0w2, FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_7_1_1,
          {and_dcpl_1007 , and_1982_rgt , and_1985_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_159 | and_dcpl_78 | or_457_cse)) ) begin
      inp_lookup_1_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs
          <= inp_lookup_1_FpMul_6U_10U_1_else_2_if_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_5_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~((and_dcpl_1247 & (inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_4_0_1[3:1]==3'b111)
        & inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_5_1 & and_dcpl_1243) | or_tmp_439
        | (chn_inp_in_crt_sva_2_739_736_1[0]) | or_dcpl_660)) ) begin
      IsNaN_6U_10U_5_land_1_lpi_1_dfm <= and_3246_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_163 | and_dcpl_78 | or_519_cse)) ) begin
      inp_lookup_2_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs
          <= inp_lookup_2_FpMul_6U_10U_1_else_2_if_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_5_land_2_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~((and_dcpl_1256 & (inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_6_4_0_1[3:2]==2'b11)
        & IsNaN_8U_23U_land_2_lpi_1_dfm_st_4 & (inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_6_4_0_1[4])
        & and_dcpl_1252) | or_tmp_439 | (chn_inp_in_crt_sva_2_739_736_1[1]) | or_dcpl_660))
        ) begin
      IsNaN_6U_10U_5_land_2_lpi_1_dfm <= and_3244_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_167 | and_dcpl_78 | or_593_cse)) ) begin
      inp_lookup_3_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs
          <= inp_lookup_3_FpMul_6U_10U_1_else_2_if_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_5_land_3_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~((and_dcpl_1265 & (inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_6_4_0_1[3:2]==2'b11)
        & IsNaN_8U_23U_land_3_lpi_1_dfm_st_4 & (inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_6_4_0_1[4])
        & and_dcpl_1261) | or_tmp_439 | (~ main_stage_v_2) | and_dcpl_78 | (chn_inp_in_crt_sva_2_739_736_1[2])))
        ) begin
      IsNaN_6U_10U_5_land_3_lpi_1_dfm <= and_3242_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_5809_cse | and_dcpl_78 | or_648_cse)) ) begin
      inp_lookup_4_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs
          <= inp_lookup_4_FpMul_6U_10U_1_else_2_if_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_5_land_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~((and_dcpl_1274 & (inp_lookup_else_if_a0_15_10_lpi_1_dfm_6_4_0_1[3:2]==2'b11)
        & IsNaN_8U_23U_land_lpi_1_dfm_st_4 & (inp_lookup_else_if_a0_15_10_lpi_1_dfm_6_4_0_1[4])
        & and_dcpl_1270) | (cfg_precision_1_sva_st_91!=2'b10) | (chn_inp_in_crt_sva_2_739_736_1[3])
        | or_dcpl_660)) ) begin
      IsNaN_6U_10U_5_land_lpi_1_dfm <= and_3240_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_8 <= 10'b0;
    end
    else if ( core_wen & ((and_dcpl_1534 & (chn_inp_in_rsci_d_mxwt[313]) & (chn_inp_in_rsci_d_mxwt[310])
        & (chn_inp_in_rsci_d_mxwt[314]) & IsDenorm_5U_10U_2_or_2_tmp & or_11_cse)
        | and_2012_rgt) & (~ mux_95_itm) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_8 <= MUX_v_10_2_2((chn_inp_in_rsci_d_mxwt[309:300]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_or_8_mx0w1,
          and_2012_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_8U_23U_1_nor_itm_2 <= 1'b0;
      IsNaN_8U_23U_1_IsNaN_8U_23U_1_nand_itm_2 <= 1'b0;
    end
    else if ( IsNaN_8U_23U_1_and_cse ) begin
      IsNaN_8U_23U_1_nor_itm_2 <= ~((chn_inp_in_rsci_d_mxwt[630:608]!=23'b00000000000000000000000));
      IsNaN_8U_23U_1_IsNaN_8U_23U_1_nand_itm_2 <= ~((chn_inp_in_rsci_d_mxwt[638:631]==8'b11111111));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_lor_6_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & FpFractionToFloat_35U_6U_10U_is_zero_FpFractionToFloat_35U_6U_10U_is_zero_or_3_cse
        & (mux_1327_nl) ) begin
      FpMul_6U_10U_2_lor_6_lpi_1_dfm_5 <= MUX_s_1_2_2(or_5873_cse, IsNaN_8U_23U_2_land_1_lpi_1_dfm_st_6,
          and_dcpl_394);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_7_land_1_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & (and_2013_rgt | and_2022_rgt | and_dcpl_394) & (~ mux_115_itm)
        ) begin
      IsNaN_6U_10U_7_land_1_lpi_1_dfm_5 <= MUX1HOT_s_1_3_2(and_3149_cse, IsNaN_6U_10U_7_land_1_lpi_1_dfm,
          nor_1869_cse, {and_2013_rgt , and_2022_rgt , and_dcpl_394});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_lor_7_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & FpFractionToFloat_35U_6U_10U_is_zero_FpFractionToFloat_35U_6U_10U_is_zero_or_2_cse
        & (mux_1329_nl) ) begin
      FpMul_6U_10U_2_lor_7_lpi_1_dfm_5 <= MUX_s_1_2_2(or_5890_cse, IsNaN_8U_23U_2_land_2_lpi_1_dfm_st_6,
          and_dcpl_402);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_7_land_2_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & (and_2023_rgt | and_2033_rgt | and_dcpl_402) & (~ mux_115_itm)
        ) begin
      IsNaN_6U_10U_7_land_2_lpi_1_dfm_5 <= MUX1HOT_s_1_3_2(and_4145_cse, IsNaN_6U_10U_7_land_2_lpi_1_dfm,
          IsNaN_8U_23U_1_land_2_lpi_1_dfm_4, {and_2023_rgt , and_2033_rgt , and_dcpl_402});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_lor_8_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & FpFractionToFloat_35U_6U_10U_is_zero_FpFractionToFloat_35U_6U_10U_is_zero_or_1_cse
        & (mux_1331_nl) ) begin
      FpMul_6U_10U_2_lor_8_lpi_1_dfm_5 <= MUX_s_1_2_2(FpMul_6U_10U_2_if_2_FpMul_6U_10U_2_if_2_or_5_tmp,
          IsNaN_8U_23U_2_land_3_lpi_1_dfm_st_6, and_dcpl_410);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_7_land_3_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & (and_2034_rgt | and_2043_rgt | and_dcpl_410) & (~ mux_115_itm)
        ) begin
      IsNaN_6U_10U_7_land_3_lpi_1_dfm_5 <= MUX1HOT_s_1_3_2(and_3249_cse, IsNaN_6U_10U_7_land_3_lpi_1_dfm,
          IsNaN_8U_23U_1_land_3_lpi_1_dfm_4, {and_2034_rgt , and_2043_rgt , and_dcpl_410});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_lor_1_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & FpFractionToFloat_35U_6U_10U_is_zero_FpFractionToFloat_35U_6U_10U_is_zero_or_cse
        & (mux_1333_nl) ) begin
      FpMul_6U_10U_2_lor_1_lpi_1_dfm_5 <= MUX_s_1_2_2(FpMul_6U_10U_2_if_2_FpMul_6U_10U_2_if_2_or_7_tmp,
          IsNaN_8U_23U_2_land_lpi_1_dfm_st_6, and_dcpl_416);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_7_land_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & (and_2044_rgt | and_2054_rgt | and_dcpl_416) & (~ mux_115_itm)
        ) begin
      IsNaN_6U_10U_7_land_lpi_1_dfm_5 <= MUX1HOT_s_1_3_2(and_3361_cse_1, IsNaN_6U_10U_7_land_lpi_1_dfm,
          IsNaN_8U_23U_1_land_lpi_1_dfm_4, {and_2044_rgt , and_2054_rgt , and_dcpl_416});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_8_reg <= 4'b0;
    end
    else if ( (mux_2001_nl) & or_11_cse & core_wen ) begin
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_8_reg <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_mux1h_11_rgt[9:6];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_8_1_reg <= 6'b0;
    end
    else if ( (~(or_5800_cse & ((cfg_precision_1_sva_st_80!=2'b10) | (chn_inp_in_crt_sva_3_739_736_1[0])
        | (~ main_stage_v_3)))) & or_11_cse & core_wen ) begin
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_8_1_reg <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_mux1h_11_rgt[5:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_10 <= 10'b0;
    end
    else if ( FpAdd_8U_23U_o_expo_and_cse & (and_2065_rgt | and_2067_rgt | and_dcpl_495
        | and_2069_rgt) & (mux_1342_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_10 <= MUX1HOT_v_10_4_2(({reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_7_itm
          , reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_7_1_itm}), FpFractionToFloat_35U_6U_10U_1_o_mant_2_lpi_1_dfm_8,
          FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_3_mx0w0, (FpMul_6U_10U_2_p_mant_20_1_2_lpi_1_dfm_3_mx0[19:10]),
          {and_2065_rgt , and_2067_rgt , and_dcpl_495 , and_2069_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_3_lpi_1_dfm_10 <= 10'b0;
    end
    else if ( core_wen & ((~((mux_1952_nl) | (fsm_output[0]))) | and_2073_rgt | and_2076_rgt
        | and_dcpl_530 | and_2078_rgt) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_3_lpi_1_dfm_10 <= MUX1HOT_v_10_4_2(FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_3_lpi_1_dfm_9,
          FpFractionToFloat_35U_6U_10U_1_o_mant_3_lpi_1_dfm_8, (FpMul_6U_10U_1_p_mant_20_1_3_lpi_1_dfm_3_mx0[19:10]),
          (FpMul_6U_10U_2_p_mant_20_1_3_lpi_1_dfm_3_mx0[19:10]), {and_2073_rgt ,
          and_2076_rgt , and_dcpl_530 , and_2078_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_8_reg <= 4'b0;
    end
    else if ( (mux_2002_nl) & or_11_cse & core_wen ) begin
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_8_reg <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_mux1h_16_rgt[9:6];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_8_1_reg <= 6'b0;
    end
    else if ( (mux_2003_nl) & or_11_cse & core_wen ) begin
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_8_1_reg <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_mux1h_16_rgt[5:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_lpi_1_dfm_7_5_1 <= 1'b0;
    end
    else if ( core_wen & FpMul_6U_10U_1_o_expo_FpMul_6U_10U_1_o_expo_or_7_cse & (mux_1345_nl)
        ) begin
      FpMul_6U_10U_1_o_expo_lpi_1_dfm_7_5_1 <= MUX1HOT_s_1_3_2(FpMul_6U_10U_1_o_expo_lpi_1_dfm_6_5_1,
          FpMul_6U_10U_2_o_expo_lpi_1_dfm_7_5_1, inp_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_1_itm_7_1,
          {and_dcpl_1617 , and_dcpl_1619 , and_dcpl_719});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_lpi_1_dfm_7_3_0_1 <= 4'b0;
    end
    else if ( core_wen & ((or_11_cse & IsNaN_6U_10U_8_land_lpi_1_dfm_4) | and_2097_rgt)
        & (mux_1346_nl) ) begin
      FpMul_6U_10U_1_o_expo_lpi_1_dfm_7_3_0_1 <= MUX_v_4_2_2(FpMul_6U_10U_1_o_expo_lpi_1_dfm_6_3_0_1,
          FpMul_6U_10U_2_o_expo_lpi_1_dfm_7_3_0_1, and_2097_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_lpi_1_dfm_7_4_1 <= 1'b0;
    end
    else if ( core_wen & FpMul_6U_10U_1_o_expo_FpMul_6U_10U_1_o_expo_or_7_cse & (~
        mux_1347_itm) ) begin
      FpMul_6U_10U_1_o_expo_lpi_1_dfm_7_4_1 <= MUX1HOT_s_1_3_2(FpAdd_8U_23U_1_o_sign_lpi_1_dfm_5,
          FpMul_6U_10U_2_o_expo_lpi_1_dfm_7_4_1, inp_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_1_itm_7_1,
          {and_dcpl_1617 , and_dcpl_1619 , and_dcpl_719});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_mant_lpi_1_dfm_9 <= 10'b0;
    end
    else if ( core_wen & ((or_5152_cse & or_11_cse) | and_dcpl_1619) & (~ mux_1347_itm)
        ) begin
      FpMul_6U_10U_1_o_mant_lpi_1_dfm_9 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_22,
          ({reg_FpMul_6U_10U_2_o_mant_lpi_1_dfm_7_reg , reg_FpMul_6U_10U_2_o_mant_lpi_1_dfm_7_1_reg}),
          and_dcpl_1619);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_7_5_1 <= 1'b0;
    end
    else if ( core_wen & FpMul_6U_10U_1_o_expo_FpMul_6U_10U_1_o_expo_or_5_cse & (~
        (mux_1350_nl)) ) begin
      FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_7_5_1 <= MUX1HOT_s_1_3_2(FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_6_5_1,
          FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_7_5_1, inp_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_1_itm_7,
          {and_dcpl_1624 , and_dcpl_1626 , and_dcpl_712});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_7_3_0_1 <= 4'b0;
    end
    else if ( core_wen & ((or_11_cse & IsNaN_6U_10U_8_land_3_lpi_1_dfm_4) | and_2104_rgt)
        & (~ (mux_1351_nl)) ) begin
      FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_7_3_0_1 <= MUX_v_4_2_2(FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_6_3_0_1,
          FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_7_3_0_1, and_2104_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_7_4_1 <= 1'b0;
    end
    else if ( core_wen & FpMul_6U_10U_1_o_expo_FpMul_6U_10U_1_o_expo_or_5_cse & (~
        (mux_1352_nl)) ) begin
      FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_7_4_1 <= MUX1HOT_s_1_3_2(FpAdd_8U_23U_1_o_sign_3_lpi_1_dfm_5,
          FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_7_4_1, inp_lookup_3_FpAdd_8U_23U_1_if_4_if_acc_1_itm_7,
          {and_dcpl_1624 , and_dcpl_1626 , and_dcpl_712});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_7_itm <= 2'b0;
    end
    else if ( and_dcpl_2487 & (~ (cfg_precision_1_sva_st_82[0])) & or_tmp_3153 &
        (cfg_precision_1_sva_st_82[1]) & (~ (chn_inp_in_crt_sva_5_739_736_1[2]))
        & or_11_cse ) begin
      reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_7_itm <= MUX_v_2_2_2(reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_6_itm,
          reg_FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_7_itm, and_dcpl_1626);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_7_1_itm <= 8'b0;
    end
    else if ( (mux_2129_nl) & and_dcpl_2487 & (~ (cfg_precision_1_sva_st_82[0]))
        & or_11_cse & (cfg_precision_1_sva_st_82[1]) ) begin
      reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_7_1_itm <= MUX1HOT_v_8_3_2(reg_FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_6_1_itm,
          reg_FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_7_1_itm, FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_2_mx0w0,
          {(FpMul_6U_10U_1_o_mant_or_nl) , and_dcpl_1626 , (FpMul_6U_10U_1_o_mant_and_8_nl)});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_7_5_1 <= 1'b0;
    end
    else if ( core_wen & FpMul_6U_10U_1_o_expo_FpMul_6U_10U_1_o_expo_or_3_cse & (mux_1359_nl)
        ) begin
      FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_7_5_1 <= MUX1HOT_s_1_3_2(FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_6_5_1,
          FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_7_5_1, inp_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_1_itm_7_1,
          {and_dcpl_1632 , and_dcpl_1634 , and_dcpl_701});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_7_3_0_1 <= 4'b0;
    end
    else if ( core_wen & ((or_11_cse & IsNaN_6U_10U_8_land_2_lpi_1_dfm_4) | and_2112_rgt)
        & (mux_1361_nl) ) begin
      FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_7_3_0_1 <= MUX_v_4_2_2(FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_6_3_0_1,
          FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_7_3_0_1, and_2112_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_7_4_1 <= 1'b0;
    end
    else if ( core_wen & FpMul_6U_10U_1_o_expo_FpMul_6U_10U_1_o_expo_or_3_cse & (~
        mux_1362_itm) ) begin
      FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_7_4_1 <= MUX1HOT_s_1_3_2(FpAdd_8U_23U_1_o_sign_2_lpi_1_dfm_5,
          FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_7_4_1, inp_lookup_2_FpAdd_8U_23U_1_if_4_if_acc_1_itm_7_1,
          {and_dcpl_1632 , and_dcpl_1634 , and_dcpl_701});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_mant_2_lpi_1_dfm_10 <= 10'b0;
    end
    else if ( core_wen & ((or_5154_cse & or_11_cse) | and_dcpl_1634) & (~ mux_1362_itm)
        ) begin
      FpMul_6U_10U_1_o_mant_2_lpi_1_dfm_10 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_22,
          ({reg_FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_7_itm , reg_FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_7_1_itm}),
          and_dcpl_1634);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_7_5_1 <= 1'b0;
    end
    else if ( core_wen & FpMul_6U_10U_1_o_expo_FpMul_6U_10U_1_o_expo_or_1_cse & (mux_1365_nl)
        ) begin
      FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_7_5_1 <= MUX1HOT_s_1_3_2(FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_6_5_1,
          FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_7_5_1, inp_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_1_itm_7_1,
          {and_dcpl_1639 , and_dcpl_1641 , and_dcpl_690});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_7_3_0_1 <= 4'b0;
    end
    else if ( core_wen & ((or_11_cse & IsNaN_6U_10U_8_land_1_lpi_1_dfm_6) | and_2119_rgt)
        & (mux_1366_nl) ) begin
      FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_7_3_0_1 <= MUX_v_4_2_2(FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_6_3_0_1,
          FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_7_3_0_1, and_2119_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_7_4_1 <= 1'b0;
    end
    else if ( core_wen & FpMul_6U_10U_1_o_expo_FpMul_6U_10U_1_o_expo_or_1_cse & (~
        mux_1367_itm) ) begin
      FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_7_4_1 <= MUX1HOT_s_1_3_2(FpAdd_8U_23U_1_o_sign_1_lpi_1_dfm_5,
          FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_7_4_1, inp_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_1_itm_7_1,
          {and_dcpl_1639 , and_dcpl_1641 , and_dcpl_690});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_mant_1_lpi_1_dfm_10 <= 10'b0;
    end
    else if ( core_wen & ((or_5155_cse & or_11_cse) | and_dcpl_1641) & (~ mux_1367_itm)
        ) begin
      FpMul_6U_10U_1_o_mant_1_lpi_1_dfm_10 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_22,
          ({reg_FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_7_itm , reg_FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_7_1_itm}),
          and_dcpl_1641);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_19 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ mux_586_itm) ) begin
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_19 <= IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_18;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_19 <= 1'b0;
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_18 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_2_aelse_and_30_cse ) begin
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_19 <= IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_18;
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_18 <= IsNaN_6U_10U_2_land_lpi_1_dfm_st_17;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_1_land_1_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_798 | and_dcpl_787 | and_dcpl_785) & (~ mux_623_itm)
        ) begin
      IsNaN_6U_10U_1_land_1_lpi_1_dfm_5 <= MUX1HOT_s_1_3_2(IsNaN_6U_10U_1_land_1_lpi_1_dfm_mx0w0,
          IsNaN_6U_10U_1_land_1_lpi_1_dfm, IsNaN_6U_10U_8_land_1_lpi_1_dfm_7, {and_dcpl_798
          , and_dcpl_787 , and_dcpl_785});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_1_land_2_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_821 | and_dcpl_810 | and_dcpl_808) & (~ mux_632_itm)
        ) begin
      IsNaN_6U_10U_1_land_2_lpi_1_dfm_5 <= MUX1HOT_s_1_3_2(IsNaN_6U_10U_1_land_2_lpi_1_dfm_mx0w0,
          IsNaN_6U_10U_1_land_2_lpi_1_dfm, IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_19,
          {and_dcpl_821 , and_dcpl_810 , and_dcpl_808});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_1_land_3_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_845 | and_dcpl_834 | and_dcpl_832) & (~ mux_623_itm)
        ) begin
      IsNaN_6U_10U_1_land_3_lpi_1_dfm_5 <= MUX1HOT_s_1_3_2(IsNaN_6U_10U_1_land_3_lpi_1_dfm_mx0w0,
          IsNaN_6U_10U_1_land_3_lpi_1_dfm, IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_19,
          {and_dcpl_845 , and_dcpl_834 , and_dcpl_832});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_1_land_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_870 | and_dcpl_859 | and_dcpl_857) & (~ mux_623_itm)
        ) begin
      IsNaN_6U_10U_1_land_lpi_1_dfm_5 <= MUX1HOT_s_1_3_2(IsNaN_6U_10U_1_land_lpi_1_dfm_mx0w0,
          IsNaN_6U_10U_1_land_lpi_1_dfm, IsNaN_6U_10U_2_land_lpi_1_dfm_st_18, {and_dcpl_870
          , and_dcpl_859 , and_dcpl_857});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_15 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1368_nl)) ) begin
      inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_15 <= inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_14;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_14 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1369_nl)) ) begin
      inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_14 <= inp_lookup_2_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_13;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_15 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1370_nl)) ) begin
      inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_15 <= inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_14;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_15 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1371_nl)) ) begin
      inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_15 <= inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_14;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_lpi_1_dfm_10 <= 10'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_6_4_1 <= 1'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_6_3_0_1 <= 4'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_lpi_1_dfm_10 <= 3'b0;
    end
    else if ( FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_8_cse ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_lpi_1_dfm_10 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_lpi_1_dfm_9;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_6_4_1 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_5_4_1;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_6_3_0_1 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_5_3_0_1;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_lpi_1_dfm_10 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_3_lpi_1_dfm_10 <= 10'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_6_4_1 <= 1'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_6_3_0_1 <= 4'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_3_lpi_1_dfm_10 <= 3'b0;
    end
    else if ( FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_9_cse ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_3_lpi_1_dfm_10 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_3_lpi_1_dfm_9;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_6_4_1 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_5_4_1;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_6_3_0_1 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_5_3_0_1;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_3_lpi_1_dfm_10 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_3_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_2_lpi_1_dfm_10 <= 10'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_6_4_1 <= 1'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_6_3_0_1 <= 4'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_2_lpi_1_dfm_10 <= 3'b0;
    end
    else if ( FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_10_cse ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_2_lpi_1_dfm_10 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_2_lpi_1_dfm_9;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_6_4_1 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_5_4_1;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_6_3_0_1 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_5_3_0_1;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_2_lpi_1_dfm_10 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_2_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_1_lpi_1_dfm_10 <= 10'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_6_4_1 <= 1'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_6_3_0_1 <= 4'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_1_lpi_1_dfm_10 <= 3'b0;
    end
    else if ( FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_11_cse ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_1_lpi_1_dfm_10 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_1_lpi_1_dfm_9;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_6_4_1 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_5_4_1;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_6_3_0_1 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_5_3_0_1;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_1_lpi_1_dfm_10 <= FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_1_lpi_1_dfm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_8_17_1_itm <= 8'b0;
    end
    else if ( or_11_cse & core_wen & main_stage_v_9 & (~ (chn_inp_in_crt_sva_9_739_736_1[3]))
        & inp_lookup_else_unequal_tmp_35 ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_8_17_1_itm <= reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_7_17_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_8_17_1_1_itm <= 9'b0;
    end
    else if ( and_dcpl_2500 & (~ (chn_inp_in_crt_sva_9_739_736_1[3])) & or_11_cse
        ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_8_17_1_1_itm <= reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_7_17_1_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_19_itm_6
          <= 1'b0;
    end
    else if ( core_wen & ((or_11_cse & (~ (chn_inp_in_crt_sva_9_739_736_1[3]))) |
        and_2125_rgt) & (mux_1384_nl) ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_19_itm_6
          <= MUX_s_1_2_2(FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_19_itm_5,
          FpMul_6U_10U_o_sign_lpi_1_dfm_5, and_2125_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_8_17_1_itm <= 8'b0;
    end
    else if ( or_11_cse & core_wen & main_stage_v_9 & (~ (chn_inp_in_crt_sva_9_739_736_1[2]))
        & inp_lookup_else_unequal_tmp_35 ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_8_17_1_itm <= reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_7_17_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_8_17_1_1_itm <= 9'b0;
    end
    else if ( and_dcpl_2500 & (~ (chn_inp_in_crt_sva_9_739_736_1[2])) & or_11_cse
        ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_8_17_1_1_itm <= reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_7_17_1_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_14_itm_6
          <= 1'b0;
    end
    else if ( core_wen & ((or_11_cse & (~ (chn_inp_in_crt_sva_9_739_736_1[2]))) |
        and_2130_rgt) & (mux_1393_nl) ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_14_itm_6
          <= MUX_s_1_2_2(FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_14_itm_5,
          FpMul_6U_10U_o_sign_3_lpi_1_dfm_5, and_2130_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_8_17_1_itm <= 8'b0;
    end
    else if ( or_11_cse & core_wen & main_stage_v_9 & (~ (chn_inp_in_crt_sva_9_739_736_1[1]))
        & inp_lookup_else_unequal_tmp_35 ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_8_17_1_itm <= reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_7_17_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_8_17_1_1_itm <= 9'b0;
    end
    else if ( and_dcpl_2500 & (~ (chn_inp_in_crt_sva_9_739_736_1[1])) & or_11_cse
        ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_8_17_1_1_itm <= reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_7_17_1_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_9_itm_6
          <= 1'b0;
    end
    else if ( core_wen & ((or_11_cse & (~ (chn_inp_in_crt_sva_9_739_736_1[1]))) |
        and_2135_rgt) & (mux_1402_nl) ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_9_itm_6
          <= MUX_s_1_2_2(FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_9_itm_5,
          FpMul_6U_10U_o_sign_2_lpi_1_dfm_5, and_2135_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_8_17_1_itm <= 8'b0;
    end
    else if ( or_11_cse & core_wen & main_stage_v_9 & (~ (chn_inp_in_crt_sva_9_739_736_1[0]))
        & inp_lookup_else_unequal_tmp_35 ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_8_17_1_itm <= reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_7_17_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_8_17_1_1_itm <= 9'b0;
    end
    else if ( and_dcpl_2500 & (~ (chn_inp_in_crt_sva_9_739_736_1[0])) & or_11_cse
        ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_8_17_1_1_itm <= reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_7_17_1_1_itm;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_4_itm_6
          <= 1'b0;
    end
    else if ( core_wen & ((or_11_cse & (~ (chn_inp_in_crt_sva_9_739_736_1[0]))) |
        and_2140_rgt) & (mux_1411_nl) ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_4_itm_6
          <= MUX_s_1_2_2(FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_4_itm_5,
          FpMul_6U_10U_o_sign_1_lpi_1_dfm_5, and_2140_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_491_itm_6 <= 1'b0;
      inp_lookup_else_mux_485_itm_10 <= 1'b0;
    end
    else if ( inp_lookup_else_and_20_cse ) begin
      inp_lookup_else_mux_491_itm_6 <= inp_lookup_else_mux_491_itm_5;
      inp_lookup_else_mux_485_itm_10 <= inp_lookup_else_mux_485_itm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_368_itm_6 <= 1'b0;
      inp_lookup_else_mux_362_itm_10 <= 1'b0;
    end
    else if ( inp_lookup_else_and_21_cse ) begin
      inp_lookup_else_mux_368_itm_6 <= inp_lookup_else_mux_368_itm_5;
      inp_lookup_else_mux_362_itm_10 <= inp_lookup_else_mux_362_itm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_245_itm_6 <= 1'b0;
      inp_lookup_else_mux_239_itm_10 <= 1'b0;
    end
    else if ( inp_lookup_else_and_22_cse ) begin
      inp_lookup_else_mux_245_itm_6 <= inp_lookup_else_mux_245_itm_5;
      inp_lookup_else_mux_239_itm_10 <= inp_lookup_else_mux_239_itm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_122_itm_6 <= 1'b0;
      inp_lookup_else_mux_116_itm_10 <= 1'b0;
    end
    else if ( inp_lookup_else_and_23_cse ) begin
      inp_lookup_else_mux_122_itm_6 <= inp_lookup_else_mux_122_itm_5;
      inp_lookup_else_mux_116_itm_10 <= inp_lookup_else_mux_116_itm_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_10_283_1 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1419_nl)) ) begin
      chn_inp_in_crt_sva_10_283_1 <= chn_inp_in_crt_sva_9_283_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_20 <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1420_nl) ) begin
      cfg_precision_1_sva_20 <= cfg_precision_1_sva_19;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_10_299_1 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1428_nl)) ) begin
      chn_inp_in_crt_sva_10_299_1 <= chn_inp_in_crt_sva_9_299_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_10_315_1 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1436_nl)) ) begin
      chn_inp_in_crt_sva_10_315_1 <= chn_inp_in_crt_sva_9_315_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_10_331_1 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1444_nl)) ) begin
      chn_inp_in_crt_sva_10_331_1 <= chn_inp_in_crt_sva_9_331_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_1_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~((~ main_stage_v_7) | (cfg_precision_1_sva_st_84!=2'b10)
        | IsNaN_6U_10U_IsNaN_6U_10U_nor_tmp | and_dcpl_78 | (~ (chn_inp_in_crt_sva_7_739_736_1[0]))))
        ) begin
      IsNaN_6U_10U_1_land_1_lpi_1_dfm <= IsNaN_6U_10U_1_land_1_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_1_land_2_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(nand_557_cse | (cfg_precision_1_sva_st_84[0]) | (~ (chn_inp_in_crt_sva_7_739_736_1[1]))
        | and_dcpl_78 | IsNaN_6U_10U_IsNaN_6U_10U_nor_1_tmp)) ) begin
      IsNaN_6U_10U_1_land_2_lpi_1_dfm <= IsNaN_6U_10U_1_land_2_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_1_land_3_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~((~ main_stage_v_7) | (cfg_precision_1_sva_st_84!=2'b10)
        | (~ (chn_inp_in_crt_sva_7_739_736_1[2])) | and_dcpl_78 | IsNaN_6U_10U_IsNaN_6U_10U_nor_2_tmp))
        ) begin
      IsNaN_6U_10U_1_land_3_lpi_1_dfm <= IsNaN_6U_10U_1_land_3_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_1_land_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_336 | (~ (cfg_precision_1_sva_st_84[1])) | (~
        (chn_inp_in_crt_sva_7_739_736_1[3])) | and_dcpl_78 | IsNaN_6U_10U_IsNaN_6U_10U_nor_3_tmp))
        ) begin
      IsNaN_6U_10U_1_land_lpi_1_dfm <= IsNaN_6U_10U_1_land_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_2010_cse | or_5873_cse | (chn_inp_in_crt_sva_1_739_395_1[341])
        | or_dcpl_8)) ) begin
      inp_lookup_1_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs
          <= inp_lookup_1_FpMul_6U_10U_2_else_2_if_acc_itm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_7_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~((and_dcpl_1545 & and_dcpl_1541 & (~ IsNaN_6U_10U_6_nor_tmp)
        & inp_lookup_1_FpMantRNE_36U_11U_1_else_and_svs_2 & (IntLeadZero_35U_1_leading_sign_35_0_rtn_1_sva_2[5])
        & FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_st_2) | or_dcpl_897 | or_dcpl_8))
        ) begin
      IsNaN_6U_10U_7_land_1_lpi_1_dfm <= and_3149_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_2010_cse | or_5890_cse | (chn_inp_in_crt_sva_1_739_395_1[342])
        | or_dcpl_8)) ) begin
      inp_lookup_2_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs
          <= inp_lookup_2_FpMul_6U_10U_2_else_2_if_acc_itm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_7_land_2_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~((and_dcpl_1556 & (FpFractionToFloat_35U_6U_10U_1_mux_40_tmp[4:3]==2'b11)
        & (~ IsNaN_6U_10U_6_nor_1_tmp) & (IntLeadZero_35U_1_leading_sign_35_0_rtn_2_sva_2[5])
        & FpFractionToFloat_35U_6U_10U_1_and_1_cse) | or_dcpl_903 | or_dcpl_8)) )
        begin
      IsNaN_6U_10U_7_land_2_lpi_1_dfm <= and_4145_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_2010_cse | FpMul_6U_10U_2_if_2_FpMul_6U_10U_2_if_2_or_5_tmp
        | (~ main_stage_v_1) | or_dcpl_906)) ) begin
      inp_lookup_3_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs
          <= inp_lookup_3_FpMul_6U_10U_2_else_2_if_acc_itm_6_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_7_land_3_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~((and_dcpl_1566 & FpFractionToFloat_35U_6U_10U_1_and_2_cse
        & (IntLeadZero_35U_1_leading_sign_35_0_rtn_3_sva_2[5]) & (FpFractionToFloat_35U_6U_10U_1_mux_41_tmp[1])
        & (FpFractionToFloat_35U_6U_10U_1_mux_41_tmp[3]) & (~ IsNaN_6U_10U_6_nor_2_tmp))
        | or_2010_cse | (~ main_stage_v_1) | or_dcpl_906)) ) begin
      IsNaN_6U_10U_7_land_3_lpi_1_dfm <= and_3249_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs
          <= 1'b0;
    end
    else if ( core_wen & (~(or_2010_cse | FpMul_6U_10U_2_if_2_FpMul_6U_10U_2_if_2_or_7_tmp
        | (~ main_stage_v_1) | or_dcpl_913)) ) begin
      inp_lookup_4_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs
          <= inp_lookup_4_FpMul_6U_10U_2_else_2_if_acc_itm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_7_land_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~((and_dcpl_1577 & (FpFractionToFloat_35U_6U_10U_1_mux_42_tmp[4:3]==2'b11)
        & (~ IsNaN_6U_10U_6_nor_3_tmp) & inp_lookup_4_FpMantRNE_36U_11U_1_else_and_svs_2
        & (IntLeadZero_35U_1_leading_sign_35_0_rtn_sva_2[5]) & FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2)
        | or_2010_cse | (~ main_stage_v_1) | or_dcpl_913)) ) begin
      IsNaN_6U_10U_7_land_lpi_1_dfm <= and_3361_cse_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1446_nl)) ) begin
      inp_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_6 <= inp_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_5 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1448_nl)) ) begin
      inp_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_5 <= IsZero_6U_10U_5_IsZero_6U_10U_5_and_1_itm_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1450_nl)) ) begin
      inp_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_6 <= inp_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_5;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_5 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1452_nl)) ) begin
      inp_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_5 <= IsZero_6U_10U_5_IsZero_6U_10U_5_and_3_itm_2;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4
          <= 1'b0;
    end
    else if ( core_wen & FpMul_6U_10U_2_oelse_1_FpMul_6U_10U_2_oelse_1_or_11_cse
        & (mux_1455_nl) ) begin
      inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4
          <= MUX_s_1_2_2(inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0,
          inp_lookup_1_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_6, and_dcpl_427);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4
          <= 1'b0;
    end
    else if ( core_wen & IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_2_cse
        & (mux_1458_nl) ) begin
      inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4
          <= MUX_s_1_2_2(inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0,
          inp_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_5, and_dcpl_464);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4
          <= 1'b0;
    end
    else if ( core_wen & IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_1_cse
        & (~ (mux_1461_nl)) ) begin
      inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4
          <= MUX_s_1_2_2(inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0,
          inp_lookup_3_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_6, and_dcpl_496);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4
          <= 1'b0;
    end
    else if ( core_wen & IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_cse
        & (mux_1464_nl) ) begin
      inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4
          <= MUX_s_1_2_2(inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_mx0w0,
          inp_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_itm_5, and_dcpl_535);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_itm_9 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_or_6_cse
        & (~ (mux_1467_nl)) ) begin
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_itm_9 <= MUX_s_1_2_2(FpMul_6U_10U_2_else_2_else_and_itm_2,
          (inp_lookup_1_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_nl), and_dcpl_565);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_1_itm_7 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_or_5_cse
        & (~ (mux_1470_nl)) ) begin
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_1_itm_7 <= MUX_s_1_2_2(FpMul_6U_10U_2_else_2_else_and_1_itm_2,
          (inp_lookup_2_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_nl), and_dcpl_583);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_itm_9 <= 1'b0;
    end
    else if ( core_wen & FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_or_4_cse
        & (~ (mux_1473_nl)) ) begin
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_itm_9 <= MUX_s_1_2_2(FpMul_6U_10U_2_else_2_else_and_2_itm_2,
          (inp_lookup_3_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_nl), and_dcpl_601);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_3_itm_7 <= 1'b0;
    end
    else if ( core_wen & FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_4_cse & (~
        (mux_1475_nl)) ) begin
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_3_itm_7 <= MUX_s_1_2_2(FpMul_6U_10U_2_else_2_else_and_3_itm_2,
          (inp_lookup_4_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_nl), and_dcpl_631);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_8_land_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1482_nl) ) begin
      IsNaN_6U_10U_8_land_lpi_1_dfm_4 <= IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_9_land_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1488_nl) ) begin
      IsNaN_6U_10U_9_land_lpi_1_dfm_6 <= ~(IsNaN_6U_10U_9_nor_3_tmp | (~(FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_5_1
          & FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_4_1 & (FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_3_0_1==4'b1111))));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_8_land_3_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1495_nl) ) begin
      IsNaN_6U_10U_8_land_3_lpi_1_dfm_4 <= IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_9_land_3_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1501_nl) ) begin
      IsNaN_6U_10U_9_land_3_lpi_1_dfm_6 <= ~(IsNaN_6U_10U_9_nor_2_tmp | (~(FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_5_1
          & FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_4_1 & (FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_3_0_1==4'b1111))));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_8_land_2_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1508_nl) ) begin
      IsNaN_6U_10U_8_land_2_lpi_1_dfm_4 <= IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_9_land_2_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1514_nl) ) begin
      IsNaN_6U_10U_9_land_2_lpi_1_dfm_6 <= ~(IsNaN_6U_10U_9_nor_1_tmp | (~(FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_5_1
          & FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_4_1 & (FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_3_0_1==4'b1111))));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_8_land_1_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1521_nl) ) begin
      IsNaN_6U_10U_8_land_1_lpi_1_dfm_6 <= IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_9_land_1_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1527_nl) ) begin
      IsNaN_6U_10U_9_land_1_lpi_1_dfm_6 <= ~(IsNaN_6U_10U_9_nor_tmp | (~(FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_5_1
          & FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_4_1 & (FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_3_0_1==4'b1111))));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_8_283_1 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1529_nl) ) begin
      chn_inp_in_crt_sva_8_283_1 <= chn_inp_in_crt_sva_7_283_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_8_299_1 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1531_nl) ) begin
      chn_inp_in_crt_sva_8_299_1 <= chn_inp_in_crt_sva_7_299_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_8_315_1 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1535_nl) ) begin
      chn_inp_in_crt_sva_8_315_1 <= chn_inp_in_crt_sva_7_315_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_8_331_1 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1539_nl) ) begin
      chn_inp_in_crt_sva_8_331_1 <= chn_inp_in_crt_sva_7_331_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_lpi_1_dfm_9 <= 10'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_5_4_1 <= 1'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_5_3_0_1 <= 4'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_lpi_1_dfm_9 <= 3'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_19_itm_5
          <= 1'b0;
    end
    else if ( FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_12_cse ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_lpi_1_dfm_9 <= MUX_v_10_2_2(({{9{IsInf_6U_23U_1_land_lpi_1_dfm_mx0w0}},
          IsInf_6U_23U_1_land_lpi_1_dfm_mx0w0}), FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_22_13_lpi_1_dfm_mx0w1,
          and_3550_nl);
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_5_4_1 <= FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_4_1
          | IsInf_6U_23U_1_land_lpi_1_dfm_mx0w0 | and_3588_cse;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_lpi_1_dfm_5_3_0_1 <= MUX_v_4_2_2((FpExpoWidthInc_6U_8U_23U_0U_1U_1_mux_44_nl),
          4'b1111, and_3588_cse);
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_lpi_1_dfm_9 <= (FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_15_nl)
          | ({{2{IsInf_6U_23U_1_land_lpi_1_dfm_mx0w0}}, IsInf_6U_23U_1_land_lpi_1_dfm_mx0w0})
          | ({{2{and_3588_cse}}, and_3588_cse});
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_19_itm_5
          <= (IsInf_6U_23U_1_aelse_mux_7_nl) & (~ and_3588_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_2_land_lpi_1_dfm_23 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1547_nl) ) begin
      IsNaN_6U_10U_2_land_lpi_1_dfm_23 <= IsNaN_6U_10U_2_land_lpi_1_dfm_22;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_3_lpi_1_dfm_9 <= 10'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_5_4_1 <= 1'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_5_3_0_1 <= 4'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_3_lpi_1_dfm_9 <= 3'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_14_itm_5
          <= 1'b0;
    end
    else if ( FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_13_cse ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_3_lpi_1_dfm_9 <= MUX_v_10_2_2(({{9{IsInf_6U_23U_1_land_3_lpi_1_dfm_mx0w0}},
          IsInf_6U_23U_1_land_3_lpi_1_dfm_mx0w0}), FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_22_13_3_lpi_1_dfm_mx0w1,
          and_3552_nl);
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_5_4_1 <= FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_4_1
          | IsInf_6U_23U_1_land_3_lpi_1_dfm_mx0w0 | and_3587_cse;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_3_lpi_1_dfm_5_3_0_1 <= MUX_v_4_2_2((FpExpoWidthInc_6U_8U_23U_0U_1U_1_mux_31_nl),
          4'b1111, and_3587_cse);
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_3_lpi_1_dfm_9 <= (FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_10_nl)
          | ({{2{IsInf_6U_23U_1_land_3_lpi_1_dfm_mx0w0}}, IsInf_6U_23U_1_land_3_lpi_1_dfm_mx0w0})
          | ({{2{and_3587_cse}}, and_3587_cse});
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_14_itm_5
          <= (IsInf_6U_23U_1_aelse_mux_5_nl) & (~ and_3587_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_23 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1555_nl) ) begin
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_23 <= IsNaN_6U_10U_2_land_3_lpi_1_dfm_22;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_2_lpi_1_dfm_9 <= 10'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_5_4_1 <= 1'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_5_3_0_1 <= 4'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_2_lpi_1_dfm_9 <= 3'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_9_itm_5
          <= 1'b0;
    end
    else if ( FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_14_cse ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_2_lpi_1_dfm_9 <= MUX_v_10_2_2(({{9{IsInf_6U_23U_1_land_2_lpi_1_dfm_mx0w0}},
          IsInf_6U_23U_1_land_2_lpi_1_dfm_mx0w0}), FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_22_13_2_lpi_1_dfm_mx0w1,
          and_3554_nl);
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_5_4_1 <= FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_4_1
          | IsInf_6U_23U_1_land_2_lpi_1_dfm_mx0w0 | and_3586_cse;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_2_lpi_1_dfm_5_3_0_1 <= MUX_v_4_2_2((FpExpoWidthInc_6U_8U_23U_0U_1U_1_mux_18_nl),
          4'b1111, and_3586_cse);
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_2_lpi_1_dfm_9 <= (FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_5_nl)
          | ({{2{IsInf_6U_23U_1_land_2_lpi_1_dfm_mx0w0}}, IsInf_6U_23U_1_land_2_lpi_1_dfm_mx0w0})
          | ({{2{and_3586_cse}}, and_3586_cse});
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_9_itm_5
          <= (IsInf_6U_23U_1_aelse_mux_3_nl) & (~ and_3586_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_1_lpi_1_dfm_9 <= 10'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_5_4_1 <= 1'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_5_3_0_1 <= 4'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_1_lpi_1_dfm_9 <= 3'b0;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_4_itm_5
          <= 1'b0;
    end
    else if ( FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_and_15_cse ) begin
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_22_13_1_lpi_1_dfm_9 <= MUX_v_10_2_2(({{9{IsInf_6U_23U_1_land_1_lpi_1_dfm_mx0w0}},
          IsInf_6U_23U_1_land_1_lpi_1_dfm_mx0w0}), FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_22_13_1_lpi_1_dfm_mx0w1,
          and_3556_nl);
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_5_4_1 <= FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_4_1
          | IsInf_6U_23U_1_land_1_lpi_1_dfm_mx0w0 | and_3585_cse;
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_4_0_1_lpi_1_dfm_5_3_0_1 <= MUX_v_4_2_2((FpExpoWidthInc_6U_8U_23U_0U_1U_1_mux_48_nl),
          4'b1111, and_3585_cse);
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_expo_7_5_1_lpi_1_dfm_9 <= (FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_nl)
          | ({{2{IsInf_6U_23U_1_land_1_lpi_1_dfm_mx0w0}}, IsInf_6U_23U_1_land_1_lpi_1_dfm_mx0w0})
          | ({{2{and_3585_cse}}, and_3585_cse});
      FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_4_itm_5
          <= (IsInf_6U_23U_1_aelse_mux_1_nl) & (~ and_3585_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_7_17_1_itm <= 8'b0;
    end
    else if ( or_11_cse & core_wen & main_stage_v_8 & (~ (chn_inp_in_crt_sva_8_739_736_1[3]))
        & inp_lookup_else_unequal_tmp_55 ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_7_17_1_itm <= IntShiftRight_69U_6U_32U_obits_fixed_mux1h_25_itm[16:9];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_7_17_1_1_itm <= 9'b0;
    end
    else if ( and_dcpl_2528 & (~ (chn_inp_in_crt_sva_8_739_736_1[3])) & or_11_cse
        ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_7_17_1_1_itm <= IntShiftRight_69U_6U_32U_obits_fixed_mux1h_25_itm[8:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_7_17_1_itm <= 8'b0;
    end
    else if ( or_11_cse & core_wen & main_stage_v_8 & (~ (chn_inp_in_crt_sva_8_739_736_1[2]))
        & inp_lookup_else_unequal_tmp_55 ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_7_17_1_itm <= IntShiftRight_69U_6U_32U_obits_fixed_mux1h_27_itm[16:9];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_7_17_1_1_itm <= 9'b0;
    end
    else if ( and_dcpl_2528 & (~ (chn_inp_in_crt_sva_8_739_736_1[2])) & or_11_cse
        ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_7_17_1_1_itm <= IntShiftRight_69U_6U_32U_obits_fixed_mux1h_27_itm[8:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_7_17_1_itm <= 8'b0;
    end
    else if ( or_11_cse & core_wen & main_stage_v_8 & (~ (chn_inp_in_crt_sva_8_739_736_1[1]))
        & inp_lookup_else_unequal_tmp_55 ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_7_17_1_itm <= IntShiftRight_69U_6U_32U_obits_fixed_mux1h_29_itm[16:9];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_7_17_1_1_itm <= 9'b0;
    end
    else if ( and_dcpl_2528 & (~ (chn_inp_in_crt_sva_8_739_736_1[1])) & or_11_cse
        ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_7_17_1_1_itm <= IntShiftRight_69U_6U_32U_obits_fixed_mux1h_29_itm[8:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_7_17_1_itm <= 8'b0;
    end
    else if ( or_11_cse & core_wen & main_stage_v_8 & (~ (chn_inp_in_crt_sva_8_739_736_1[0]))
        & inp_lookup_else_unequal_tmp_55 ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_7_17_1_itm <= IntShiftRight_69U_6U_32U_obits_fixed_mux1h_31_itm[16:9];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_7_17_1_1_itm <= 9'b0;
    end
    else if ( and_dcpl_2528 & (~ (chn_inp_in_crt_sva_8_739_736_1[0])) & or_11_cse
        ) begin
      reg_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_7_17_1_1_itm <= IntShiftRight_69U_6U_32U_obits_fixed_mux1h_31_itm[8:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_lpi_1_dfm_16 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1564_nl) ) begin
      IntSaturation_51U_32U_o_lpi_1_dfm_16 <= IntSaturation_51U_32U_o_lpi_1_dfm_15;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_3_lpi_1_dfm_16 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1567_nl) ) begin
      IntSaturation_51U_32U_o_3_lpi_1_dfm_16 <= IntSaturation_51U_32U_o_3_lpi_1_dfm_15;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_2_lpi_1_dfm_16 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1570_nl) ) begin
      IntSaturation_51U_32U_o_2_lpi_1_dfm_16 <= IntSaturation_51U_32U_o_2_lpi_1_dfm_15;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_1_lpi_1_dfm_16 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1573_nl) ) begin
      IntSaturation_51U_32U_o_1_lpi_1_dfm_16 <= IntSaturation_51U_32U_o_1_lpi_1_dfm_15;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_19 <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1574_nl) ) begin
      cfg_precision_1_sva_19 <= cfg_precision_1_sva_18;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_485_itm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ mux_1558_itm) ) begin
      inp_lookup_else_mux_485_itm_9 <= inp_lookup_else_mux_485_itm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_491_itm_5 <= 1'b0;
    end
    else if ( core_wen & IntShiftRight_69U_6U_32U_obits_fixed_inp_lookup_else_or_7_cse
        & (~ mux_1558_itm) ) begin
      inp_lookup_else_mux_491_itm_5 <= MUX_s_1_2_2((IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_12[0]),
          (FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_9_0_lpi_1_dfm_2_mx0[0]), and_2194_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_362_itm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ mux_1559_itm) ) begin
      inp_lookup_else_mux_362_itm_9 <= inp_lookup_else_mux_362_itm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_368_itm_5 <= 1'b0;
    end
    else if ( core_wen & IntShiftRight_69U_6U_32U_obits_fixed_inp_lookup_else_or_7_cse
        & (~ mux_1559_itm) ) begin
      inp_lookup_else_mux_368_itm_5 <= MUX_s_1_2_2((IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_12[0]),
          (FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_9_0_3_lpi_1_dfm_2_mx0[0]), and_2194_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_239_itm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ mux_1560_itm) ) begin
      inp_lookup_else_mux_239_itm_9 <= inp_lookup_else_mux_239_itm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_245_itm_5 <= 1'b0;
    end
    else if ( core_wen & IntShiftRight_69U_6U_32U_obits_fixed_inp_lookup_else_or_7_cse
        & (~ mux_1560_itm) ) begin
      inp_lookup_else_mux_245_itm_5 <= MUX_s_1_2_2((IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_12[0]),
          (FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_9_0_2_lpi_1_dfm_2_mx0[0]), and_2194_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_116_itm_9 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ mux_1561_itm) ) begin
      inp_lookup_else_mux_116_itm_9 <= inp_lookup_else_mux_116_itm_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_122_itm_5 <= 1'b0;
    end
    else if ( core_wen & IntShiftRight_69U_6U_32U_obits_fixed_inp_lookup_else_or_7_cse
        & (~ mux_1561_itm) ) begin
      inp_lookup_else_mux_122_itm_5 <= MUX_s_1_2_2((IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_12[0]),
          (FpExpoWidthInc_6U_8U_23U_0U_1U_1_o_mant_9_0_1_lpi_1_dfm_2_mx0[0]), and_2194_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_qr_lpi_1_dfm_3_0 <= 4'b0;
      reg_FpAdd_6U_10U_qr_lpi_1_dfm_5_4_tmp <= 1'b0;
      reg_FpAdd_6U_10U_qr_lpi_1_dfm_5_4_tmp_1 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_and_41_cse ) begin
      FpAdd_6U_10U_qr_lpi_1_dfm_3_0 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_27,
          FpMul_6U_10U_o_expo_lpi_1_dfm_6_3_0_1, and_dcpl_1731);
      reg_FpAdd_6U_10U_qr_lpi_1_dfm_5_4_tmp <= MUX_s_1_2_2(reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_15_tmp,
          reg_FpMul_6U_10U_o_expo_lpi_1_dfm_6_5_4_tmp, and_dcpl_1731);
      reg_FpAdd_6U_10U_qr_lpi_1_dfm_5_4_tmp_1 <= MUX_s_1_2_2(reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_15_tmp_1,
          reg_FpMul_6U_10U_o_expo_lpi_1_dfm_6_5_4_tmp_1, and_dcpl_1731);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_12 <= 18'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1579_nl)) ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_12 <= IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_11;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_12 <= 18'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1580_nl)) ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_12 <= IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_11;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_12 <= 18'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1581_nl)) ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_12 <= IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_11;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_12 <= 18'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1582_nl)) ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_12 <= IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_11;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_3_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_3_0 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_3 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_3_1 <= chn_inp_in_rsci_d_mxwt[346];
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_3_0 <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_3_0_mx0w0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_3 <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_3_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_3_0 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_3 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_3_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_3_1 <= chn_inp_in_rsci_d_mxwt[362];
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_3_0 <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_3_0_mx0w0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_3 <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_3_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_3_0 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_3_lpi_1_dfm_3 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_6_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_3_1 <= chn_inp_in_rsci_d_mxwt[378];
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_3_0 <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_3_0_mx0w0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_3_lpi_1_dfm_3 <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_3_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_3_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_3_0 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_3 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_and_9_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_3_1 <= chn_inp_in_rsci_d_mxwt[394];
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_3_0 <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_3_0_mx0w0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_3 <= FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_7_283_1 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1583_nl) ) begin
      chn_inp_in_crt_sva_7_283_1 <= chn_inp_in_crt_sva_6_283_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_7_331_1 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1584_nl) ) begin
      chn_inp_in_crt_sva_7_331_1 <= chn_inp_in_crt_sva_6_331_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_7_299_1 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1585_nl) ) begin
      chn_inp_in_crt_sva_7_299_1 <= chn_inp_in_crt_sva_6_299_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_7_315_1 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1588_nl) ) begin
      chn_inp_in_crt_sva_7_315_1 <= chn_inp_in_crt_sva_6_315_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_lpi_1_dfm_15 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1590_nl) ) begin
      IntSaturation_51U_32U_o_lpi_1_dfm_15 <= IntSaturation_51U_32U_o_lpi_1_dfm_14;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_3_lpi_1_dfm_15 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1592_nl) ) begin
      IntSaturation_51U_32U_o_3_lpi_1_dfm_15 <= IntSaturation_51U_32U_o_3_lpi_1_dfm_14;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_2_lpi_1_dfm_15 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1595_nl) ) begin
      IntSaturation_51U_32U_o_2_lpi_1_dfm_15 <= IntSaturation_51U_32U_o_2_lpi_1_dfm_14;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_1_lpi_1_dfm_15 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1597_nl) ) begin
      IntSaturation_51U_32U_o_1_lpi_1_dfm_15 <= IntSaturation_51U_32U_o_1_lpi_1_dfm_14;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_18 <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1598_nl) ) begin
      cfg_precision_1_sva_18 <= cfg_precision_1_sva_17;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_485_itm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1599_nl)) ) begin
      inp_lookup_else_mux_485_itm_8 <= inp_lookup_else_mux_485_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_362_itm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1600_nl)) ) begin
      inp_lookup_else_mux_362_itm_8 <= inp_lookup_else_mux_362_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_239_itm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1601_nl)) ) begin
      inp_lookup_else_mux_239_itm_8 <= inp_lookup_else_mux_239_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_116_itm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1602_nl)) ) begin
      inp_lookup_else_mux_116_itm_8 <= inp_lookup_else_mux_116_itm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsInf_6U_23U_1_land_1_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_295 | and_dcpl_78 | (chn_inp_in_crt_sva_8_739_736_1[0])))
        ) begin
      IsInf_6U_23U_1_land_1_lpi_1_dfm <= IsInf_6U_23U_1_land_1_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsInf_6U_23U_1_land_2_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(nand_544_cse | (chn_inp_in_crt_sva_8_739_736_1[1]) |
        and_dcpl_78 | (cfg_precision_1_sva_st_85[0]))) ) begin
      IsInf_6U_23U_1_land_2_lpi_1_dfm <= IsInf_6U_23U_1_land_2_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsInf_6U_23U_1_land_3_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_295 | and_dcpl_78 | (chn_inp_in_crt_sva_8_739_736_1[2])))
        ) begin
      IsInf_6U_23U_1_land_3_lpi_1_dfm <= IsInf_6U_23U_1_land_3_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsInf_6U_23U_1_land_lpi_1_dfm <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_295 | and_dcpl_78 | (chn_inp_in_crt_sva_8_739_736_1[3])))
        ) begin
      IsInf_6U_23U_1_land_lpi_1_dfm <= IsInf_6U_23U_1_land_lpi_1_dfm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_3 <= 10'b0;
    end
    else if ( core_wen & ((and_dcpl_1760 & and_dcpl_1758 & (fsm_output[1])) | (and_dcpl_1764
        & and_dcpl_1758) | FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_3_mx0c1)
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_3 <= MUX_v_10_2_2((chn_inp_in_rsci_d_mxwt[341:332]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_or_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_3_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_3 <= 10'b0;
    end
    else if ( core_wen & ((and_dcpl_1773 & and_dcpl_1772 & (fsm_output[1])) | (and_dcpl_1777
        & and_dcpl_1772) | FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_3_mx0c1)
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_3 <= MUX_v_10_2_2((chn_inp_in_rsci_d_mxwt[357:348]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_or_4_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_3_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_3_lpi_1_dfm_3 <= 10'b0;
    end
    else if ( core_wen & ((and_dcpl_1786 & and_dcpl_1785 & (fsm_output[1])) | (and_dcpl_1790
        & and_dcpl_1785) | FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_3_lpi_1_dfm_3_mx0c1)
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_3_lpi_1_dfm_3 <= MUX_v_10_2_2((chn_inp_in_rsci_d_mxwt[373:364]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_or_8_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_3_lpi_1_dfm_3_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_3 <= 10'b0;
    end
    else if ( core_wen & ((and_dcpl_1799 & and_dcpl_1798 & (fsm_output[1])) | (and_dcpl_1803
        & and_dcpl_1798) | FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_3_mx0c1)
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_3 <= MUX_v_10_2_2((chn_inp_in_rsci_d_mxwt[389:380]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_FpExpoWidthInc_5U_6U_10U_1U_1U_3_or_12_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_3_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_itm_8 <= 1'b0;
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_itm_8 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_19 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_19 <= 10'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_19 <= 10'b0;
    end
    else if ( IsZero_6U_10U_1_and_12_cse ) begin
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_itm_8 <= IsZero_6U_10U_1_IsZero_6U_10U_1_and_itm_7;
      IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_itm_8 <= IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_itm_7;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_19 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_18;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_19 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_18;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_19 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_18;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_22 <= 10'b0;
    end
    else if ( core_wen & FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_3_cse & (mux_1605_nl)
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_22 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_21,
          FpMul_6U_10U_1_FpMul_6U_10U_1_FpMul_6U_10U_1_nor_4_itm, FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_46_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_22 <= 10'b0;
    end
    else if ( core_wen & FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_2_cse & (mux_1608_nl)
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_22 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_21,
          FpMul_6U_10U_1_FpMul_6U_10U_1_FpMul_6U_10U_1_nor_5_itm, FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_45_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_22 <= 10'b0;
    end
    else if ( core_wen & IsNaN_8U_23U_2_aelse_IsNaN_8U_23U_2_aelse_or_cse & (mux_1612_nl)
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_22 <= MUX_v_10_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_21,
          FpMul_6U_10U_1_FpMul_6U_10U_1_FpMul_6U_10U_1_nor_7_itm, FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_44_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_6_283_1 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1613_nl) ) begin
      chn_inp_in_crt_sva_6_283_1 <= chn_inp_in_crt_sva_5_283_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_6_299_1 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1614_nl) ) begin
      chn_inp_in_crt_sva_6_299_1 <= chn_inp_in_crt_sva_5_299_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_6_315_1 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1615_nl) ) begin
      chn_inp_in_crt_sva_6_315_1 <= chn_inp_in_crt_sva_5_315_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_6_331_1 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1616_nl) ) begin
      chn_inp_in_crt_sva_6_331_1 <= chn_inp_in_crt_sva_5_331_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_11 <= 18'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1617_nl)) ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_11 <= IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_11 <= 18'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1618_nl)) ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_11 <= IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_11 <= 18'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1619_nl)) ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_11 <= IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_11 <= 18'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1620_nl)) ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_11 <= IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_10;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_lpi_1_dfm_14 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1622_nl) ) begin
      IntSaturation_51U_32U_o_lpi_1_dfm_14 <= IntSaturation_51U_32U_o_lpi_1_dfm_13;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_3_lpi_1_dfm_14 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1624_nl) ) begin
      IntSaturation_51U_32U_o_3_lpi_1_dfm_14 <= IntSaturation_51U_32U_o_3_lpi_1_dfm_13;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_2_lpi_1_dfm_14 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1629_nl) ) begin
      IntSaturation_51U_32U_o_2_lpi_1_dfm_14 <= IntSaturation_51U_32U_o_2_lpi_1_dfm_13;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_1_lpi_1_dfm_14 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1632_nl) ) begin
      IntSaturation_51U_32U_o_1_lpi_1_dfm_14 <= IntSaturation_51U_32U_o_1_lpi_1_dfm_13;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_17 <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1633_nl) ) begin
      cfg_precision_1_sva_17 <= cfg_precision_1_sva_16;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_485_itm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1634_nl)) ) begin
      inp_lookup_else_mux_485_itm_7 <= inp_lookup_else_mux_485_itm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_362_itm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1635_nl)) ) begin
      inp_lookup_else_mux_362_itm_7 <= inp_lookup_else_mux_362_itm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_239_itm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1636_nl)) ) begin
      inp_lookup_else_mux_239_itm_7 <= inp_lookup_else_mux_239_itm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_116_itm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1637_nl)) ) begin
      inp_lookup_else_mux_116_itm_7 <= inp_lookup_else_mux_116_itm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_21 <= 10'b0;
    end
    else if ( core_wen & (and_2284_rgt | and_2287_rgt | and_2289_rgt) & (mux_1640_nl)
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_21 <= MUX1HOT_v_10_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_20,
          (FpMul_6U_10U_1_p_mant_20_1_1_lpi_1_dfm_3_mx0[19:10]), inp_lookup_else_if_a0_9_0_1_lpi_1_dfm_10,
          {and_2284_rgt , and_2287_rgt , and_2289_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_21 <= 10'b0;
    end
    else if ( core_wen & (and_2291_rgt | and_2294_rgt | and_2296_rgt) & (mux_1643_nl)
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_21 <= MUX1HOT_v_10_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_20,
          (FpMul_6U_10U_1_p_mant_20_1_2_lpi_1_dfm_3_mx0[19:10]), inp_lookup_else_if_a0_9_0_2_lpi_1_dfm_10,
          {and_2291_rgt , and_2294_rgt , and_2296_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_21 <= 10'b0;
    end
    else if ( core_wen & (and_2298_rgt | and_2301_rgt | and_2303_rgt) & (mux_1646_nl)
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_21 <= MUX1HOT_v_10_3_2(FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_20,
          (FpMul_6U_10U_1_p_mant_20_1_lpi_1_dfm_3_mx0[19:10]), inp_lookup_else_if_a0_9_0_lpi_1_dfm_10,
          {and_2298_rgt , and_2301_rgt , and_2303_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_5_283_1 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1647_nl) ) begin
      chn_inp_in_crt_sva_5_283_1 <= chn_inp_in_crt_sva_4_283_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_5_331_1 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1648_nl) ) begin
      chn_inp_in_crt_sva_5_331_1 <= chn_inp_in_crt_sva_4_331_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_5_299_1 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1649_nl) ) begin
      chn_inp_in_crt_sva_5_299_1 <= chn_inp_in_crt_sva_4_299_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_5_315_1 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1650_nl) ) begin
      chn_inp_in_crt_sva_5_315_1 <= chn_inp_in_crt_sva_4_315_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_o_sign_1_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & (or_5766_rgt | or_5767_rgt | and_dcpl_655) & not_tmp_1029
        ) begin
      FpAdd_8U_23U_1_o_sign_1_lpi_1_dfm_5 <= MUX1HOT_s_1_3_2((chn_inp_in_crt_sva_4_127_0_1[31]),
          (~ FpAdd_8U_23U_o_sign_1_lpi_1_dfm_8), FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_3_4_mx1w1,
          {or_5766_rgt , or_5767_rgt , and_dcpl_655});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_o_sign_2_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & (or_5764_rgt | or_5765_rgt | and_dcpl_663) & not_tmp_1046
        ) begin
      FpAdd_8U_23U_1_o_sign_2_lpi_1_dfm_5 <= MUX1HOT_s_1_3_2((chn_inp_in_crt_sva_4_127_0_1[63]),
          (~ FpAdd_8U_23U_o_sign_2_lpi_1_dfm_8), FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_3_4_mx1w1,
          {or_5764_rgt , or_5765_rgt , and_dcpl_663});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_o_sign_3_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & (or_5762_rgt | or_5763_rgt | and_dcpl_671) & not_tmp_1063
        ) begin
      FpAdd_8U_23U_1_o_sign_3_lpi_1_dfm_5 <= MUX1HOT_s_1_3_2((chn_inp_in_crt_sva_4_127_0_1[95]),
          (~ FpAdd_8U_23U_o_sign_3_lpi_1_dfm_9), FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_4_mx1w1,
          {or_5762_rgt , or_5763_rgt , and_dcpl_671});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_1_o_sign_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( core_wen & (or_5760_rgt | or_5761_rgt | and_dcpl_679) & not_tmp_1080
        ) begin
      FpAdd_8U_23U_1_o_sign_lpi_1_dfm_5 <= MUX1HOT_s_1_3_2((chn_inp_in_crt_sva_4_127_0_1[127]),
          (~ FpAdd_8U_23U_o_sign_lpi_1_dfm_9), FpMul_6U_10U_1_o_expo_lpi_1_dfm_3_4_mx0w1,
          {or_5760_rgt , or_5761_rgt , and_dcpl_679});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_10 <= 18'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1652_nl)) ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_10 <= IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_10 <= 18'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1654_nl)) ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_10 <= IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_10 <= 18'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1656_nl)) ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_10 <= IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_10 <= 18'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1658_nl)) ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_10 <= IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_9;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_lpi_1_dfm_13 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1660_nl) ) begin
      IntSaturation_51U_32U_o_lpi_1_dfm_13 <= IntSaturation_51U_32U_o_lpi_1_dfm_12;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_3_lpi_1_dfm_13 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1662_nl) ) begin
      IntSaturation_51U_32U_o_3_lpi_1_dfm_13 <= IntSaturation_51U_32U_o_3_lpi_1_dfm_12;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_2_lpi_1_dfm_13 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1664_nl) ) begin
      IntSaturation_51U_32U_o_2_lpi_1_dfm_13 <= IntSaturation_51U_32U_o_2_lpi_1_dfm_12;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_1_lpi_1_dfm_13 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1666_nl) ) begin
      IntSaturation_51U_32U_o_1_lpi_1_dfm_13 <= IntSaturation_51U_32U_o_1_lpi_1_dfm_12;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_precision_1_sva_16 <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1667_nl) ) begin
      cfg_precision_1_sva_16 <= cfg_precision_1_sva_st_82;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_485_itm_6 <= 1'b0;
    end
    else if ( core_wen & (and_2320_cse | IntShiftRight_69U_6U_32U_obits_fixed_or_6_rgt
        | IntShiftRight_69U_6U_32U_obits_fixed_or_7_rgt) & (~ (mux_1668_nl)) ) begin
      inp_lookup_else_mux_485_itm_6 <= MUX1HOT_s_1_3_2((IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_9[17]),
          FpMul_6U_10U_2_o_sign_lpi_1_dfm_8, FpMul_6U_10U_1_o_sign_lpi_1_dfm_8, {and_2320_cse
          , IntShiftRight_69U_6U_32U_obits_fixed_or_6_rgt , IntShiftRight_69U_6U_32U_obits_fixed_or_7_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_362_itm_6 <= 1'b0;
    end
    else if ( core_wen & (and_2320_cse | IntShiftRight_69U_6U_32U_obits_fixed_or_4_rgt
        | IntShiftRight_69U_6U_32U_obits_fixed_or_5_rgt) & (~ (mux_1669_nl)) ) begin
      inp_lookup_else_mux_362_itm_6 <= MUX1HOT_s_1_3_2((IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_9[17]),
          FpMul_6U_10U_2_o_sign_3_lpi_1_dfm_8, FpMul_6U_10U_1_o_sign_3_lpi_1_dfm_8,
          {and_2320_cse , IntShiftRight_69U_6U_32U_obits_fixed_or_4_rgt , IntShiftRight_69U_6U_32U_obits_fixed_or_5_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_239_itm_6 <= 1'b0;
    end
    else if ( core_wen & (and_2320_cse | IntShiftRight_69U_6U_32U_obits_fixed_or_2_rgt
        | IntShiftRight_69U_6U_32U_obits_fixed_or_3_rgt) & (~ (mux_1670_nl)) ) begin
      inp_lookup_else_mux_239_itm_6 <= MUX1HOT_s_1_3_2((IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_9[17]),
          FpMul_6U_10U_2_o_sign_2_lpi_1_dfm_8, FpMul_6U_10U_1_o_sign_2_lpi_1_dfm_8,
          {and_2320_cse , IntShiftRight_69U_6U_32U_obits_fixed_or_2_rgt , IntShiftRight_69U_6U_32U_obits_fixed_or_3_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_else_mux_116_itm_6 <= 1'b0;
    end
    else if ( core_wen & (and_2320_cse | IntShiftRight_69U_6U_32U_obits_fixed_or_rgt
        | IntShiftRight_69U_6U_32U_obits_fixed_or_1_rgt) & (~ (mux_1671_nl)) ) begin
      inp_lookup_else_mux_116_itm_6 <= MUX1HOT_s_1_3_2((IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_9[17]),
          FpMul_6U_10U_2_o_sign_1_lpi_1_dfm_8, FpMul_6U_10U_1_o_sign_1_lpi_1_dfm_8,
          {and_2320_cse , IntShiftRight_69U_6U_32U_obits_fixed_or_rgt , IntShiftRight_69U_6U_32U_obits_fixed_or_1_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_9 <= 18'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1673_nl)) ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_9 <= IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_9 <= 18'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1675_nl)) ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_9 <= IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_9 <= 18'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1677_nl)) ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_9 <= IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_9 <= 18'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1679_nl)) ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_9 <= IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_8;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_6_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_6_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_15 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_6_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_6_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_18 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_100_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_6_1_1 <= MUX_s_1_2_2((chn_inp_in_rsci_d_mxwt[410]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3_1, and_dcpl_1854);
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_6_0_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3_0_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3_0, and_dcpl_1854);
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_15 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3, and_dcpl_1854);
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_6_1_1 <= MUX_s_1_2_2((chn_inp_in_rsci_d_mxwt[282]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_3_1, and_dcpl_1854);
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_6_0_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_3_0_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_3_0, and_dcpl_1854);
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_18 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_3, and_dcpl_1854);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_6_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_6_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_15 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_6_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_6_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_18 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_103_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_6_1_1 <= MUX_s_1_2_2((chn_inp_in_rsci_d_mxwt[426]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3_1, and_dcpl_1857);
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_6_0_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3_0_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3_0, and_dcpl_1857);
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_15 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3, and_dcpl_1857);
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_6_1_1 <= MUX_s_1_2_2((chn_inp_in_rsci_d_mxwt[298]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_3_1, and_dcpl_1857);
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_6_0_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_3_0_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_3_0, and_dcpl_1857);
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_18 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_3, and_dcpl_1857);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_6_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_6_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_15 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_6_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_6_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_18 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_106_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_6_1_1 <= MUX_s_1_2_2((chn_inp_in_rsci_d_mxwt[442]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3_1, and_dcpl_1860);
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_6_0_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3_0_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3_0, and_dcpl_1860);
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_15 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3, and_dcpl_1860);
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_6_1_1 <= MUX_s_1_2_2((chn_inp_in_rsci_d_mxwt[314]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_3_1, and_dcpl_1860);
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_6_0_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_3_0_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_3_0, and_dcpl_1860);
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_18 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_3, and_dcpl_1860);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_6_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_6_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_15 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_6_1_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_6_0_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_18 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_109_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_6_1_1 <= MUX_s_1_2_2((chn_inp_in_rsci_d_mxwt[458]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3_1, and_dcpl_1863);
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_6_0_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3_0_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3_0, and_dcpl_1863);
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_15 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_3, and_dcpl_1863);
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_6_1_1 <= MUX_s_1_2_2((chn_inp_in_rsci_d_mxwt[330]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_3_1, and_dcpl_1863);
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_6_0_1 <= MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_3_0_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_3_0, and_dcpl_1863);
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_18 <= MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_3_mx0w0,
          FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_3, and_dcpl_1863);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_20 <= 10'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1682_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_20 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_19;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_20 <= 10'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1685_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_20 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_19;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_20 <= 10'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1688_nl) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_20 <= FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_19;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_4_283_1 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1689_nl) ) begin
      chn_inp_in_crt_sva_4_283_1 <= chn_inp_in_crt_sva_3_331_268_1[15];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_4_331_1 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1691_nl) ) begin
      chn_inp_in_crt_sva_4_331_1 <= chn_inp_in_crt_sva_3_331_268_1[63];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_4_299_1 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1692_nl) ) begin
      chn_inp_in_crt_sva_4_299_1 <= chn_inp_in_crt_sva_3_331_268_1[31];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_inp_in_crt_sva_4_315_1 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1693_nl) ) begin
      chn_inp_in_crt_sva_4_315_1 <= chn_inp_in_crt_sva_3_331_268_1[47];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_11 <= 1'b0;
    end
    else if ( core_wen & FpMul_6U_10U_1_oelse_1_IsNaN_8U_23U_2_aelse_or_4_cse & (~
        (mux_1697_nl)) ) begin
      inp_lookup_4_FpAdd_6U_10U_IsZero_6U_10U_2_nand_itm_11 <= MUX_s_1_2_2(FpMul_6U_10U_2_lor_1_lpi_1_dfm_st_4,
          (inp_lookup_4_FpMul_6U_10U_1_p_mant_p1_mul_tmp[21]), and_dcpl_631);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_o_sign_1_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (((IsNaN_6U_10U_5_land_1_lpi_1_dfm_5 ^ (chn_inp_in_crt_sva_3_739_736_1[0]))
        & or_11_cse) | and_2342_rgt) & (mux_1703_nl) ) begin
      FpAdd_8U_23U_o_sign_1_lpi_1_dfm_8 <= MUX_s_1_2_2(FpAdd_8U_23U_o_sign_1_lpi_1_dfm_5,
          FpMantRNE_22U_11U_1_else_carry_1_sva, and_2342_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_o_sign_2_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (((IsNaN_6U_10U_5_land_2_lpi_1_dfm_5 ^ (chn_inp_in_crt_sva_3_739_736_1[1]))
        & or_11_cse) | and_2345_rgt) & (~ (mux_1711_nl)) ) begin
      FpAdd_8U_23U_o_sign_2_lpi_1_dfm_8 <= MUX_s_1_2_2(FpAdd_8U_23U_o_sign_2_lpi_1_dfm_5,
          FpMantRNE_22U_11U_1_else_carry_2_sva, and_2345_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_o_sign_3_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (((IsNaN_6U_10U_5_land_3_lpi_1_dfm_5 ^ (chn_inp_in_crt_sva_3_739_736_1[2]))
        & or_11_cse) | and_2348_rgt) & (~ (mux_1719_nl)) ) begin
      FpAdd_8U_23U_o_sign_3_lpi_1_dfm_9 <= MUX_s_1_2_2(FpAdd_8U_23U_o_sign_3_lpi_1_dfm_8,
          FpMantRNE_22U_11U_1_else_carry_3_sva, and_2348_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_o_sign_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_630 | and_2350_rgt | and_2351_rgt) & (mux_1729_nl)
        ) begin
      FpAdd_8U_23U_o_sign_lpi_1_dfm_9 <= MUX1HOT_s_1_3_2(FpAdd_8U_23U_o_sign_lpi_1_dfm_8,
          FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_8_0, FpMantRNE_22U_11U_1_else_carry_sva_mx0w1,
          {and_dcpl_630 , and_2350_rgt , and_2351_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_lpi_1_dfm_12 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1731_nl) ) begin
      IntSaturation_51U_32U_o_lpi_1_dfm_12 <= IntSaturation_51U_32U_o_lpi_1_dfm_11;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_3_lpi_1_dfm_12 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1733_nl) ) begin
      IntSaturation_51U_32U_o_3_lpi_1_dfm_12 <= IntSaturation_51U_32U_o_3_lpi_1_dfm_11;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_2_lpi_1_dfm_12 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1735_nl) ) begin
      IntSaturation_51U_32U_o_2_lpi_1_dfm_12 <= IntSaturation_51U_32U_o_2_lpi_1_dfm_11;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_1_lpi_1_dfm_12 <= 32'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1737_nl) ) begin
      IntSaturation_51U_32U_o_1_lpi_1_dfm_12 <= IntSaturation_51U_32U_o_1_lpi_1_dfm_11;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_o_sign_1_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1744_nl) ) begin
      FpMul_6U_10U_2_o_sign_1_lpi_1_dfm_8 <= FpMul_6U_10U_2_o_sign_1_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_sign_1_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1752_nl) ) begin
      FpMul_6U_10U_1_o_sign_1_lpi_1_dfm_8 <= FpMul_6U_10U_1_o_sign_1_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_o_sign_2_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1759_nl) ) begin
      FpMul_6U_10U_2_o_sign_2_lpi_1_dfm_8 <= FpMul_6U_10U_2_o_sign_2_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_sign_2_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1767_nl) ) begin
      FpMul_6U_10U_1_o_sign_2_lpi_1_dfm_8 <= FpMul_6U_10U_1_o_sign_2_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_o_sign_3_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1774_nl) ) begin
      FpMul_6U_10U_2_o_sign_3_lpi_1_dfm_8 <= FpMul_6U_10U_2_o_sign_3_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_sign_3_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1782_nl) ) begin
      FpMul_6U_10U_1_o_sign_3_lpi_1_dfm_8 <= FpMul_6U_10U_1_o_sign_3_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_2_o_sign_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1789_nl) ) begin
      FpMul_6U_10U_2_o_sign_lpi_1_dfm_8 <= FpMul_6U_10U_2_o_sign_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMul_6U_10U_1_o_sign_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1797_nl) ) begin
      FpMul_6U_10U_1_o_sign_lpi_1_dfm_8 <= FpMul_6U_10U_1_o_sign_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_o_sign_1_lpi_1_dfm_5 <= 1'b0;
      FpAdd_8U_23U_o_sign_2_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( FpAdd_8U_23U_o_sign_and_cse ) begin
      FpAdd_8U_23U_o_sign_1_lpi_1_dfm_5 <= FpAdd_8U_23U_o_sign_1_lpi_1_dfm_7;
      FpAdd_8U_23U_o_sign_2_lpi_1_dfm_5 <= FpAdd_8U_23U_o_sign_2_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_o_sign_3_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1802_nl)) ) begin
      FpAdd_8U_23U_o_sign_3_lpi_1_dfm_8 <= FpAdd_8U_23U_o_sign_3_lpi_1_dfm_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3_0 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_3_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_3_0 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_3 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3_1 <= chn_inp_in_rsci_d_mxwt[426];
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3_0 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3_0_mx0w0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_3_1 <= chn_inp_in_rsci_d_mxwt[298];
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_3_0 <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_3_0_mx0w0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_3 <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_2_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3_0 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_3_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_3_0 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_3 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_3_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3_1 <= chn_inp_in_rsci_d_mxwt[458];
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3_0 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3_0_mx0w0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_3 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_3_1 <= chn_inp_in_rsci_d_mxwt[330];
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_3_0 <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_3_0_mx0w0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_3 <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_15 <= 10'b0;
    end
    else if ( core_wen & (and_2358_rgt | and_2359_rgt | and_dcpl_1854) & mux_tmp_6
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_15 <= MUX1HOT_v_10_3_2((chn_inp_in_rsci_d_mxwt[405:396]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_3, {and_2358_rgt , and_2359_rgt
          , and_dcpl_1854});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_15 <= 10'b0;
    end
    else if ( core_wen & (and_2367_rgt | and_2368_rgt | and_dcpl_1857) & mux_tmp_6
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_15 <= MUX1HOT_v_10_3_2((chn_inp_in_rsci_d_mxwt[421:412]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_4_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_3, {and_2367_rgt , and_2368_rgt
          , and_dcpl_1857});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_15 <= 10'b0;
    end
    else if ( core_wen & (and_2375_rgt | and_2376_rgt | and_dcpl_1860) & mux_tmp_6
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_15 <= MUX1HOT_v_10_3_2((chn_inp_in_rsci_d_mxwt[437:428]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_8_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_3, {and_2375_rgt , and_2376_rgt
          , and_dcpl_1860});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_15 <= 10'b0;
    end
    else if ( core_wen & (and_2384_rgt | and_2385_rgt | and_dcpl_1863) & mux_tmp_6
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_15 <= MUX1HOT_v_10_3_2((chn_inp_in_rsci_d_mxwt[453:444]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_12_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_3, {and_2384_rgt , and_2385_rgt
          , and_dcpl_1863});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_8 <= 18'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1805_nl)) ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_8 <= IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_lpi_1_dfm_11 <= 32'b0;
    end
    else if ( core_wen & (IntSaturation_51U_32U_o_IntSaturation_51U_32U_o_nor_rgt
        | IntSaturation_51U_32U_and_7_rgt | IntSaturation_51U_32U_o_and_7_rgt) &
        (mux_1808_nl) ) begin
      IntSaturation_51U_32U_o_lpi_1_dfm_11 <= MUX1HOT_v_32_3_2((inp_lookup_if_else_o_acc_psp_sva[31:0]),
          32'b10000000000000000000000000000000, 32'b1111111111111111111111111111111,
          {IntSaturation_51U_32U_o_IntSaturation_51U_32U_o_nor_rgt , IntSaturation_51U_32U_and_7_rgt
          , IntSaturation_51U_32U_o_and_7_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_8 <= 18'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1810_nl)) ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_8 <= IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_3_lpi_1_dfm_11 <= 32'b0;
    end
    else if ( core_wen & (IntSaturation_51U_32U_o_IntSaturation_51U_32U_o_nor_1_rgt
        | IntSaturation_51U_32U_and_5_rgt | IntSaturation_51U_32U_o_and_5_rgt) &
        (mux_1812_nl) ) begin
      IntSaturation_51U_32U_o_3_lpi_1_dfm_11 <= MUX1HOT_v_32_3_2((inp_lookup_if_else_o_acc_psp_3_sva[31:0]),
          32'b10000000000000000000000000000000, 32'b1111111111111111111111111111111,
          {IntSaturation_51U_32U_o_IntSaturation_51U_32U_o_nor_1_rgt , IntSaturation_51U_32U_and_5_rgt
          , IntSaturation_51U_32U_o_and_5_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_8 <= 18'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1814_nl)) ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_8 <= IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_2_lpi_1_dfm_11 <= 32'b0;
    end
    else if ( core_wen & (IntSaturation_51U_32U_o_IntSaturation_51U_32U_o_nor_2_rgt
        | IntSaturation_51U_32U_and_3_rgt | IntSaturation_51U_32U_o_and_3_rgt) &
        (mux_1816_nl) ) begin
      IntSaturation_51U_32U_o_2_lpi_1_dfm_11 <= MUX1HOT_v_32_3_2((inp_lookup_if_else_o_acc_psp_2_sva[31:0]),
          32'b10000000000000000000000000000000, 32'b1111111111111111111111111111111,
          {IntSaturation_51U_32U_o_IntSaturation_51U_32U_o_nor_2_rgt , IntSaturation_51U_32U_and_3_rgt
          , IntSaturation_51U_32U_o_and_3_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_8 <= 18'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1818_nl)) ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_8 <= IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_7;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_51U_32U_o_1_lpi_1_dfm_11 <= 32'b0;
    end
    else if ( core_wen & (IntSaturation_51U_32U_o_IntSaturation_51U_32U_o_nor_3_rgt
        | IntSaturation_51U_32U_and_1_rgt | IntSaturation_51U_32U_o_and_1_rgt) &
        (mux_1820_nl) ) begin
      IntSaturation_51U_32U_o_1_lpi_1_dfm_11 <= MUX1HOT_v_32_3_2((inp_lookup_if_else_o_acc_psp_1_sva[31:0]),
          32'b10000000000000000000000000000000, 32'b1111111111111111111111111111111,
          {IntSaturation_51U_32U_o_IntSaturation_51U_32U_o_nor_3_rgt , IntSaturation_51U_32U_and_1_rgt
          , IntSaturation_51U_32U_o_and_1_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_18 <= 10'b0;
    end
    else if ( core_wen & ((or_11_cse & (chn_inp_in_rsci_d_mxwt[282:278]==5'b11111)
        & IsDenorm_5U_10U_2_or_tmp) | and_2392_rgt) & (~ mux_93_cse) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_1_lpi_1_dfm_18 <= MUX_v_10_2_2((chn_inp_in_rsci_d_mxwt[277:268]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_or_mx0w1,
          and_2392_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_18 <= 10'b0;
    end
    else if ( core_wen & ((or_11_cse & (chn_inp_in_rsci_d_mxwt[298:294]==5'b11111)
        & IsDenorm_5U_10U_2_or_1_tmp) | and_2399_rgt) & (~ mux_93_cse) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_2_lpi_1_dfm_18 <= MUX_v_10_2_2((chn_inp_in_rsci_d_mxwt[293:284]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_or_4_mx0w1,
          and_2399_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_18 <= 10'b0;
    end
    else if ( core_wen & (and_2404_rgt | and_2405_rgt | and_dcpl_1860) & mux_tmp_6
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_18 <= MUX1HOT_v_10_3_2((chn_inp_in_rsci_d_mxwt[309:300]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_or_8_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_3, {and_2404_rgt ,
          and_2405_rgt , and_dcpl_1860});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_18 <= 10'b0;
    end
    else if ( core_wen & ((or_11_cse & (chn_inp_in_rsci_d_mxwt[330:326]==5'b11111)
        & IsDenorm_5U_10U_2_or_3_tmp) | and_2412_rgt) & (~ mux_93_cse) ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_lpi_1_dfm_18 <= MUX_v_10_2_2((chn_inp_in_rsci_d_mxwt[325:316]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_or_12_mx0w1,
          and_2412_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_o_sign_1_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_1230 | and_dcpl_1232 | and_dcpl_393) & (~ (mux_1824_nl))
        ) begin
      FpAdd_8U_23U_o_sign_1_lpi_1_dfm_7 <= MUX1HOT_s_1_3_2((chn_inp_in_crt_sva_1_739_395_1[116]),
          FpAdd_8U_23U_else_6_mux_mx0w1, FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_6_0_1,
          {and_dcpl_1230 , and_dcpl_1232 , and_dcpl_393});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_o_sign_2_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (and_2414_rgt | and_2416_rgt | and_dcpl_401) & (~ (mux_1828_nl))
        ) begin
      FpAdd_8U_23U_o_sign_2_lpi_1_dfm_7 <= MUX1HOT_s_1_3_2((chn_inp_in_crt_sva_1_739_395_1[148]),
          FpAdd_8U_23U_else_6_mux_3_mx0w1, FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_6_0_1,
          {and_2414_rgt , and_2416_rgt , and_dcpl_401});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_o_sign_3_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_1224 | and_dcpl_1226 | and_dcpl_409) & (~ (mux_1831_nl))
        ) begin
      FpAdd_8U_23U_o_sign_3_lpi_1_dfm_7 <= MUX1HOT_s_1_3_2((chn_inp_in_crt_sva_1_739_395_1[180]),
          FpAdd_8U_23U_else_6_mux_6_mx0w1, FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_6_0_1,
          {and_dcpl_1224 , and_dcpl_1226 , and_dcpl_409});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_o_sign_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (and_2417_rgt | and_2418_rgt | and_2419_rgt) & mux_tmp_50
        ) begin
      FpAdd_8U_23U_o_sign_lpi_1_dfm_7 <= MUX1HOT_s_1_3_2((chn_inp_in_crt_sva_1_739_395_1[212]),
          FpAdd_8U_23U_else_6_mux_9_mx0w1, FpAdd_8U_23U_o_sign_lpi_1_dfm_1, {and_2417_rgt
          , and_2418_rgt , and_2419_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_7 <= 18'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1833_nl)) ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_7 <= nl_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_7[17:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_7 <= 18'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1835_nl)) ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_7 <= nl_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_7[17:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_7 <= 18'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1837_nl)) ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_7 <= nl_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_7[17:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_7 <= 18'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (~ (mux_1840_nl)) ) begin
      IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_7 <= nl_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_7[17:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_8U_23U_o_sign_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( core_wen & (FpAdd_8U_23U_o_sign_lpi_1_dfm_1_mx0c0 | FpAdd_8U_23U_o_sign_lpi_1_dfm_1_mx0c1
        | FpAdd_8U_23U_o_sign_lpi_1_dfm_1_mx0c2) ) begin
      FpAdd_8U_23U_o_sign_lpi_1_dfm_1 <= MUX1HOT_s_1_3_2((chn_inp_in_crt_sva_1_739_395_1[212]),
          FpAdd_8U_23U_else_6_mux_9_mx0w1, (inp_lookup_4_IsZero_6U_10U_1_IsZero_6U_10U_1_nor_nl),
          {FpAdd_8U_23U_o_sign_lpi_1_dfm_1_mx0c0 , FpAdd_8U_23U_o_sign_lpi_1_dfm_1_mx0c1
          , FpAdd_8U_23U_o_sign_lpi_1_dfm_1_mx0c2});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_3 <= 10'b0;
    end
    else if ( core_wen & ((and_dcpl_1961 & IsDenorm_5U_10U_or_tmp & (chn_inp_in_rsci_d_mxwt[407:406]==2'b11)
        & and_dcpl_1957 & (fsm_output[1])) | (and_dcpl_1759 & (chn_inp_in_rsci_d_mxwt[736])
        & IsDenorm_5U_10U_or_tmp & chn_inp_out_rsci_bawt & reg_chn_inp_out_rsci_ld_core_psct_cse
        & (chn_inp_in_rsci_d_mxwt[407:406]==2'b11) & and_dcpl_1957) | FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_3_mx0c1)
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_3 <= MUX_v_10_2_2((chn_inp_in_rsci_d_mxwt[405:396]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_3_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3_0 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_3_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_3_0 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_3 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_6_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3_1 <= chn_inp_in_rsci_d_mxwt[410];
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3_0 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3_0_mx0w0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_3_1 <= chn_inp_in_rsci_d_mxwt[282];
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_3_0 <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_1_lpi_1_dfm_3_0_mx0w0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_3 <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_1_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_3 <= 10'b0;
    end
    else if ( core_wen & ((and_dcpl_1980 & and_dcpl_1979 & (fsm_output[1])) | (and_dcpl_1984
        & and_dcpl_1979) | FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_3_mx0c1)
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_3 <= MUX_v_10_2_2((chn_inp_in_rsci_d_mxwt[421:412]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_4_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_2_lpi_1_dfm_3_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_3 <= 10'b0;
    end
    else if ( core_wen & ((and_dcpl_1993 & (chn_inp_in_rsci_d_mxwt[442]) & (chn_inp_in_rsci_d_mxwt[441])
        & (chn_inp_in_rsci_d_mxwt[438]) & and_dcpl_1989 & (fsm_output[1])) | (and_dcpl_1759
        & (chn_inp_in_rsci_d_mxwt[738]) & (chn_inp_in_rsci_d_mxwt[442]) & chn_inp_out_rsci_bawt
        & reg_chn_inp_out_rsci_ld_core_psct_cse & (chn_inp_in_rsci_d_mxwt[441]) &
        (chn_inp_in_rsci_d_mxwt[438]) & and_dcpl_1989) | FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_3_mx0c1)
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_3 <= MUX_v_10_2_2((chn_inp_in_rsci_d_mxwt[437:428]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_8_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_3_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3_0 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3 <= 4'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_3_1 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_3_0 <= 1'b0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_3 <= 4'b0;
    end
    else if ( FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_and_9_cse ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3_1 <= chn_inp_in_rsci_d_mxwt[442];
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3_0 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3_0_mx0w0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3 <= FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_3_1 <= chn_inp_in_rsci_d_mxwt[314];
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_3_0 <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_3_0_mx0w0;
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_3 <= FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_3_0_3_lpi_1_dfm_3_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_3 <= 10'b0;
    end
    else if ( core_wen & ((and_dcpl_1953 & and_dcpl_2011 & (fsm_output[1])) | (and_dcpl_2015
        & and_dcpl_2011) | FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_3_mx0c1)
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_3 <= MUX_v_10_2_2((chn_inp_in_rsci_d_mxwt[453:444]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_FpExpoWidthInc_5U_6U_10U_1U_1U_or_12_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_lpi_1_dfm_3_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2 <= 1'b0;
    end
    else if ( core_wen & (and_2497_rgt | and_dcpl_394 | and_2499_rgt | and_2501_rgt)
        & (mux_1845_nl) ) begin
      inp_lookup_1_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2 <= MUX1HOT_s_1_4_2((inp_lookup_1_IntShiftRight_69U_6U_32U_obits_fixed_or_nl),
          (inp_lookup_1_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_nl), inp_lookup_1_FpMul_6U_10U_2_else_2_if_acc_itm_6,
          inp_lookup_1_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs,
          {and_2497_rgt , and_dcpl_394 , and_2499_rgt , and_2501_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2 <= 1'b0;
    end
    else if ( core_wen & (and_2503_rgt | and_dcpl_402 | and_2505_rgt | and_2507_rgt)
        & (mux_1850_nl) ) begin
      inp_lookup_2_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2 <= MUX1HOT_s_1_4_2((inp_lookup_2_IntShiftRight_69U_6U_32U_obits_fixed_or_nl),
          (inp_lookup_2_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_nl), inp_lookup_2_FpMul_6U_10U_2_else_2_if_acc_itm_6,
          inp_lookup_2_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs,
          {and_2503_rgt , and_dcpl_402 , and_2505_rgt , and_2507_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2 <= 1'b0;
    end
    else if ( core_wen & (and_2509_rgt | and_dcpl_410 | and_2511_rgt | and_2513_rgt)
        & (mux_1855_nl) ) begin
      inp_lookup_3_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2 <= MUX1HOT_s_1_4_2((inp_lookup_3_IntShiftRight_69U_6U_32U_obits_fixed_or_nl),
          (inp_lookup_3_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_nl), inp_lookup_3_FpMul_6U_10U_2_else_2_if_acc_itm_6_1,
          inp_lookup_3_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs,
          {and_2509_rgt , and_dcpl_410 , and_2511_rgt , and_2513_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2 <= 1'b0;
    end
    else if ( core_wen & (and_2515_rgt | and_dcpl_416 | and_2517_rgt | and_2519_rgt)
        & (mux_1860_nl) ) begin
      inp_lookup_4_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2 <= MUX1HOT_s_1_4_2((inp_lookup_4_IntShiftRight_69U_6U_32U_obits_fixed_or_nl),
          (inp_lookup_4_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_nl), inp_lookup_4_FpMul_6U_10U_2_else_2_if_acc_itm_6,
          inp_lookup_4_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs,
          {and_2515_rgt , and_dcpl_416 , and_2517_rgt , and_2519_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_inp_lookup_1_else_else_a0_acc_reg <= 1'b0;
    end
    else if ( or_11_cse & core_wen & (~(nor_1798_cse | (chn_inp_in_rsci_d_mxwt[736])))
        ) begin
      reg_inp_lookup_1_else_else_a0_acc_reg <= inp_lookup_else_else_a0_mux1h_rgt[35];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_inp_lookup_1_else_else_a0_acc_1_reg <= 1'b0;
    end
    else if ( or_11_cse & core_wen & (~ (chn_inp_in_rsci_d_mxwt[736])) ) begin
      reg_inp_lookup_1_else_else_a0_acc_1_reg <= inp_lookup_else_else_a0_mux1h_rgt[34];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_1_else_else_b1_mul_itm_2 <= 51'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1861_nl) ) begin
      inp_lookup_1_else_else_b1_mul_itm_2 <= nl_inp_lookup_1_else_else_b1_mul_itm_2[50:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_inp_lookup_2_else_else_a0_acc_reg <= 1'b0;
    end
    else if ( or_11_cse & core_wen & (~(nor_1798_cse | (chn_inp_in_rsci_d_mxwt[737])))
        ) begin
      reg_inp_lookup_2_else_else_a0_acc_reg <= inp_lookup_else_else_a0_mux1h_1_rgt[35];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_inp_lookup_2_else_else_a0_acc_1_reg <= 1'b0;
    end
    else if ( or_11_cse & core_wen & (~ (chn_inp_in_rsci_d_mxwt[737])) ) begin
      reg_inp_lookup_2_else_else_a0_acc_1_reg <= inp_lookup_else_else_a0_mux1h_1_rgt[34];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_2_else_else_b1_mul_itm_2 <= 51'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1862_nl) ) begin
      inp_lookup_2_else_else_b1_mul_itm_2 <= nl_inp_lookup_2_else_else_b1_mul_itm_2[50:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_inp_lookup_3_else_else_a0_acc_reg <= 1'b0;
    end
    else if ( or_11_cse & core_wen & (~(nor_1798_cse | (chn_inp_in_rsci_d_mxwt[738])))
        ) begin
      reg_inp_lookup_3_else_else_a0_acc_reg <= inp_lookup_else_else_a0_mux1h_2_rgt[35];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_inp_lookup_3_else_else_a0_acc_1_reg <= 1'b0;
    end
    else if ( or_11_cse & core_wen & (~ (chn_inp_in_rsci_d_mxwt[738])) ) begin
      reg_inp_lookup_3_else_else_a0_acc_1_reg <= inp_lookup_else_else_a0_mux1h_2_rgt[34];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_3_else_else_b1_mul_itm_2 <= 51'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1863_nl) ) begin
      inp_lookup_3_else_else_b1_mul_itm_2 <= nl_inp_lookup_3_else_else_b1_mul_itm_2[50:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_inp_lookup_4_else_else_a0_acc_reg <= 1'b0;
    end
    else if ( or_11_cse & core_wen & (~(nor_1798_cse | (chn_inp_in_rsci_d_mxwt[739])))
        ) begin
      reg_inp_lookup_4_else_else_a0_acc_reg <= inp_lookup_else_else_a0_mux1h_3_rgt[35];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_inp_lookup_4_else_else_a0_acc_1_reg <= 1'b0;
    end
    else if ( or_11_cse & core_wen & (~ (chn_inp_in_rsci_d_mxwt[739])) ) begin
      reg_inp_lookup_4_else_else_a0_acc_1_reg <= inp_lookup_else_else_a0_mux1h_3_rgt[34];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      inp_lookup_4_else_else_b1_mul_itm_2 <= 51'b0;
    end
    else if ( core_wen & (~ and_dcpl_78) & (mux_1864_nl) ) begin
      inp_lookup_4_else_else_b1_mul_itm_2 <= nl_inp_lookup_4_else_else_b1_mul_itm_2[50:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_3 <= 10'b0;
    end
    else if ( core_wen & ((and_dcpl_1927 & and_dcpl_1993 & (fsm_output[1])) | (and_dcpl_1927
        & and_dcpl_2005) | FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_3_mx0c1)
        ) begin
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_3 <= MUX_v_10_2_2((chn_inp_in_rsci_d_mxwt[309:300]),
          FpExpoWidthInc_5U_6U_10U_1U_1U_2_FpExpoWidthInc_5U_6U_10U_1U_1U_2_or_8_mx0w1,
          FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_3_lpi_1_dfm_3_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMantRNE_36U_11U_1_else_ac_int_cctor_tmp <= 10'b0;
    end
    else if ( (mux_2130_nl) & or_11_cse & (~(and_dcpl_383 | (cfg_precision_rsci_d[0])))
        & (cfg_precision_rsci_d[1]) & chn_inp_in_rsci_bawt & (~ (chn_inp_in_rsci_d_mxwt[739]))
        & core_wen ) begin
      reg_FpMantRNE_36U_11U_1_else_ac_int_cctor_tmp <= FpMantRNE_36U_11U_1_else_ac_int_cctor_sva_mx0w0[10:1];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMantRNE_36U_11U_1_else_ac_int_cctor_4_tmp <= 10'b0;
    end
    else if ( (mux_2131_nl) & or_11_cse & (~ and_dcpl_313) & chn_inp_in_rsci_bawt
        & (cfg_precision_rsci_d==2'b10) & (~ (chn_inp_in_rsci_d_mxwt[738])) & core_wen
        ) begin
      reg_FpMantRNE_36U_11U_1_else_ac_int_cctor_4_tmp <= FpMantRNE_36U_11U_1_else_ac_int_cctor_4_sva_mx0w0[10:1];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMantRNE_36U_11U_1_else_ac_int_cctor_3_tmp <= 10'b0;
    end
    else if ( (mux_2132_nl) & or_11_cse & (~(and_dcpl_243 | (cfg_precision_rsci_d[0])))
        & (cfg_precision_rsci_d[1]) & chn_inp_in_rsci_bawt & (~ (chn_inp_in_rsci_d_mxwt[737]))
        & core_wen ) begin
      reg_FpMantRNE_36U_11U_1_else_ac_int_cctor_3_tmp <= FpMantRNE_36U_11U_1_else_ac_int_cctor_3_sva_mx0w0[10:1];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpMantRNE_36U_11U_1_else_ac_int_cctor_2_tmp <= 10'b0;
    end
    else if ( (mux_2133_nl) & or_11_cse & (~(and_dcpl_173 | (cfg_precision_rsci_d[0])))
        & (cfg_precision_rsci_d[1]) & chn_inp_in_rsci_bawt & (~ (chn_inp_in_rsci_d_mxwt[736]))
        & core_wen ) begin
      reg_FpMantRNE_36U_11U_1_else_ac_int_cctor_2_tmp <= FpMantRNE_36U_11U_1_else_ac_int_cctor_2_sva_mx0w0[10:1];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_8U_23U_o_expo_1_lpi_1_dfm_12_tmp <= 2'b0;
      reg_FpAdd_8U_23U_o_expo_1_lpi_1_dfm_12_tmp_1 <= 6'b0;
    end
    else if ( FpAdd_8U_23U_o_expo_and_14_ssc ) begin
      reg_FpAdd_8U_23U_o_expo_1_lpi_1_dfm_12_tmp <= reg_FpAdd_8U_23U_o_expo_1_lpi_1_dfm_11_reg;
      reg_FpAdd_8U_23U_o_expo_1_lpi_1_dfm_12_tmp_1 <= reg_FpAdd_8U_23U_o_expo_1_lpi_1_dfm_11_1_reg;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_8U_23U_o_expo_2_lpi_1_dfm_12_tmp <= 2'b0;
      reg_FpAdd_8U_23U_o_expo_2_lpi_1_dfm_12_tmp_1 <= 6'b0;
    end
    else if ( FpAdd_8U_23U_o_expo_and_13_ssc ) begin
      reg_FpAdd_8U_23U_o_expo_2_lpi_1_dfm_12_tmp <= reg_FpAdd_8U_23U_o_expo_2_lpi_1_dfm_11_reg;
      reg_FpAdd_8U_23U_o_expo_2_lpi_1_dfm_12_tmp_1 <= reg_FpAdd_8U_23U_o_expo_2_lpi_1_dfm_11_1_reg;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpAdd_8U_23U_o_expo_lpi_1_dfm_12_tmp <= 2'b0;
      reg_FpAdd_8U_23U_o_expo_lpi_1_dfm_12_tmp_1 <= 6'b0;
    end
    else if ( FpAdd_8U_23U_o_expo_and_12_ssc ) begin
      reg_FpAdd_8U_23U_o_expo_lpi_1_dfm_12_tmp <= reg_FpAdd_8U_23U_o_expo_lpi_1_dfm_11_reg;
      reg_FpAdd_8U_23U_o_expo_lpi_1_dfm_12_tmp_1 <= reg_FpAdd_8U_23U_o_expo_lpi_1_dfm_11_1_reg;
    end
  end
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_mux_5_nl = MUX_v_4_2_2(FpAdd_6U_10U_o_expo_1_lpi_1_dfm_7_3_0,
      4'b1110, IsInf_6U_23U_land_1_lpi_1_dfm_mx0w0);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_4_nl =
      MUX_v_4_2_2((FpExpoWidthInc_6U_8U_23U_0U_1U_mux_5_nl), 4'b1111, IsNaN_6U_23U_IsNaN_6U_23U_nor_tmp);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_20_nl =
      (FpAdd_6U_10U_o_expo_1_lpi_1_dfm_7_5_4[0]) | IsInf_6U_23U_land_1_lpi_1_dfm_mx1
      | IsNaN_6U_23U_land_1_lpi_1_dfm_mx2;
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_mux_18_nl = MUX_v_4_2_2(FpAdd_6U_10U_o_expo_2_lpi_1_dfm_7_3_0,
      4'b1110, IsInf_6U_23U_land_2_lpi_1_dfm_mx0w0);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_9_nl =
      MUX_v_4_2_2((FpExpoWidthInc_6U_8U_23U_0U_1U_mux_18_nl), 4'b1111, IsNaN_6U_23U_IsNaN_6U_23U_nor_1_tmp);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_21_nl =
      (FpAdd_6U_10U_o_expo_2_lpi_1_dfm_7_5_4[0]) | IsInf_6U_23U_land_2_lpi_1_dfm_mx1
      | IsNaN_6U_23U_land_2_lpi_1_dfm_mx2;
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_mux_31_nl = MUX_v_4_2_2(FpAdd_6U_10U_o_expo_3_lpi_1_dfm_7_3_0,
      4'b1110, IsInf_6U_23U_land_3_lpi_1_dfm_mx0w0);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_14_nl =
      MUX_v_4_2_2((FpExpoWidthInc_6U_8U_23U_0U_1U_mux_31_nl), 4'b1111, IsNaN_6U_23U_IsNaN_6U_23U_nor_2_tmp);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_22_nl =
      (FpAdd_6U_10U_o_expo_3_lpi_1_dfm_7_5_4[0]) | IsInf_6U_23U_land_3_lpi_1_dfm_mx1
      | IsNaN_6U_23U_land_3_lpi_1_dfm_mx1;
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_mux_44_nl = MUX_v_4_2_2(FpAdd_6U_10U_o_expo_lpi_1_dfm_7_3_0,
      4'b1110, IsInf_6U_23U_land_lpi_1_dfm_mx0w0);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_19_nl =
      MUX_v_4_2_2((FpExpoWidthInc_6U_8U_23U_0U_1U_mux_44_nl), 4'b1111, IsNaN_6U_23U_IsNaN_6U_23U_nor_3_tmp);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_23_nl =
      (FpAdd_6U_10U_o_expo_lpi_1_dfm_7_5_4[0]) | IsInf_6U_23U_land_lpi_1_dfm_mx1
      | IsNaN_6U_23U_land_lpi_1_dfm_mx1;
  assign nor_1802_nl = ~(inp_lookup_asn_110 | or_5836_tmp);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_4_nl =
      IsInf_6U_23U_land_1_lpi_1_dfm_mx1 & (~ IsNaN_6U_23U_land_1_lpi_1_dfm_mx2);
  assign inp_lookup_or_nl = ((~ IsNaN_6U_23U_3_land_1_lpi_1_dfm_10) & inp_lookup_and_8_m1c)
      | (IsNaN_6U_23U_3_land_1_lpi_1_dfm_10 & inp_lookup_and_8_m1c);
  assign inp_lookup_and_82_nl = inp_lookup_and_10_m1c & (~ and_3545_tmp);
  assign nl_inp_lookup_1_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl = conv_u2u_2_3({1'b1
      , (FpAdd_6U_10U_o_expo_1_lpi_1_dfm_7_5_4[1])}) + 3'b1;
  assign inp_lookup_1_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl = nl_inp_lookup_1_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl[2:0];
  assign IsZero_6U_23U_aelse_IsZero_6U_23U_or_3_nl = (FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_22_13_1_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_9_0_1_lpi_1_dfm!=10'b0000000000)
      | (FpAdd_6U_10U_o_expo_1_lpi_1_dfm_7_5_4!=2'b00) | (FpAdd_6U_10U_o_expo_1_lpi_1_dfm_7_3_0!=4'b0000);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_nl = MUX_v_3_2_2(3'b000,
      (inp_lookup_1_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl), (IsZero_6U_23U_aelse_IsZero_6U_23U_or_3_nl));
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_3_nl =
      (FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_nl) | ({{2{IsInf_6U_23U_land_1_lpi_1_dfm_mx0w0}},
      IsInf_6U_23U_land_1_lpi_1_dfm_mx0w0}) | ({{2{IsNaN_6U_23U_IsNaN_6U_23U_nor_tmp}},
      IsNaN_6U_23U_IsNaN_6U_23U_nor_tmp});
  assign nor_1803_nl = ~(inp_lookup_asn_126 | or_5838_tmp);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_9_nl =
      IsInf_6U_23U_land_2_lpi_1_dfm_mx1 & (~ IsNaN_6U_23U_land_2_lpi_1_dfm_mx2);
  assign inp_lookup_or_1_nl = ((~ IsNaN_6U_23U_3_land_2_lpi_1_dfm_10) & inp_lookup_and_28_m1c)
      | (IsNaN_6U_23U_3_land_2_lpi_1_dfm_10 & inp_lookup_and_28_m1c);
  assign inp_lookup_and_86_nl = inp_lookup_and_30_m1c & (~ and_3546_tmp);
  assign nl_inp_lookup_2_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl = conv_u2u_2_3({1'b1
      , (FpAdd_6U_10U_o_expo_2_lpi_1_dfm_7_5_4[1])}) + 3'b1;
  assign inp_lookup_2_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl = nl_inp_lookup_2_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl[2:0];
  assign IsZero_6U_23U_aelse_IsZero_6U_23U_or_2_nl = (FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_22_13_2_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_9_0_2_lpi_1_dfm!=10'b0000000000)
      | (FpAdd_6U_10U_o_expo_2_lpi_1_dfm_7_5_4!=2'b00) | (FpAdd_6U_10U_o_expo_2_lpi_1_dfm_7_3_0!=4'b0000);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_5_nl =
      MUX_v_3_2_2(3'b000, (inp_lookup_2_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl),
      (IsZero_6U_23U_aelse_IsZero_6U_23U_or_2_nl));
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_8_nl =
      (FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_5_nl) |
      ({{2{IsInf_6U_23U_land_2_lpi_1_dfm_mx0w0}}, IsInf_6U_23U_land_2_lpi_1_dfm_mx0w0})
      | ({{2{IsNaN_6U_23U_IsNaN_6U_23U_nor_1_tmp}}, IsNaN_6U_23U_IsNaN_6U_23U_nor_1_tmp});
  assign nor_1804_nl = ~(inp_lookup_asn_118 | or_5840_tmp);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_14_nl
      = IsInf_6U_23U_land_3_lpi_1_dfm_mx1 & (~ IsNaN_6U_23U_land_3_lpi_1_dfm_mx1);
  assign inp_lookup_or_2_nl = ((~ IsNaN_6U_23U_3_land_3_lpi_1_dfm_10) & inp_lookup_and_48_m1c)
      | (IsNaN_6U_23U_3_land_3_lpi_1_dfm_10 & inp_lookup_and_48_m1c);
  assign inp_lookup_and_90_nl = inp_lookup_and_50_m1c & (~ and_3547_tmp);
  assign nl_inp_lookup_3_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl = conv_u2u_2_3({1'b1
      , (FpAdd_6U_10U_o_expo_3_lpi_1_dfm_7_5_4[1])}) + 3'b1;
  assign inp_lookup_3_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl = nl_inp_lookup_3_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl[2:0];
  assign IsZero_6U_23U_aelse_IsZero_6U_23U_or_1_nl = (FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_22_13_3_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_9_0_3_lpi_1_dfm!=10'b0000000000)
      | (FpAdd_6U_10U_o_expo_3_lpi_1_dfm_7_5_4!=2'b00) | (FpAdd_6U_10U_o_expo_3_lpi_1_dfm_7_3_0!=4'b0000);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_10_nl
      = MUX_v_3_2_2(3'b000, (inp_lookup_3_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl),
      (IsZero_6U_23U_aelse_IsZero_6U_23U_or_1_nl));
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_13_nl =
      (FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_10_nl) |
      ({{2{IsInf_6U_23U_land_3_lpi_1_dfm_mx0w0}}, IsInf_6U_23U_land_3_lpi_1_dfm_mx0w0})
      | ({{2{IsNaN_6U_23U_IsNaN_6U_23U_nor_2_tmp}}, IsNaN_6U_23U_IsNaN_6U_23U_nor_2_tmp});
  assign nor_1805_nl = ~(inp_lookup_asn_102 | or_5842_tmp);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_19_nl
      = IsInf_6U_23U_land_lpi_1_dfm_mx1 & (~ IsNaN_6U_23U_land_lpi_1_dfm_mx1);
  assign inp_lookup_or_3_nl = ((~ IsNaN_6U_23U_3_land_lpi_1_dfm_10) & inp_lookup_and_68_m1c)
      | (IsNaN_6U_23U_3_land_lpi_1_dfm_10 & inp_lookup_and_68_m1c);
  assign inp_lookup_and_94_nl = inp_lookup_and_70_m1c & (~ and_3548_tmp);
  assign nl_inp_lookup_4_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl = conv_u2u_2_3({1'b1
      , (FpAdd_6U_10U_o_expo_lpi_1_dfm_7_5_4[1])}) + 3'b1;
  assign inp_lookup_4_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl = nl_inp_lookup_4_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl[2:0];
  assign IsZero_6U_23U_aelse_IsZero_6U_23U_or_nl = (FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_22_13_lpi_1_dfm!=10'b0000000000)
      | (FpMantWidthInc_6U_10U_23U_0U_1U_o_mant_9_0_lpi_1_dfm!=10'b0000000000) |
      (FpAdd_6U_10U_o_expo_lpi_1_dfm_7_5_4!=2'b00) | (FpAdd_6U_10U_o_expo_lpi_1_dfm_7_3_0!=4'b0000);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_15_nl
      = MUX_v_3_2_2(3'b000, (inp_lookup_4_FpExpoWidthInc_6U_8U_23U_0U_1U_else_acc_nl),
      (IsZero_6U_23U_aelse_IsZero_6U_23U_or_nl));
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_or_18_nl =
      (FpExpoWidthInc_6U_8U_23U_0U_1U_FpExpoWidthInc_6U_8U_23U_0U_1U_and_15_nl) |
      ({{2{IsInf_6U_23U_land_lpi_1_dfm_mx0w0}}, IsInf_6U_23U_land_lpi_1_dfm_mx0w0})
      | ({{2{IsNaN_6U_23U_IsNaN_6U_23U_nor_3_tmp}}, IsNaN_6U_23U_IsNaN_6U_23U_nor_3_tmp});
  assign inp_lookup_if_mux_600_nl = MUX_s_1_2_2((FpExpoWidthInc_6U_8U_23U_0U_1U_o_mant_9_0_1_lpi_1_dfm_2_mx0[0]),
      (IntSaturation_51U_32U_o_1_lpi_1_dfm_12_30_0_1[0]), inp_lookup_if_unequal_tmp_19);
  assign inp_lookup_if_mux_601_nl = MUX_s_1_2_2((FpExpoWidthInc_6U_8U_23U_0U_1U_o_mant_9_0_2_lpi_1_dfm_2_mx0[0]),
      (IntSaturation_51U_32U_o_2_lpi_1_dfm_12_30_0_1[0]), inp_lookup_if_unequal_tmp_19);
  assign inp_lookup_if_mux_602_nl = MUX_s_1_2_2((FpExpoWidthInc_6U_8U_23U_0U_1U_o_mant_9_0_3_lpi_1_dfm_2_mx0[0]),
      (IntSaturation_51U_32U_o_3_lpi_1_dfm_12_30_0_1[0]), inp_lookup_if_unequal_tmp_19);
  assign inp_lookup_if_mux_603_nl = MUX_s_1_2_2((FpExpoWidthInc_6U_8U_23U_0U_1U_o_mant_9_0_lpi_1_dfm_2_mx0[0]),
      (IntSaturation_51U_32U_o_lpi_1_dfm_12_30_0_1[0]), inp_lookup_if_unequal_tmp_19);
  assign inp_lookup_1_FpAdd_6U_10U_IsZero_6U_10U_2_nand_nl = ~(inp_lookup_1_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_2
      & inp_lookup_1_IsZero_6U_10U_5_IsZero_6U_10U_5_nor_2);
  assign IsZero_6U_10U_7_IsZero_6U_10U_7_and_nl = (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_3_mx1==10'b0000000000)
      & (~((chn_inp_in_rsci_d_mxwt[346]) | FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_3_0_mx0w0
      | (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_3_mx0w0!=4'b0000)));
  assign IsZero_6U_10U_5_IsZero_6U_10U_5_and_nl = inp_lookup_1_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_2
      & inp_lookup_1_IsZero_6U_10U_5_IsZero_6U_10U_5_nor_2;
  assign IsZero_6U_10U_1_IsZero_6U_10U_1_and_nl = (FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_1_lpi_1_dfm_3_mx1==10'b0000000000)
      & (~((chn_inp_in_rsci_d_mxwt[410]) | FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_3_0_mx0w0
      | (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_3_mx0w0!=4'b0000)));
  assign nor_1721_nl = ~((chn_inp_in_rsci_d_mxwt[736]) | (~ chn_inp_in_rsci_bawt)
      | (cfg_precision_rsci_d!=2'b10) | not_tmp_34);
  assign nor_1722_nl = ~((~ main_stage_v_1) | (chn_inp_in_crt_sva_1_739_395_1[341])
      | (~((inp_lookup_1_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_3!=35'b00000000000000000000000000000000000)))
      | (cfg_precision_1_sva_st_90!=2'b10));
  assign mux_80_nl = MUX_s_1_2_2((nor_1722_nl), (nor_1721_nl), or_11_cse);
  assign FpFractionToFloat_35U_6U_10U_1_if_else_else_FpFractionToFloat_35U_6U_10U_1_if_else_else_and_nl
      = MUX_v_10_2_2(10'b0000000000, (FpMantRNE_36U_11U_1_else_ac_int_cctor_2_sva_mx0w0[9:0]),
      inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_itm_5);
  assign FpFractionToFloat_35U_6U_10U_1_o_mant_and_nl = (~ and_dcpl_173) & FpFractionToFloat_35U_6U_10U_1_o_mant_1_lpi_1_dfm_6_mx0c1;
  assign FpFractionToFloat_35U_6U_10U_1_o_mant_and_10_nl = and_dcpl_173 & FpFractionToFloat_35U_6U_10U_1_o_mant_1_lpi_1_dfm_6_mx0c1;
  assign inp_lookup_2_IsZero_6U_10U_1_IsZero_6U_10U_1_nor_nl = ~((chn_inp_in_rsci_d_mxwt[426])
      | FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_3_0_mx0w0 | (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_3_mx0w0!=4'b0000));
  assign inp_lookup_2_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_nl = (chn_inp_in_rsci_d_mxwt[62:32]!=31'b0000000000000000000000000000000);
  assign IsZero_6U_10U_5_IsZero_6U_10U_5_and_1_nl = inp_lookup_2_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_mx0w0
      & inp_lookup_2_IsZero_6U_10U_5_IsZero_6U_10U_5_nor_mx0w1;
  assign nor_1717_nl = ~((chn_inp_in_rsci_d_mxwt[737]) | (~ chn_inp_in_rsci_bawt)
      | (cfg_precision_rsci_d!=2'b10) | not_tmp_45);
  assign nor_1718_nl = ~((~ main_stage_v_1) | (chn_inp_in_crt_sva_1_739_395_1[342])
      | (~((inp_lookup_2_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_3!=35'b00000000000000000000000000000000000)))
      | (cfg_precision_1_sva_st_90!=2'b10));
  assign mux_86_nl = MUX_s_1_2_2((nor_1718_nl), (nor_1717_nl), or_11_cse);
  assign inp_lookup_2_FpAdd_8U_23U_IsZero_8U_23U_1_or_nl = (chn_inp_in_rsci_d_mxwt[670:640]!=31'b0000000000000000000000000000000);
  assign IsZero_6U_10U_7_IsZero_6U_10U_7_and_1_nl = (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_3_mx1==10'b0000000000)
      & (~((chn_inp_in_rsci_d_mxwt[362]) | FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_2_lpi_1_dfm_3_0_mx0w0
      | (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_2_lpi_1_dfm_3_mx0w0!=4'b0000)));
  assign nand_nl = ~(main_stage_v_1 & (~ or_2010_cse));
  assign mux_92_nl = MUX_s_1_2_2((nand_nl), or_tmp_6, or_11_cse);
  assign FpFractionToFloat_35U_6U_10U_1_if_else_else_FpFractionToFloat_35U_6U_10U_1_if_else_else_and_1_nl
      = MUX_v_10_2_2(10'b0000000000, (FpMantRNE_36U_11U_1_else_ac_int_cctor_3_sva_mx0w0[9:0]),
      inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_itm_5);
  assign FpFractionToFloat_35U_6U_10U_1_o_mant_and_8_nl = (~ and_dcpl_243) & FpFractionToFloat_35U_6U_10U_1_o_mant_2_lpi_1_dfm_6_mx0c1;
  assign FpFractionToFloat_35U_6U_10U_1_o_mant_and_9_nl = and_dcpl_243 & FpFractionToFloat_35U_6U_10U_1_o_mant_2_lpi_1_dfm_6_mx0c1;
  assign inp_lookup_3_FpAdd_6U_10U_IsZero_6U_10U_2_nand_nl = ~(inp_lookup_3_IsZero_6U_10U_2_aif_IsZero_6U_10U_2_aelse_nor_2
      & inp_lookup_3_IsZero_6U_10U_5_IsZero_6U_10U_5_nor_2);
  assign IsZero_6U_10U_7_IsZero_6U_10U_7_and_2_nl = (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_3_lpi_1_dfm_3_mx1==10'b0000000000)
      & (~((chn_inp_in_rsci_d_mxwt[378]) | FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_3_lpi_1_dfm_3_0_mx0w0
      | (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_3_lpi_1_dfm_3_mx0w0!=4'b0000)));
  assign IsZero_6U_10U_5_IsZero_6U_10U_5_and_2_nl = inp_lookup_3_IsZero_6U_10U_2_aif_IsZero_6U_10U_2_aelse_nor_2
      & inp_lookup_3_IsZero_6U_10U_5_IsZero_6U_10U_5_nor_2;
  assign IsZero_6U_10U_1_IsZero_6U_10U_1_and_2_nl = (FpExpoWidthInc_5U_6U_10U_1U_1U_o_mant_3_lpi_1_dfm_3_mx1==10'b0000000000)
      & (~((chn_inp_in_rsci_d_mxwt[442]) | FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_3_0_mx0w0
      | (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_3_mx0w0!=4'b0000)));
  assign nor_1715_nl = ~((chn_inp_in_rsci_d_mxwt[738]) | (cfg_precision_rsci_d!=2'b10)
      | (~(chn_inp_in_rsci_bawt & or_79_cse)));
  assign nor_1716_nl = ~((~ main_stage_v_1) | (chn_inp_in_crt_sva_1_739_395_1[343])
      | (cfg_precision_1_sva_st_90[0]) | (~((cfg_precision_1_sva_st_90[1]) & or_82_cse)));
  assign mux_94_nl = MUX_s_1_2_2((nor_1716_nl), (nor_1715_nl), or_11_cse);
  assign FpFractionToFloat_35U_6U_10U_1_if_else_else_FpFractionToFloat_35U_6U_10U_1_if_else_else_and_2_nl
      = MUX_v_10_2_2(10'b0000000000, (FpMantRNE_36U_11U_1_else_ac_int_cctor_4_sva_mx0w0[9:0]),
      inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_itm_5);
  assign FpFractionToFloat_35U_6U_10U_1_o_mant_and_6_nl = (~ and_dcpl_313) & FpFractionToFloat_35U_6U_10U_1_o_mant_3_lpi_1_dfm_6_mx0c1;
  assign FpFractionToFloat_35U_6U_10U_1_o_mant_and_7_nl = and_dcpl_313 & FpFractionToFloat_35U_6U_10U_1_o_mant_3_lpi_1_dfm_6_mx0c1;
  assign nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_nl = ({1'b1 , (chn_inp_in_rsci_d_mxwt[598:576])})
      + conv_u2u_23_24(~ (chn_inp_in_rsci_d_mxwt[726:704])) + 24'b1;
  assign FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_nl = nl_FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_nl[23:0];
  assign nl_FpAdd_8U_23U_is_a_greater_acc_3_nl = ({1'b1 , (chn_inp_in_rsci_d_mxwt[734:727])})
      + conv_u2u_8_9(~ (chn_inp_in_rsci_d_mxwt[606:599])) + 9'b1;
  assign FpAdd_8U_23U_is_a_greater_acc_3_nl = nl_FpAdd_8U_23U_is_a_greater_acc_3_nl[8:0];
  assign FpAdd_8U_23U_is_a_greater_FpAdd_8U_23U_is_a_greater_or_3_nl = (~((readslicef_24_1_23((FpAdd_8U_23U_is_a_greater_oif_aelse_acc_3_nl)))
      | ((chn_inp_in_rsci_d_mxwt[606:599]) != (chn_inp_in_rsci_d_mxwt[734:727]))))
      | (readslicef_9_1_8((FpAdd_8U_23U_is_a_greater_acc_3_nl)));
  assign inp_lookup_4_FpAdd_8U_23U_1_IsZero_8U_23U_2_or_nl = (chn_inp_in_rsci_d_mxwt[126:96]!=31'b0000000000000000000000000000000);
  assign IsZero_6U_10U_5_IsZero_6U_10U_5_and_3_nl = inp_lookup_4_IsZero_6U_10U_5_aif_IsZero_6U_10U_5_aelse_nor_mx0w0
      & inp_lookup_4_IsZero_6U_10U_5_IsZero_6U_10U_5_nor_mx0w1;
  assign nor_1760_nl = ~((chn_inp_in_rsci_d_mxwt[739]) | (~ chn_inp_in_rsci_bawt)
      | (cfg_precision_rsci_d!=2'b10) | not_tmp_69);
  assign nor_1761_nl = ~((chn_inp_in_crt_sva_1_739_395_1[344]) | nor_1713_cse | (~
      main_stage_v_1) | (cfg_precision_1_sva_st_90!=2'b10));
  assign mux_99_nl = MUX_s_1_2_2((nor_1761_nl), (nor_1760_nl), or_11_cse);
  assign inp_lookup_4_FpAdd_8U_23U_IsZero_8U_23U_1_or_nl = (chn_inp_in_rsci_d_mxwt[734:704]!=31'b0000000000000000000000000000000);
  assign IsZero_6U_10U_7_IsZero_6U_10U_7_and_3_nl = (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_3_mx1==10'b0000000000)
      & (~((chn_inp_in_rsci_d_mxwt[394]) | FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_3_0_mx0w0
      | (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_3_mx0w0!=4'b0000)));
  assign nand_2_nl = ~(main_stage_v_1 & nor_1336_cse_1);
  assign mux_104_nl = MUX_s_1_2_2(or_tmp_8, (nand_2_nl), chn_inp_in_crt_sva_1_739_395_1[344]);
  assign mux_105_nl = MUX_s_1_2_2((mux_104_nl), or_tmp_6, or_11_cse);
  assign FpFractionToFloat_35U_6U_10U_1_if_else_else_FpFractionToFloat_35U_6U_10U_1_if_else_else_and_3_nl
      = MUX_v_10_2_2(10'b0000000000, (FpMantRNE_36U_11U_1_else_ac_int_cctor_sva_mx0w0[9:0]),
      inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_else_else_if_acc_itm_5);
  assign FpFractionToFloat_35U_6U_10U_1_o_mant_and_4_nl = (~ and_dcpl_383) & FpFractionToFloat_35U_6U_10U_1_o_mant_lpi_1_dfm_6_mx0c1;
  assign FpFractionToFloat_35U_6U_10U_1_o_mant_and_5_nl = and_dcpl_383 & FpFractionToFloat_35U_6U_10U_1_o_mant_lpi_1_dfm_6_mx0c1;
  assign FpFractionToFloat_35U_6U_10U_if_else_else_FpFractionToFloat_35U_6U_10U_if_else_else_and_nl
      = MUX_v_10_2_2(10'b0000000000, (FpMantRNE_36U_11U_else_ac_int_cctor_2_sva[9:0]),
      inp_lookup_1_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_itm_5_1);
  assign nor_1707_nl = ~((cfg_precision_1_sva_st_90!=2'b10) | (chn_inp_in_crt_sva_1_739_395_1[341])
      | (~(main_stage_v_1 & IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_13 & ((inp_lookup_1_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_3!=35'b00000000000000000000000000000000000))
      & (inp_lookup_1_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_itm_5_1 |
      inp_lookup_1_FpMantRNE_36U_11U_else_and_tmp))));
  assign nor_1708_nl = ~((~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[0])
      | (cfg_precision_1_sva_st_91!=2'b10) | FpFractionToFloat_35U_6U_10U_is_zero_1_lpi_1_dfm_5
      | (~(IsNaN_8U_23U_land_1_lpi_1_dfm_st_4 & ((inp_lookup_1_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_4!=35'b00000000000000000000000000000000000)))));
  assign mux_111_nl = MUX_s_1_2_2((nor_1708_nl), (nor_1707_nl), or_11_cse);
  assign or_156_nl = (inp_lookup_1_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_3!=35'b00000000000000000000000000000000000)
      | (chn_inp_in_crt_sva_1_739_395_1[341]);
  assign mux_112_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_1_739_395_1[341]), (or_156_nl),
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_13);
  assign nor_1703_nl = ~((~ main_stage_v_1) | (cfg_precision_1_sva_st_90[0]) | (~((cfg_precision_1_sva_st_90[1])
      & (mux_112_nl))));
  assign nor_1704_nl = ~((~((inp_lookup_1_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_4!=35'b00000000000000000000000000000000000)
      | (chn_inp_in_crt_sva_2_739_736_1[0]))) | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10));
  assign mux_113_nl = MUX_s_1_2_2(and_3393_cse, (nor_1704_nl), IsNaN_8U_23U_land_1_lpi_1_dfm_st_4);
  assign mux_114_nl = MUX_s_1_2_2((mux_113_nl), (nor_1703_nl), or_11_cse);
  assign IsNaN_6U_10U_6_IsNaN_6U_10U_6_nor_nl = ~(IsNaN_6U_10U_6_nor_tmp | (~(FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_3_5_mx0w0
      & (FpFractionToFloat_35U_6U_10U_1_o_expo_1_lpi_1_dfm_3_4_0_mx0w0==5'b11111))));
  assign nor_1893_nl = ~(inp_lookup_1_FpMul_6U_10U_2_else_2_if_acc_itm_6 | (~ or_tmp_4611));
  assign mux_2043_nl = MUX_s_1_2_2((nor_1893_nl), or_tmp_4611, or_5873_cse);
  assign nor_1894_nl = ~(inp_lookup_1_FpMul_6U_10U_2_else_2_if_acc_itm_6 | (~ or_tmp_4615));
  assign mux_2044_nl = MUX_s_1_2_2((nor_1894_nl), or_tmp_4615, or_5873_cse);
  assign mux_2045_nl = MUX_s_1_2_2((mux_2044_nl), (mux_2043_nl), FpFractionToFloat_35U_6U_10U_1_o_mant_1_lpi_1_dfm_6[9]);
  assign and_4147_nl = (~(FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_6_1_1
      & FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_1_lpi_1_dfm_6_0_1 & (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_1_lpi_1_dfm_9==4'b1111)))
      & or_tmp_4620;
  assign and_4148_nl = ((FpFractionToFloat_35U_6U_10U_1_o_mant_1_lpi_1_dfm_6!=10'b0000000000))
      & (FpFractionToFloat_35U_6U_10U_1_mux_tmp[4:3]==2'b11) & (IntLeadZero_35U_1_leading_sign_35_0_rtn_1_sva_2[5])
      & inp_lookup_1_FpMantRNE_36U_11U_1_else_and_svs_2 & FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_st_2
      & (FpFractionToFloat_35U_6U_10U_1_mux_tmp[2:0]==3'b111);
  assign mux_2046_nl = MUX_s_1_2_2((and_4147_nl), or_tmp_4620, and_4148_nl);
  assign mux_2047_nl = MUX_s_1_2_2(or_tmp_4620, (mux_2046_nl), or_5882_cse);
  assign nl_inp_lookup_1_FpFractionToFloat_35U_6U_10U_if_else_else_else_acc_nl =
      (~ (IntLeadZero_35U_leading_sign_35_0_rtn_1_sva_2[4:0])) + 5'b11111;
  assign inp_lookup_1_FpFractionToFloat_35U_6U_10U_if_else_else_else_acc_nl = nl_inp_lookup_1_FpFractionToFloat_35U_6U_10U_if_else_else_else_acc_nl[4:0];
  assign FpFractionToFloat_35U_6U_10U_if_else_mux_nl = MUX_v_5_2_2((inp_lookup_1_FpFractionToFloat_35U_6U_10U_if_else_else_else_acc_nl),
      (~ (IntLeadZero_35U_leading_sign_35_0_rtn_1_sva_2[4:0])), inp_lookup_1_FpMantRNE_36U_11U_else_and_tmp);
  assign FpFractionToFloat_35U_6U_10U_nor_nl = ~(MUX_v_5_2_2((FpFractionToFloat_35U_6U_10U_if_else_mux_nl),
      5'b11111, FpFractionToFloat_35U_6U_10U_is_zero_1_lpi_1_dfm_mx0w0));
  assign or_205_nl = (~ main_stage_v_1) | (chn_inp_in_crt_sva_1_739_395_1[341]) |
      (cfg_precision_1_sva_st_90[0]) | not_tmp_101;
  assign mux_126_nl = MUX_s_1_2_2(or_5800_cse, (or_205_nl), or_11_cse);
  assign or_208_nl = nor_1896_cse | (~ main_stage_v_1) | (chn_inp_in_crt_sva_1_739_395_1[341])
      | (cfg_precision_1_sva_st_90[0]) | not_tmp_101;
  assign mux_127_nl = MUX_s_1_2_2((or_208_nl), (mux_126_nl), IsNaN_8U_23U_land_1_lpi_1_dfm_st_4);
  assign FpFractionToFloat_35U_6U_10U_if_else_else_FpFractionToFloat_35U_6U_10U_if_else_else_and_1_nl
      = MUX_v_10_2_2(10'b0000000000, (FpMantRNE_36U_11U_else_ac_int_cctor_3_sva[9:0]),
      inp_lookup_2_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_itm_5_1);
  assign nor_1690_nl = ~((cfg_precision_1_sva_st_90!=2'b10) | (chn_inp_in_crt_sva_1_739_395_1[342])
      | (~(main_stage_v_1 & IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_13 & ((inp_lookup_2_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_3!=35'b00000000000000000000000000000000000))
      & (inp_lookup_2_FpMantRNE_36U_11U_else_and_tmp | inp_lookup_2_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_itm_5_1))));
  assign nor_1691_nl = ~((~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[1])
      | (cfg_precision_1_sva_st_91!=2'b10) | FpFractionToFloat_35U_6U_10U_is_zero_2_lpi_1_dfm_5
      | (~(IsNaN_8U_23U_land_2_lpi_1_dfm_st_4 & ((inp_lookup_2_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_4!=35'b00000000000000000000000000000000000)))));
  assign mux_134_nl = MUX_s_1_2_2((nor_1691_nl), (nor_1690_nl), or_11_cse);
  assign or_226_nl = (inp_lookup_2_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_3!=35'b00000000000000000000000000000000000)
      | (chn_inp_in_crt_sva_1_739_395_1[342]);
  assign mux_135_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_1_739_395_1[342]), (or_226_nl),
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_13);
  assign nor_1686_nl = ~((~ main_stage_v_1) | (cfg_precision_1_sva_st_90[0]) | (~((cfg_precision_1_sva_st_90[1])
      & (mux_135_nl))));
  assign nor_1687_nl = ~((~((inp_lookup_2_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_4!=35'b00000000000000000000000000000000000)
      | (chn_inp_in_crt_sva_2_739_736_1[1]))) | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10));
  assign mux_136_nl = MUX_s_1_2_2(and_3391_cse, (nor_1687_nl), IsNaN_8U_23U_land_2_lpi_1_dfm_st_4);
  assign mux_137_nl = MUX_s_1_2_2((mux_136_nl), (nor_1686_nl), or_11_cse);
  assign IsZero_6U_10U_1_IsZero_6U_10U_1_and_1_nl = inp_lookup_2_IsZero_6U_10U_1_aif_IsZero_6U_10U_1_aelse_nor_itm_2
      & FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_2_lpi_1_dfm_6_0_1;
  assign IsNaN_6U_10U_6_IsNaN_6U_10U_6_nor_1_nl = ~(IsNaN_6U_10U_6_nor_1_tmp | (~(FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_3_5_mx0w0
      & (FpFractionToFloat_35U_6U_10U_1_o_expo_2_lpi_1_dfm_3_4_0_mx0w0==5'b11111))));
  assign nor_1889_nl = ~(inp_lookup_2_FpMul_6U_10U_2_else_2_if_acc_itm_6 | (~ or_tmp_4625));
  assign mux_2048_nl = MUX_s_1_2_2((nor_1889_nl), or_tmp_4625, or_5890_cse);
  assign nor_1890_nl = ~((~(inp_lookup_2_FpMul_6U_10U_2_oelse_1_acc_itm_7 | IsZero_6U_10U_7_IsZero_6U_10U_7_and_1_itm_2
      | IsZero_6U_10U_6_IsZero_6U_10U_6_nor_1_tmp | (~ inp_lookup_2_FpMul_6U_10U_2_else_2_if_acc_itm_6)))
      | nor_tmp_708);
  assign and_4146_nl = (FpFractionToFloat_35U_6U_10U_1_mux_40_tmp==5'b11111) & (IntLeadZero_35U_1_leading_sign_35_0_rtn_2_sva_2[5])
      & inp_lookup_2_FpMantRNE_36U_11U_1_else_and_svs_2 & FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_st_2;
  assign mux_2049_nl = MUX_s_1_2_2((nor_1890_nl), (mux_2048_nl), and_4146_nl);
  assign mux_2050_nl = MUX_s_1_2_2(or_5896_cse, (mux_2049_nl), or_5889_cse);
  assign and_3610_nl = ((FpFractionToFloat_35U_6U_10U_1_o_mant_2_lpi_1_dfm_6!=10'b0000000000))
      & (FpFractionToFloat_35U_6U_10U_1_mux_40_tmp==5'b11111) & (IntLeadZero_35U_1_leading_sign_35_0_rtn_2_sva_2[5])
      & inp_lookup_2_FpMantRNE_36U_11U_1_else_and_svs_2 & FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_st_2
      & or_5896_cse;
  assign mux_2051_nl = MUX_s_1_2_2(or_5896_cse, (and_3610_nl), and_4145_cse);
  assign nl_inp_lookup_2_FpFractionToFloat_35U_6U_10U_if_else_else_else_acc_nl =
      (~ (IntLeadZero_35U_leading_sign_35_0_rtn_2_sva_2[4:0])) + 5'b11111;
  assign inp_lookup_2_FpFractionToFloat_35U_6U_10U_if_else_else_else_acc_nl = nl_inp_lookup_2_FpFractionToFloat_35U_6U_10U_if_else_else_else_acc_nl[4:0];
  assign FpFractionToFloat_35U_6U_10U_if_else_mux_16_nl = MUX_v_5_2_2((inp_lookup_2_FpFractionToFloat_35U_6U_10U_if_else_else_else_acc_nl),
      (~ (IntLeadZero_35U_leading_sign_35_0_rtn_2_sva_2[4:0])), inp_lookup_2_FpMantRNE_36U_11U_else_and_tmp);
  assign FpFractionToFloat_35U_6U_10U_nor_1_nl = ~(MUX_v_5_2_2((FpFractionToFloat_35U_6U_10U_if_else_mux_16_nl),
      5'b11111, FpFractionToFloat_35U_6U_10U_is_zero_2_lpi_1_dfm_mx0w0));
  assign or_269_nl = (~ main_stage_v_1) | (chn_inp_in_crt_sva_1_739_395_1[342]) |
      (cfg_precision_1_sva_st_90[0]) | not_tmp_126;
  assign mux_148_nl = MUX_s_1_2_2(or_tmp_234, (or_269_nl), or_11_cse);
  assign or_272_nl = nor_1896_cse | (~ main_stage_v_1) | (chn_inp_in_crt_sva_1_739_395_1[342])
      | (cfg_precision_1_sva_st_90[0]) | not_tmp_126;
  assign mux_149_nl = MUX_s_1_2_2((or_272_nl), (mux_148_nl), IsNaN_8U_23U_land_2_lpi_1_dfm_st_4);
  assign FpFractionToFloat_35U_6U_10U_if_else_else_FpFractionToFloat_35U_6U_10U_if_else_else_and_2_nl
      = MUX_v_10_2_2(10'b0000000000, (FpMantRNE_36U_11U_else_ac_int_cctor_4_sva[9:0]),
      inp_lookup_3_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_itm_5_1);
  assign nor_1671_nl = ~((cfg_precision_1_sva_st_90!=2'b10) | (chn_inp_in_crt_sva_1_739_395_1[343])
      | (~(main_stage_v_1 & IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_13 & or_82_cse & (inp_lookup_3_FpMantRNE_36U_11U_else_and_tmp
      | inp_lookup_3_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_itm_5_1))));
  assign nor_1672_nl = ~((~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[2])
      | (cfg_precision_1_sva_st_91!=2'b10) | FpFractionToFloat_35U_6U_10U_is_zero_3_lpi_1_dfm_5
      | (~(IsNaN_8U_23U_land_3_lpi_1_dfm_st_4 & ((inp_lookup_3_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_4!=35'b00000000000000000000000000000000000)))));
  assign mux_156_nl = MUX_s_1_2_2((nor_1672_nl), (nor_1671_nl), or_11_cse);
  assign nor_1665_nl = ~((~((inp_lookup_3_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_3!=35'b00000000000000000000000000000000000)
      | (chn_inp_in_crt_sva_1_739_395_1[343]))) | (~ main_stage_v_1) | (cfg_precision_1_sva_st_90!=2'b10));
  assign mux_157_nl = MUX_s_1_2_2(and_3389_cse, (nor_1665_nl), IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_13);
  assign nor_1668_nl = ~((~((inp_lookup_3_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_4!=35'b00000000000000000000000000000000000)
      | (chn_inp_in_crt_sva_2_739_736_1[2]))) | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10));
  assign mux_158_nl = MUX_s_1_2_2(and_3401_cse, (nor_1668_nl), IsNaN_8U_23U_land_3_lpi_1_dfm_st_4);
  assign mux_159_nl = MUX_s_1_2_2((mux_158_nl), (mux_157_nl), or_11_cse);
  assign IsNaN_6U_10U_6_IsNaN_6U_10U_6_nor_2_nl = ~(IsNaN_6U_10U_6_nor_2_tmp | (~(FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_3_5_mx0w0
      & (FpFractionToFloat_35U_6U_10U_1_o_expo_3_lpi_1_dfm_3_4_0_mx0w0==5'b11111))));
  assign nl_inp_lookup_3_FpFractionToFloat_35U_6U_10U_if_else_else_else_acc_nl =
      (~ (IntLeadZero_35U_leading_sign_35_0_rtn_3_sva_2[4:0])) + 5'b11111;
  assign inp_lookup_3_FpFractionToFloat_35U_6U_10U_if_else_else_else_acc_nl = nl_inp_lookup_3_FpFractionToFloat_35U_6U_10U_if_else_else_else_acc_nl[4:0];
  assign FpFractionToFloat_35U_6U_10U_if_else_mux_17_nl = MUX_v_5_2_2((inp_lookup_3_FpFractionToFloat_35U_6U_10U_if_else_else_else_acc_nl),
      (~ (IntLeadZero_35U_leading_sign_35_0_rtn_3_sva_2[4:0])), inp_lookup_3_FpMantRNE_36U_11U_else_and_tmp);
  assign FpFractionToFloat_35U_6U_10U_nor_2_nl = ~(MUX_v_5_2_2((FpFractionToFloat_35U_6U_10U_if_else_mux_17_nl),
      5'b11111, FpFractionToFloat_35U_6U_10U_is_zero_3_lpi_1_dfm_mx0w0));
  assign or_339_nl = (chn_inp_in_crt_sva_1_739_395_1[343]) | (~ main_stage_v_1) |
      (cfg_precision_1_sva_st_90[0]) | not_tmp_152;
  assign mux_168_nl = MUX_s_1_2_2(or_tmp_306, (or_339_nl), or_11_cse);
  assign or_342_nl = nor_1896_cse | (chn_inp_in_crt_sva_1_739_395_1[343]) | (~ main_stage_v_1)
      | (cfg_precision_1_sva_st_90[0]) | not_tmp_152;
  assign mux_169_nl = MUX_s_1_2_2((or_342_nl), (mux_168_nl), IsNaN_8U_23U_land_3_lpi_1_dfm_st_4);
  assign FpFractionToFloat_35U_6U_10U_if_else_else_FpFractionToFloat_35U_6U_10U_if_else_else_and_3_nl
      = MUX_v_10_2_2(10'b0000000000, (FpMantRNE_36U_11U_else_ac_int_cctor_sva[9:0]),
      inp_lookup_4_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_itm_5_1);
  assign nor_1656_nl = ~(nor_1713_cse | (chn_inp_in_crt_sva_1_739_395_1[344]) | (~
      main_stage_v_1) | (~ FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2) | (cfg_precision_1_sva_st_90[0])
      | (~((cfg_precision_1_sva_st_90[1]) & (inp_lookup_4_FpMantRNE_36U_11U_else_and_tmp
      | inp_lookup_4_FpFractionToFloat_35U_6U_10U_if_else_else_if_acc_itm_5_1))));
  assign nor_1658_nl = ~(FpFractionToFloat_35U_6U_10U_is_zero_lpi_1_dfm_5 | (~ main_stage_v_2)
      | (~ IsNaN_8U_23U_land_lpi_1_dfm_st_4) | (chn_inp_in_crt_sva_2_739_736_1[3])
      | (cfg_precision_1_sva_st_91[0]) | (~((cfg_precision_1_sva_st_91[1]) & or_356_cse)));
  assign mux_175_nl = MUX_s_1_2_2((nor_1658_nl), (nor_1656_nl), or_11_cse);
  assign or_360_nl = (inp_lookup_4_chn_inp_in_fraction_slc_chn_inp_in_crt_267_128_2_itm_3!=35'b00000000000000000000000000000000000)
      | (chn_inp_in_crt_sva_1_739_395_1[344]);
  assign mux_176_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_1_739_395_1[344]), (or_360_nl),
      FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2);
  assign nor_1654_nl = ~((~ main_stage_v_1) | (cfg_precision_1_sva_st_90[0]) | (~((cfg_precision_1_sva_st_90[1])
      & (mux_176_nl))));
  assign nor_1655_nl = ~((~ main_stage_v_2) | (cfg_precision_1_sva_st_91[0]) | (~((cfg_precision_1_sva_st_91[1])
      & ((chn_inp_in_crt_sva_2_739_736_1[3]) | (or_356_cse & IsNaN_8U_23U_land_lpi_1_dfm_st_4)))));
  assign mux_177_nl = MUX_s_1_2_2((nor_1655_nl), (nor_1654_nl), or_11_cse);
  assign IsZero_6U_10U_1_IsZero_6U_10U_1_and_3_nl = inp_lookup_4_IsZero_6U_10U_1_aif_IsZero_6U_10U_1_aelse_nor_itm_2
      & FpAdd_8U_23U_o_sign_lpi_1_dfm_1;
  assign IsNaN_6U_10U_6_IsNaN_6U_10U_6_nor_3_nl = ~(IsNaN_6U_10U_6_nor_3_tmp | (~(FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_3_5_mx0w0
      & (FpFractionToFloat_35U_6U_10U_1_o_expo_lpi_1_dfm_3_4_0_mx0w0==5'b11111))));
  assign and_4143_nl = (~(FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_6_1_1
      & FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_5_4_lpi_1_dfm_6_0_1 & (FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_expo_3_0_lpi_1_dfm_9==4'b1111)))
      & or_tmp_4637;
  assign and_4144_nl = or_6160_cse & (FpFractionToFloat_35U_6U_10U_1_mux_42_tmp==5'b11111)
      & (IntLeadZero_35U_1_leading_sign_35_0_rtn_sva_2[5]) & inp_lookup_4_FpMantRNE_36U_11U_1_else_and_svs_2
      & FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2;
  assign mux_2052_nl = MUX_s_1_2_2((and_4143_nl), or_tmp_4637, and_4144_nl);
  assign mux_2053_nl = MUX_s_1_2_2(or_tmp_4637, (mux_2052_nl), or_5904_cse);
  assign and_3622_nl = or_6160_cse & (FpFractionToFloat_35U_6U_10U_1_mux_42_tmp==5'b11111)
      & (IntLeadZero_35U_1_leading_sign_35_0_rtn_sva_2[5]) & inp_lookup_4_FpMantRNE_36U_11U_1_else_and_svs_2
      & FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2 & or_tmp_4637;
  assign mux_2054_nl = MUX_s_1_2_2(or_tmp_4637, (and_3622_nl), and_3361_cse_1);
  assign nl_inp_lookup_4_FpFractionToFloat_35U_6U_10U_if_else_else_else_acc_nl =
      (~ (IntLeadZero_35U_leading_sign_35_0_rtn_sva_2[4:0])) + 5'b11111;
  assign inp_lookup_4_FpFractionToFloat_35U_6U_10U_if_else_else_else_acc_nl = nl_inp_lookup_4_FpFractionToFloat_35U_6U_10U_if_else_else_else_acc_nl[4:0];
  assign FpFractionToFloat_35U_6U_10U_if_else_mux_18_nl = MUX_v_5_2_2((inp_lookup_4_FpFractionToFloat_35U_6U_10U_if_else_else_else_acc_nl),
      (~ (IntLeadZero_35U_leading_sign_35_0_rtn_sva_2[4:0])), inp_lookup_4_FpMantRNE_36U_11U_else_and_tmp);
  assign FpFractionToFloat_35U_6U_10U_nor_3_nl = ~(MUX_v_5_2_2((FpFractionToFloat_35U_6U_10U_if_else_mux_18_nl),
      5'b11111, FpFractionToFloat_35U_6U_10U_is_zero_lpi_1_dfm_mx0w0));
  assign nor_1644_nl = ~((chn_inp_in_crt_sva_1_739_395_1[344]) | (~ main_stage_v_1)
      | (~ FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2) | (cfg_precision_1_sva_st_90!=2'b10));
  assign nor_1645_nl = ~((~ main_stage_v_2) | (~ IsNaN_8U_23U_land_lpi_1_dfm_st_4)
      | (chn_inp_in_crt_sva_2_739_736_1[3]) | (cfg_precision_1_sva_st_91!=2'b10));
  assign mux_187_nl = MUX_s_1_2_2((nor_1645_nl), (nor_1644_nl), or_11_cse);
  assign nor_1641_nl = ~((~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ main_stage_v_3) | (~ (chn_inp_in_crt_sva_3_739_736_1[0])) | (cfg_precision_1_sva_st_80!=2'b10)
      | (FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_3_49_1_1[48]) | FpMul_6U_10U_1_lor_6_lpi_1_dfm_5
      | inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4);
  assign nor_1642_nl = ~((z_out[49]) | (~ main_stage_v_2) | (~ (chn_inp_in_crt_sva_2_739_736_1[0]))
      | (cfg_precision_1_sva_st_91!=2'b10));
  assign nor_1643_nl = ~((~ main_stage_v_3) | (~ (chn_inp_in_crt_sva_3_739_736_1[0]))
      | (cfg_precision_1_sva_st_80!=2'b10) | (FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_3_49_1_1[48])
      | FpMul_6U_10U_1_lor_6_lpi_1_dfm_5 | inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4);
  assign mux_188_nl = MUX_s_1_2_2((nor_1643_nl), (nor_1642_nl), or_11_cse);
  assign mux_189_nl = MUX_s_1_2_2((mux_188_nl), (nor_1641_nl), FpNormalize_8U_49U_if_FpNormalize_8U_49U_if_nand_tmp);
  assign mux_1870_nl = MUX_s_1_2_2(nand_772_cse, or_4340_cse, main_stage_v_3);
  assign FpAdd_8U_23U_o_mant_not_nl = ~ (fsm_output[0]);
  assign and_3421_nl = MUX_v_23_2_2(23'b00000000000000000000000, FpAdd_8U_23U_FpAdd_8U_23U_or_4_itm,
      (FpAdd_8U_23U_o_mant_not_nl));
  assign and_894_nl = and_dcpl_423 & (chn_inp_in_crt_sva_2_739_736_1[0]) & and_dcpl_419
      & (fsm_output[1]);
  assign mux_2210_nl = MUX_s_1_2_2(mux_tmp, or_tmp_4811, nor_1961_cse);
  assign nor_1977_nl = ~((cfg_precision_1_sva_st_90[1]) | (~ mux_tmp));
  assign mux_2211_nl = MUX_s_1_2_2((nor_1977_nl), mux_tmp, or_6241_cse);
  assign and_4228_nl = nand_602_cse_1 & mux_tmp;
  assign mux_2212_nl = MUX_s_1_2_2((and_4228_nl), (mux_2211_nl), main_stage_v_1);
  assign mux_2213_nl = MUX_s_1_2_2((mux_2212_nl), (mux_2210_nl), main_stage_v_2);
  assign mux_2214_nl = MUX_s_1_2_2((fsm_output[0]), or_tmp_4811, nor_1961_cse);
  assign mux_2215_nl = MUX_s_1_2_2(not_tmp_3015, (fsm_output[0]), or_6241_cse);
  assign and_4237_nl = nand_602_cse_1 & (fsm_output[0]);
  assign mux_2216_nl = MUX_s_1_2_2((and_4237_nl), (mux_2215_nl), main_stage_v_1);
  assign mux_2217_nl = MUX_s_1_2_2((mux_2216_nl), (mux_2214_nl), main_stage_v_2);
  assign mux_2218_nl = MUX_s_1_2_2((mux_2217_nl), (mux_2213_nl), main_stage_v_3);
  assign and_4229_nl = (fsm_output[0]) & or_4340_cse;
  assign or_6247_nl = (~ (chn_inp_in_crt_sva_2_739_736_1[0])) | (cfg_precision_1_sva_st_91[0]);
  assign mux_2219_nl = MUX_s_1_2_2(nor_1978_cse, (fsm_output[0]), or_6247_nl);
  assign or_6249_nl = (~ main_stage_v_1) | (~ (chn_inp_in_crt_sva_1_739_395_1[341]))
      | (cfg_precision_1_sva_st_90[0]);
  assign mux_2220_nl = MUX_s_1_2_2(not_tmp_3015, (fsm_output[0]), or_6249_nl);
  assign mux_2221_nl = MUX_s_1_2_2((mux_2220_nl), (mux_2219_nl), main_stage_v_2);
  assign mux_2222_nl = MUX_s_1_2_2((mux_2221_nl), (and_4229_nl), main_stage_v_3);
  assign mux_2223_nl = MUX_s_1_2_2((mux_2222_nl), (mux_2218_nl), or_11_cse);
  assign or_6250_nl = (~ main_stage_v_3) | IsNaN_6U_10U_6_land_1_lpi_1_dfm_5 | IsNaN_6U_10U_7_land_1_lpi_1_dfm_6;
  assign mux_2224_nl = MUX_s_1_2_2(or_tmp_4815, (fsm_output[0]), or_6250_nl);
  assign mux_2225_nl = MUX_s_1_2_2((mux_2224_nl), (mux_2223_nl), fsm_output[1]);
  assign nand_684_nl = ~(main_stage_v_3 & (chn_inp_in_crt_sva_3_739_736_1[0]) & (cfg_precision_1_sva_st_80==2'b10));
  assign mux_196_nl = MUX_s_1_2_2((nand_684_nl), nand_772_cse, or_11_cse);
  assign nl_inp_lookup_1_FpNormalize_8U_49U_else_acc_nl = reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_7_1_itm
      + ({2'b11 , (~ libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_8)})
      + 8'b1;
  assign inp_lookup_1_FpNormalize_8U_49U_else_acc_nl = nl_inp_lookup_1_FpNormalize_8U_49U_else_acc_nl[7:0];
  assign FpNormalize_8U_49U_oelse_not_4_nl = ~ FpNormalize_8U_49U_if_FpNormalize_8U_49U_if_nand_tmp;
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_nl = MUX_v_8_2_2(8'b00000000,
      (inp_lookup_1_FpNormalize_8U_49U_else_acc_nl), (FpNormalize_8U_49U_oelse_not_4_nl));
  assign nl_inp_lookup_1_FpAdd_8U_23U_if_3_if_acc_nl = reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_1_lpi_1_dfm_7_1_itm
      + 8'b1;
  assign inp_lookup_1_FpAdd_8U_23U_if_3_if_acc_nl = nl_inp_lookup_1_FpAdd_8U_23U_if_3_if_acc_nl[7:0];
  assign or_5922_nl = (~ (chn_inp_in_crt_sva_1_739_395_1[341])) | (cfg_precision_1_sva_st_90!=2'b10);
  assign mux_191_nl = MUX_s_1_2_2(nand_602_cse_1, (or_5922_nl), main_stage_v_1);
  assign or_433_nl = main_stage_v_2 | (mux_191_nl);
  assign or_5925_nl = (~ (chn_inp_in_crt_sva_2_739_736_1[0])) | (cfg_precision_1_sva_st_91!=2'b10);
  assign mux_2057_nl = MUX_s_1_2_2(nand_694_cse, (or_5925_nl), main_stage_v_2);
  assign or_436_nl = main_stage_v_3 | (mux_2057_nl);
  assign mux_200_nl = MUX_s_1_2_2((or_436_nl), (or_433_nl), or_11_cse);
  assign and_3359_nl = ((chn_inp_in_crt_sva_2_739_736_1!=4'b0000)) & main_stage_v_2;
  assign and_3360_nl = ((chn_inp_in_crt_sva_3_739_736_1!=4'b0000)) & main_stage_v_3;
  assign mux_201_nl = MUX_s_1_2_2((and_3360_nl), (and_3359_nl), or_11_cse);
  assign inp_lookup_1_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_1_sva[30:1]),
      30'b111111111111111111111111111111, IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_ovfl_1_sva));
  assign inp_lookup_1_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_nl
      = ~((~((IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_1_sva[0]) | IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_ovfl_1_sva))
      | IntSignedShiftRight_50U_5U_32U_obits_fixed_and_unfl_1_sva);
  assign mux_206_nl = MUX_s_1_2_2(and_tmp_33, and_tmp_29, or_11_cse);
  assign mux_207_nl = MUX_s_1_2_2((mux_206_nl), mux_tmp_127, and_3358_cse);
  assign mux_208_nl = MUX_s_1_2_2((mux_207_nl), mux_tmp_127, nor_35_cse);
  assign nor_1639_nl = ~((~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | and_tmp_34);
  assign and_3356_nl = inp_lookup_1_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs
      & (inp_lookup_1_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21]);
  assign mux_216_nl = MUX_s_1_2_2(or_tmp_463, (nor_1639_nl), and_3356_nl);
  assign mux_217_nl = MUX_s_1_2_2((mux_216_nl), or_tmp_463, FpMul_6U_10U_2_lor_6_lpi_1_dfm_st_3);
  assign mux_218_nl = MUX_s_1_2_2(nand_tmp_14, (~ (mux_217_nl)), cfg_precision_1_sva_st_91[1]);
  assign mux_219_nl = MUX_s_1_2_2((mux_218_nl), nand_tmp_14, or_461_cse);
  assign mux_220_nl = MUX_s_1_2_2(nand_tmp_14, (~ or_tmp_463), cfg_precision_1_sva_st_90[1]);
  assign or_468_nl = (chn_inp_in_crt_sva_1_739_395_1[341]) | (cfg_precision_1_sva_st_90[0]);
  assign mux_221_nl = MUX_s_1_2_2((mux_220_nl), nand_tmp_14, or_468_nl);
  assign nand_15_nl = ~(main_stage_v_3 & (~ or_tmp_461));
  assign mux_222_nl = MUX_s_1_2_2((nand_15_nl), or_471_cse, or_11_cse);
  assign mux_223_nl = MUX_s_1_2_2((mux_222_nl), (mux_221_nl), main_stage_v_1);
  assign mux_224_nl = MUX_s_1_2_2((mux_223_nl), (mux_219_nl), main_stage_v_2);
  assign or_474_nl = (~ inp_lookup_1_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4)
      | FpMul_6U_10U_2_lor_6_lpi_1_dfm_st_4 | (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[0])
      | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_225_nl = MUX_s_1_2_2((or_474_nl), or_5800_cse, or_11_cse);
  assign or_476_nl = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ inp_lookup_1_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4)
      | FpMul_6U_10U_2_lor_6_lpi_1_dfm_st_4 | (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[0])
      | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_226_nl = MUX_s_1_2_2((or_476_nl), (mux_225_nl), nor_44_cse);
  assign or_478_nl = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | FpMul_6U_10U_2_lor_6_lpi_1_dfm_st_4 | (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[0])
      | (cfg_precision_1_sva_st_80!=2'b10);
  assign or_481_nl = FpMul_6U_10U_2_lor_6_lpi_1_dfm_st_4 | (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[0])
      | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_227_nl = MUX_s_1_2_2((or_481_nl), or_5800_cse, or_11_cse);
  assign mux_228_nl = MUX_s_1_2_2((mux_227_nl), (or_478_nl), FpMul_6U_10U_2_lor_6_lpi_1_dfm_st_3);
  assign or_483_nl = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ main_stage_v_3) | (~ (chn_inp_in_crt_sva_3_739_736_1[1])) | (FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_3_49_1_1[48])
      | FpMul_6U_10U_1_lor_7_lpi_1_dfm_5 | (cfg_precision_1_sva_st_80!=2'b10) | inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4;
  assign or_485_nl = (~ main_stage_v_3) | (~ (chn_inp_in_crt_sva_3_739_736_1[1]))
      | (FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_3_49_1_1[48]) | FpMul_6U_10U_1_lor_7_lpi_1_dfm_5
      | (cfg_precision_1_sva_st_80!=2'b10) | inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4;
  assign mux_229_nl = MUX_s_1_2_2((or_485_nl), nand_358_cse, or_11_cse);
  assign or_482_nl = FpNormalize_8U_49U_if_FpNormalize_8U_49U_if_nand_1_tmp | (z_out_1[49]);
  assign mux_230_nl = MUX_s_1_2_2((mux_229_nl), (or_483_nl), or_482_nl);
  assign or_4352_nl = (~ (chn_inp_in_crt_sva_3_739_736_1[1])) | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_1874_nl = MUX_s_1_2_2(nand_358_cse, (or_4352_nl), main_stage_v_3);
  assign FpAdd_8U_23U_o_mant_not_1_nl = ~ (fsm_output[0]);
  assign and_3422_nl = MUX_v_23_2_2(23'b00000000000000000000000, FpAdd_8U_23U_FpAdd_8U_23U_or_5_itm,
      (FpAdd_8U_23U_o_mant_not_1_nl));
  assign and_931_nl = and_dcpl_423 & (chn_inp_in_crt_sva_2_739_736_1[1]) & and_dcpl_419
      & (fsm_output[1]);
  assign mux_2227_nl = MUX_s_1_2_2(or_tmp_4831, mux_tmp_2075, or_6252_cse);
  assign nor_1976_nl = ~((cfg_precision_1_sva_st_90[1]) | (~ mux_tmp_2075));
  assign mux_2228_nl = MUX_s_1_2_2((nor_1976_nl), mux_tmp_2075, or_6257_cse);
  assign and_4231_nl = nand_728_cse_1 & mux_tmp_2075;
  assign mux_2229_nl = MUX_s_1_2_2((and_4231_nl), (mux_2228_nl), main_stage_v_1);
  assign mux_2230_nl = MUX_s_1_2_2((mux_2229_nl), (mux_2227_nl), main_stage_v_2);
  assign mux_2231_nl = MUX_s_1_2_2(or_tmp_4831, (fsm_output[0]), or_6252_cse);
  assign mux_2232_nl = MUX_s_1_2_2(not_tmp_3015, (fsm_output[0]), or_6257_cse);
  assign and_4239_nl = nand_728_cse_1 & (fsm_output[0]);
  assign mux_2233_nl = MUX_s_1_2_2((and_4239_nl), (mux_2232_nl), main_stage_v_1);
  assign mux_2234_nl = MUX_s_1_2_2((mux_2233_nl), (mux_2231_nl), main_stage_v_2);
  assign mux_2235_nl = MUX_s_1_2_2((mux_2234_nl), (mux_2230_nl), main_stage_v_3);
  assign and_4232_nl = (fsm_output[0]) & or_tmp_4829;
  assign and_4240_nl = or_6252_cse & (fsm_output[0]);
  assign or_6265_nl = (~ main_stage_v_1) | (~ (chn_inp_in_crt_sva_1_739_395_1[342]))
      | (cfg_precision_1_sva_st_90[0]);
  assign mux_2236_nl = MUX_s_1_2_2(not_tmp_3015, (fsm_output[0]), or_6265_nl);
  assign mux_2237_nl = MUX_s_1_2_2((mux_2236_nl), (and_4240_nl), main_stage_v_2);
  assign mux_2238_nl = MUX_s_1_2_2((mux_2237_nl), (and_4232_nl), main_stage_v_3);
  assign mux_2239_nl = MUX_s_1_2_2((mux_2238_nl), (mux_2235_nl), or_11_cse);
  assign or_6266_nl = (~ main_stage_v_3) | IsNaN_6U_10U_6_land_2_lpi_1_dfm_5 | IsNaN_6U_10U_7_land_2_lpi_1_dfm_6;
  assign mux_2240_nl = MUX_s_1_2_2(or_tmp_4830, (fsm_output[0]), or_6266_nl);
  assign mux_2241_nl = MUX_s_1_2_2((mux_2240_nl), (mux_2239_nl), fsm_output[1]);
  assign nand_599_nl = ~(main_stage_v_3 & (chn_inp_in_crt_sva_3_739_736_1[1]) & (cfg_precision_1_sva_st_80==2'b10));
  assign mux_236_nl = MUX_s_1_2_2((nand_599_nl), nand_358_cse, or_11_cse);
  assign nl_inp_lookup_2_FpNormalize_8U_49U_else_acc_nl = reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_7_1_itm
      + ({2'b11 , (~ libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_9)})
      + 8'b1;
  assign inp_lookup_2_FpNormalize_8U_49U_else_acc_nl = nl_inp_lookup_2_FpNormalize_8U_49U_else_acc_nl[7:0];
  assign FpNormalize_8U_49U_oelse_not_5_nl = ~ FpNormalize_8U_49U_if_FpNormalize_8U_49U_if_nand_1_tmp;
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_2_nl = MUX_v_8_2_2(8'b00000000,
      (inp_lookup_2_FpNormalize_8U_49U_else_acc_nl), (FpNormalize_8U_49U_oelse_not_5_nl));
  assign nl_inp_lookup_2_FpAdd_8U_23U_if_3_if_acc_nl = reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_2_lpi_1_dfm_7_1_itm
      + 8'b1;
  assign inp_lookup_2_FpAdd_8U_23U_if_3_if_acc_nl = nl_inp_lookup_2_FpAdd_8U_23U_if_3_if_acc_nl[7:0];
  assign or_5933_nl = (~ (chn_inp_in_crt_sva_1_739_395_1[342])) | (cfg_precision_1_sva_st_90!=2'b10);
  assign mux_231_nl = MUX_s_1_2_2(nand_728_cse_1, (or_5933_nl), main_stage_v_1);
  assign or_498_nl = main_stage_v_2 | (mux_231_nl);
  assign mux_2062_nl = MUX_s_1_2_2(or_tmp_213, or_6252_cse, main_stage_v_2);
  assign or_499_nl = main_stage_v_3 | (mux_2062_nl);
  assign mux_238_nl = MUX_s_1_2_2((or_499_nl), (or_498_nl), or_11_cse);
  assign inp_lookup_2_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_2_sva[30:1]),
      30'b111111111111111111111111111111, IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_ovfl_2_sva));
  assign inp_lookup_2_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_nl
      = ~((~((IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_2_sva[0]) | IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_ovfl_2_sva))
      | IntSignedShiftRight_50U_5U_32U_obits_fixed_and_unfl_2_sva);
  assign mux_244_nl = MUX_s_1_2_2(and_tmp_38, and_tmp_35, or_11_cse);
  assign mux_245_nl = MUX_s_1_2_2(mux_tmp_165, (mux_244_nl), or_507_cse);
  assign mux_246_nl = MUX_s_1_2_2((mux_245_nl), mux_tmp_165, and_3355_cse);
  assign nor_1637_nl = ~((~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | and_tmp_39);
  assign and_3352_nl = inp_lookup_2_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs
      & (inp_lookup_2_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21]);
  assign mux_254_nl = MUX_s_1_2_2(or_tmp_525, (nor_1637_nl), and_3352_nl);
  assign mux_255_nl = MUX_s_1_2_2((mux_254_nl), or_tmp_525, FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_3);
  assign mux_256_nl = MUX_s_1_2_2(nand_tmp_16, (~ (mux_255_nl)), cfg_precision_1_sva_st_91[1]);
  assign mux_257_nl = MUX_s_1_2_2((mux_256_nl), nand_tmp_16, or_523_cse);
  assign mux_258_nl = MUX_s_1_2_2(nand_tmp_16, (~ or_tmp_525), cfg_precision_1_sva_st_90[1]);
  assign or_530_nl = (chn_inp_in_crt_sva_1_739_395_1[342]) | (cfg_precision_1_sva_st_90[0]);
  assign mux_259_nl = MUX_s_1_2_2((mux_258_nl), nand_tmp_16, or_530_nl);
  assign nor_1638_nl = ~((~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (main_stage_v_3 & (~ or_tmp_523)));
  assign mux_260_nl = MUX_s_1_2_2(nand_tmp_16, (nor_1638_nl), chn_inp_in_rsci_bawt);
  assign or_531_nl = (chn_inp_in_rsci_d_mxwt[737]) | (cfg_precision_rsci_d!=2'b10);
  assign mux_261_nl = MUX_s_1_2_2((mux_260_nl), nand_tmp_16, or_531_nl);
  assign mux_262_nl = MUX_s_1_2_2((mux_261_nl), (mux_259_nl), main_stage_v_1);
  assign mux_263_nl = MUX_s_1_2_2((mux_262_nl), (mux_257_nl), main_stage_v_2);
  assign or_535_nl = (~ inp_lookup_2_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4)
      | FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_4 | (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[1])
      | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_264_nl = MUX_s_1_2_2((or_535_nl), or_tmp_238, or_11_cse);
  assign nor_1959_nl = ~((~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[1])
      | (cfg_precision_1_sva_st_91!=2'b10) | FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_3);
  assign nor_1960_nl = ~(FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_4 | (~ main_stage_v_3)
      | (chn_inp_in_crt_sva_3_739_736_1[1]) | (cfg_precision_1_sva_st_80!=2'b10));
  assign mux_265_nl = MUX_s_1_2_2((nor_1960_nl), (nor_1959_nl), or_11_cse);
  assign or_539_nl = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ main_stage_v_3) | (~ (chn_inp_in_crt_sva_3_739_736_1[2])) | (FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_3_49_1_1[48])
      | (cfg_precision_1_sva_st_80!=2'b10) | FpMul_6U_10U_1_lor_8_lpi_1_dfm_5 | inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4;
  assign or_541_nl = (~ main_stage_v_3) | (~ (chn_inp_in_crt_sva_3_739_736_1[2]))
      | (FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_3_49_1_1[48]) | (cfg_precision_1_sva_st_80!=2'b10)
      | FpMul_6U_10U_1_lor_8_lpi_1_dfm_5 | inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4;
  assign mux_266_nl = MUX_s_1_2_2((or_541_nl), or_tmp_277, or_11_cse);
  assign or_538_nl = FpNormalize_8U_49U_if_FpNormalize_8U_49U_if_nand_2_tmp | (z_out_2[49]);
  assign mux_267_nl = MUX_s_1_2_2((mux_266_nl), (or_539_nl), or_538_nl);
  assign or_4363_nl = (~ (chn_inp_in_crt_sva_3_739_736_1[2])) | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_1880_nl = MUX_s_1_2_2(or_tmp_277, (or_4363_nl), main_stage_v_3);
  assign FpAdd_8U_23U_o_mant_not_2_nl = ~ (fsm_output[0]);
  assign and_3423_nl = MUX_v_23_2_2(23'b00000000000000000000000, FpAdd_8U_23U_FpAdd_8U_23U_or_6_itm,
      (FpAdd_8U_23U_o_mant_not_2_nl));
  assign and_969_nl = and_dcpl_498 & and_dcpl_496 & (fsm_output[1]);
  assign mux_2243_nl = MUX_s_1_2_2(mux_tmp_2091, or_tmp_4843, nor_1967_cse);
  assign nor_1974_nl = ~((cfg_precision_1_sva_st_90[1]) | (~ mux_tmp_2091));
  assign mux_2244_nl = MUX_s_1_2_2((nor_1974_nl), mux_tmp_2091, or_6272_cse);
  assign and_4234_nl = nand_598_cse & mux_tmp_2091;
  assign mux_2245_nl = MUX_s_1_2_2((and_4234_nl), (mux_2244_nl), main_stage_v_1);
  assign mux_2246_nl = MUX_s_1_2_2((mux_2245_nl), (mux_2243_nl), main_stage_v_2);
  assign mux_2247_nl = MUX_s_1_2_2((fsm_output[0]), or_tmp_4843, nor_1967_cse);
  assign mux_2248_nl = MUX_s_1_2_2(not_tmp_3015, (fsm_output[0]), or_6272_cse);
  assign and_4242_nl = nand_598_cse & (fsm_output[0]);
  assign mux_2249_nl = MUX_s_1_2_2((and_4242_nl), (mux_2248_nl), main_stage_v_1);
  assign mux_2250_nl = MUX_s_1_2_2((mux_2249_nl), (mux_2247_nl), main_stage_v_2);
  assign mux_2251_nl = MUX_s_1_2_2((mux_2250_nl), (mux_2246_nl), main_stage_v_3);
  assign and_4235_nl = (fsm_output[0]) & or_tmp_4845;
  assign or_6278_nl = (~ (chn_inp_in_crt_sva_2_739_736_1[2])) | (cfg_precision_1_sva_st_91[0]);
  assign mux_2252_nl = MUX_s_1_2_2(nor_1978_cse, (fsm_output[0]), or_6278_nl);
  assign or_6280_nl = (~ main_stage_v_1) | (~ (chn_inp_in_crt_sva_1_739_395_1[343]))
      | (cfg_precision_1_sva_st_90[0]);
  assign mux_2253_nl = MUX_s_1_2_2(not_tmp_3015, (fsm_output[0]), or_6280_nl);
  assign mux_2254_nl = MUX_s_1_2_2((mux_2253_nl), (mux_2252_nl), main_stage_v_2);
  assign mux_2255_nl = MUX_s_1_2_2((mux_2254_nl), (and_4235_nl), main_stage_v_3);
  assign mux_2256_nl = MUX_s_1_2_2((mux_2255_nl), (mux_2251_nl), or_11_cse);
  assign or_6281_nl = (~ main_stage_v_3) | IsNaN_6U_10U_6_land_3_lpi_1_dfm_5 | IsNaN_6U_10U_7_land_3_lpi_1_dfm_6;
  assign mux_2257_nl = MUX_s_1_2_2(or_tmp_4846, (fsm_output[0]), or_6281_nl);
  assign mux_2258_nl = MUX_s_1_2_2((mux_2257_nl), (mux_2256_nl), fsm_output[1]);
  assign nand_597_nl = ~(main_stage_v_3 & (chn_inp_in_crt_sva_3_739_736_1[2]) & (cfg_precision_1_sva_st_80==2'b10));
  assign mux_273_nl = MUX_s_1_2_2((nand_597_nl), or_tmp_277, or_11_cse);
  assign nl_inp_lookup_3_FpNormalize_8U_49U_else_acc_nl = reg_FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_7_1_itm
      + ({2'b11 , (~ libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_10)})
      + 8'b1;
  assign inp_lookup_3_FpNormalize_8U_49U_else_acc_nl = nl_inp_lookup_3_FpNormalize_8U_49U_else_acc_nl[7:0];
  assign FpNormalize_8U_49U_oelse_not_6_nl = ~ FpNormalize_8U_49U_if_FpNormalize_8U_49U_if_nand_2_tmp;
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_4_nl = MUX_v_8_2_2(8'b00000000,
      (inp_lookup_3_FpNormalize_8U_49U_else_acc_nl), (FpNormalize_8U_49U_oelse_not_6_nl));
  assign nl_inp_lookup_3_FpAdd_8U_23U_if_3_if_acc_nl = reg_FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_mant_3_lpi_1_dfm_7_1_itm
      + 8'b1;
  assign inp_lookup_3_FpAdd_8U_23U_if_3_if_acc_nl = nl_inp_lookup_3_FpAdd_8U_23U_if_3_if_acc_nl[7:0];
  assign or_557_nl = main_stage_v_3 | (~ (chn_inp_in_crt_sva_2_739_736_1[2])) | (cfg_precision_1_sva_st_91!=2'b10)
      | (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt;
  assign or_560_nl = (~ (chn_inp_in_crt_sva_1_739_395_1[343])) | (cfg_precision_1_sva_st_90[0])
      | (~((cfg_precision_1_sva_st_90[1]) & ((~ main_stage_v_3) | (~ reg_chn_inp_out_rsci_ld_core_psct_cse)
      | chn_inp_out_rsci_bawt)));
  assign or_563_nl = (~ (chn_inp_in_rsci_d_mxwt[738])) | (cfg_precision_rsci_d!=2'b10)
      | (~(chn_inp_in_rsci_bawt & or_11_cse));
  assign mux_275_nl = MUX_s_1_2_2((or_563_nl), (or_560_nl), main_stage_v_1);
  assign mux_276_nl = MUX_s_1_2_2((mux_275_nl), (or_557_nl), main_stage_v_2);
  assign inp_lookup_3_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_3_sva[30:1]),
      30'b111111111111111111111111111111, IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_ovfl_3_sva));
  assign inp_lookup_3_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_nl
      = ~((~((IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_3_sva[0]) | IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_ovfl_3_sva))
      | IntSignedShiftRight_50U_5U_32U_obits_fixed_and_unfl_3_sva);
  assign mux_282_nl = MUX_s_1_2_2(and_tmp_45, and_tmp_42, or_11_cse);
  assign mux_283_nl = MUX_s_1_2_2((mux_282_nl), mux_tmp_203, nor_55_cse);
  assign mux_284_nl = MUX_s_1_2_2((mux_283_nl), mux_tmp_203, and_3351_cse);
  assign nor_1632_nl = ~((~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | and_tmp_49);
  assign and_3347_nl = inp_lookup_3_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs
      & (inp_lookup_3_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21]);
  assign mux_299_nl = MUX_s_1_2_2(or_tmp_599, (nor_1632_nl), and_3347_nl);
  assign mux_300_nl = MUX_s_1_2_2((mux_299_nl), or_tmp_599, FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_3);
  assign mux_301_nl = MUX_s_1_2_2(nand_tmp_20, (~ (mux_300_nl)), cfg_precision_1_sva_st_91[1]);
  assign mux_302_nl = MUX_s_1_2_2((mux_301_nl), nand_tmp_20, or_597_cse);
  assign mux_303_nl = MUX_s_1_2_2(nand_tmp_20, (~ or_tmp_599), cfg_precision_1_sva_st_90[1]);
  assign mux_304_nl = MUX_s_1_2_2((mux_303_nl), nand_tmp_20, or_604_cse);
  assign nor_1633_nl = ~((~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (main_stage_v_3 & (~ or_tmp_597)));
  assign mux_305_nl = MUX_s_1_2_2(nand_tmp_20, (nor_1633_nl), chn_inp_in_rsci_bawt);
  assign or_605_nl = (chn_inp_in_rsci_d_mxwt[738]) | (cfg_precision_rsci_d!=2'b10);
  assign mux_306_nl = MUX_s_1_2_2((mux_305_nl), nand_tmp_20, or_605_nl);
  assign mux_307_nl = MUX_s_1_2_2((mux_306_nl), (mux_304_nl), main_stage_v_1);
  assign mux_308_nl = MUX_s_1_2_2((mux_307_nl), (mux_302_nl), main_stage_v_2);
  assign or_609_nl = (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[2]) | (~
      inp_lookup_3_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4)
      | FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_4 | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_309_nl = MUX_s_1_2_2((or_609_nl), or_tmp_306, or_11_cse);
  assign or_610_nl = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[2]) | (~ inp_lookup_3_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4)
      | FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_4 | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_310_nl = MUX_s_1_2_2((or_610_nl), (mux_309_nl), nor_67_cse);
  assign or_611_nl = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[2]) | FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_4
      | (cfg_precision_1_sva_st_80!=2'b10);
  assign or_613_nl = (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[2]) | FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_4
      | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_311_nl = MUX_s_1_2_2((or_613_nl), or_tmp_306, or_11_cse);
  assign mux_312_nl = MUX_s_1_2_2((mux_311_nl), (or_611_nl), FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_3);
  assign nor_1630_nl = ~((~ main_stage_v_2) | (~ (chn_inp_in_crt_sva_2_739_736_1[3]))
      | (cfg_precision_1_sva_st_91!=2'b10) | FpNormalize_8U_49U_if_FpNormalize_8U_49U_if_nand_3_tmp
      | (z_out_3[49]));
  assign nor_1631_nl = ~((~ main_stage_v_3) | (~ (chn_inp_in_crt_sva_3_739_736_1[3]))
      | (cfg_precision_1_sva_st_80!=2'b10) | (FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_3_49_1_1[48])
      | FpMul_6U_10U_1_lor_1_lpi_1_dfm_5 | inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4);
  assign mux_313_nl = MUX_s_1_2_2((nor_1631_nl), (nor_1630_nl), or_11_cse);
  assign mux_314_nl = MUX_s_1_2_2(nand_661_cse, nand_701_cse, or_11_cse);
  assign nl_inp_lookup_4_FpNormalize_8U_49U_else_acc_nl = reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_7_1_itm
      + ({2'b11 , (~ libraries_leading_sign_49_0_78e877fc94067377fcee479dbb0ed8e083a3_11)})
      + 8'b1;
  assign inp_lookup_4_FpNormalize_8U_49U_else_acc_nl = nl_inp_lookup_4_FpNormalize_8U_49U_else_acc_nl[7:0];
  assign FpNormalize_8U_49U_oelse_not_7_nl = ~ FpNormalize_8U_49U_if_FpNormalize_8U_49U_if_nand_3_tmp;
  assign FpNormalize_8U_49U_FpNormalize_8U_49U_and_6_nl = MUX_v_8_2_2(8'b00000000,
      (inp_lookup_4_FpNormalize_8U_49U_else_acc_nl), (FpNormalize_8U_49U_oelse_not_7_nl));
  assign nl_inp_lookup_4_FpAdd_8U_23U_if_3_if_acc_nl = reg_FpExpoWidthInc_5U_6U_10U_1U_1U_3_o_mant_lpi_1_dfm_7_1_itm
      + 8'b1;
  assign inp_lookup_4_FpAdd_8U_23U_if_3_if_acc_nl = nl_inp_lookup_4_FpAdd_8U_23U_if_3_if_acc_nl[7:0];
  assign mux_316_nl = MUX_s_1_2_2(or_tmp_621, or_2010_cse, main_stage_v_1);
  assign or_624_nl = main_stage_v_1 | (~ (chn_inp_in_rsci_d_mxwt[739])) | (~ chn_inp_in_rsci_bawt)
      | (cfg_precision_rsci_d!=2'b10);
  assign mux_317_nl = MUX_s_1_2_2((or_624_nl), (mux_316_nl), chn_inp_in_crt_sva_1_739_395_1[344]);
  assign or_625_nl = main_stage_v_2 | (mux_317_nl);
  assign or_627_nl = (~ (chn_inp_in_crt_sva_2_739_736_1[3])) | (cfg_precision_1_sva_st_91!=2'b10);
  assign mux_318_nl = MUX_s_1_2_2(or_tmp_347, (or_627_nl), main_stage_v_2);
  assign or_628_nl = main_stage_v_3 | (mux_318_nl);
  assign mux_319_nl = MUX_s_1_2_2((or_628_nl), (or_625_nl), or_11_cse);
  assign inp_lookup_4_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_2_nl = ~(MUX_v_30_2_2((IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_sva[30:1]),
      30'b111111111111111111111111111111, IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_ovfl_sva));
  assign inp_lookup_4_IntSignedShiftRight_50U_5U_32U_obits_fixed_IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_1_nl
      = ~((~((IntSignedShiftRight_50U_5U_32U_obits_fixed_acc_sat_sva[0]) | IntSignedShiftRight_50U_5U_32U_obits_fixed_nor_ovfl_sva))
      | IntSignedShiftRight_50U_5U_32U_obits_fixed_and_unfl_sva);
  assign mux_1992_nl = MUX_s_1_2_2(mux_tmp_250, (~ mux_tmp_247), main_stage_v_2);
  assign mux_331_nl = MUX_s_1_2_2((mux_1992_nl), mux_tmp_250, chn_inp_in_crt_sva_2_739_736_1[3]);
  assign mux_330_nl = MUX_s_1_2_2(mux_tmp_250, (~ mux_tmp_247), main_stage_v_2);
  assign or_637_nl = inp_lookup_4_FpMul_6U_10U_1_oelse_1_acc_itm_7_1 | FpMul_6U_10U_1_if_2_FpMul_6U_10U_1_if_2_or_6_tmp
      | (~ inp_lookup_4_FpMul_6U_10U_1_else_2_if_acc_itm_6_1) | (chn_inp_in_crt_sva_2_739_736_1[3]);
  assign mux_332_nl = MUX_s_1_2_2((mux_330_nl), mux_tmp_250, or_637_nl);
  assign mux_333_nl = MUX_s_1_2_2((mux_332_nl), (mux_331_nl), and_3345_cse);
  assign mux_334_nl = MUX_s_1_2_2(mux_tmp_251, (~ (mux_333_nl)), cfg_precision_1_sva_st_91[1]);
  assign mux_335_nl = MUX_s_1_2_2((mux_334_nl), mux_tmp_251, cfg_precision_1_sva_st_91[0]);
  assign nor_1626_nl = ~((~((~(FpMul_6U_10U_2_lor_1_lpi_1_dfm_st_3 | (~ inp_lookup_4_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs)
      | (~ (inp_lookup_4_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21])))) | (chn_inp_in_crt_sva_2_739_736_1[3])))
      | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10));
  assign nor_1628_nl = ~((~ main_stage_v_3) | (cfg_precision_1_sva_st_80[0]) | (~((cfg_precision_1_sva_st_80[1])
      & ((~(FpMul_6U_10U_2_lor_1_lpi_1_dfm_st_4 | (~ inp_lookup_4_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4)
      | (~ inp_lookup_4_FpMul_6U_10U_2_else_2_else_slc_FpMul_6U_10U_2_p_mant_p1_21_itm_2)))
      | (chn_inp_in_crt_sva_3_739_736_1[3])))));
  assign mux_347_nl = MUX_s_1_2_2((nor_1628_nl), (nor_1626_nl), or_11_cse);
  assign or_663_nl = (~ main_stage_v_3) | (~ inp_lookup_4_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4)
      | FpMul_6U_10U_2_lor_1_lpi_1_dfm_st_4 | (chn_inp_in_crt_sva_3_739_736_1[3])
      | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_348_nl = MUX_s_1_2_2((or_663_nl), or_tmp_374, or_11_cse);
  assign nor_1957_nl = ~(FpMul_6U_10U_2_lor_1_lpi_1_dfm_st_3 | (~ main_stage_v_2)
      | (chn_inp_in_crt_sva_2_739_736_1[3]) | (cfg_precision_1_sva_st_91!=2'b10));
  assign nor_1958_nl = ~((~ main_stage_v_3) | FpMul_6U_10U_2_lor_1_lpi_1_dfm_st_4
      | (chn_inp_in_crt_sva_3_739_736_1[3]) | (cfg_precision_1_sva_st_80!=2'b10));
  assign mux_349_nl = MUX_s_1_2_2((nor_1958_nl), (nor_1957_nl), or_11_cse);
  assign or_667_nl = (cfg_precision_1_sva_st_80!=2'b10) | FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_3;
  assign mux_350_nl = MUX_s_1_2_2((or_667_nl), or_tmp_440, chn_inp_in_crt_sva_3_739_736_1[0]);
  assign and_3342_nl = main_stage_v_3 & (~ (mux_350_nl));
  assign and_3343_nl = main_stage_v_4 & (~((~((~ FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_4)
      | (chn_inp_in_crt_sva_4_739_736_1[0]))) | (cfg_precision_1_sva_st_81!=2'b10)));
  assign mux_351_nl = MUX_s_1_2_2((and_3343_nl), (and_3342_nl), or_11_cse);
  assign FpMul_6U_10U_1_FpMul_6U_10U_1_and_nl = (inp_lookup_1_FpMul_6U_10U_1_else_2_else_if_if_acc_1_itm_5_1
      | (~ FpMul_6U_10U_1_p_mant_p1_1_sva_mx2_21)) & inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4;
  assign or_697_nl = (chn_inp_in_crt_sva_3_739_736_1[0]) | (cfg_precision_1_sva_st_80[0])
      | not_tmp_282;
  assign mux_357_nl = MUX_s_1_2_2(or_471_cse, or_683_cse, main_stage_v_1);
  assign mux_358_nl = MUX_s_1_2_2((mux_357_nl), or_tmp_679, main_stage_v_2);
  assign mux_368_nl = MUX_s_1_2_2((mux_358_nl), (or_697_nl), main_stage_v_3);
  assign or_699_nl = (chn_inp_in_crt_sva_4_739_736_1[0]) | (cfg_precision_1_sva_st_81!=2'b10)
      | (~ IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_16);
  assign or_687_nl = (chn_inp_in_crt_sva_3_739_736_1[0]) | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_360_nl = MUX_s_1_2_2(or_tmp_21, or_tmp_679, main_stage_v_2);
  assign mux_361_nl = MUX_s_1_2_2((mux_360_nl), (or_687_nl), main_stage_v_3);
  assign mux_369_nl = MUX_s_1_2_2((mux_361_nl), (or_699_nl), main_stage_v_4);
  assign mux_370_nl = MUX_s_1_2_2((mux_369_nl), (mux_368_nl), or_11_cse);
  assign nor_1619_nl = ~((~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | and_tmp_54);
  assign or_704_nl = (~ IsNaN_6U_10U_5_land_1_lpi_1_dfm_5) | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_15;
  assign mux_371_nl = MUX_s_1_2_2((nor_1619_nl), or_tmp_704, or_704_nl);
  assign mux_372_nl = MUX_s_1_2_2(nand_tmp_29, (~ (mux_371_nl)), cfg_precision_1_sva_st_80[1]);
  assign or_700_nl = (chn_inp_in_crt_sva_3_739_736_1[0]) | (cfg_precision_1_sva_st_80[0]);
  assign mux_373_nl = MUX_s_1_2_2((mux_372_nl), nand_tmp_29, or_700_nl);
  assign mux_374_nl = MUX_s_1_2_2(nand_tmp_29, (~ or_tmp_704), cfg_precision_1_sva_st_91[1]);
  assign mux_375_nl = MUX_s_1_2_2((mux_374_nl), nand_tmp_29, or_461_cse);
  assign mux_376_nl = MUX_s_1_2_2((~ or_tmp_704), nand_tmp_29, or_683_cse);
  assign nor_1620_nl = ~((~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (main_stage_v_4 & (~ or_tmp_701)));
  assign mux_377_nl = MUX_s_1_2_2((nor_1620_nl), nand_tmp_29, or_471_cse);
  assign mux_378_nl = MUX_s_1_2_2((mux_377_nl), (mux_376_nl), main_stage_v_1);
  assign mux_379_nl = MUX_s_1_2_2((mux_378_nl), (mux_375_nl), main_stage_v_2);
  assign mux_380_nl = MUX_s_1_2_2((mux_379_nl), (mux_373_nl), main_stage_v_3);
  assign and_3337_nl = main_stage_v_3 & (~((~((chn_inp_in_crt_sva_3_739_736_1[1])
      | (~ FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_3))) | (cfg_precision_1_sva_st_80!=2'b10)));
  assign and_3338_nl = main_stage_v_4 & (~((~((chn_inp_in_crt_sva_4_739_736_1[1])
      | (~ FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_4))) | (cfg_precision_1_sva_st_81!=2'b10)));
  assign mux_382_nl = MUX_s_1_2_2((and_3338_nl), (and_3337_nl), or_11_cse);
  assign FpMul_6U_10U_1_FpMul_6U_10U_1_and_16_nl = (inp_lookup_2_FpMul_6U_10U_1_else_2_else_if_if_acc_1_itm_5_1
      | (~ FpMul_6U_10U_1_p_mant_p1_2_sva_mx2_21)) & inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4;
  assign FpMul_6U_10U_2_o_mant_or_nl = FpAdd_8U_23U_or_1_cse | and_dcpl_593;
  assign or_749_nl = (chn_inp_in_crt_sva_3_739_736_1[1]) | (cfg_precision_1_sva_st_80!=2'b10)
      | (~ IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_15);
  assign mux_401_nl = MUX_s_1_2_2(mux_400_cse, or_tmp_736, main_stage_v_2);
  assign mux_408_nl = MUX_s_1_2_2((mux_401_nl), (or_749_nl), main_stage_v_3);
  assign or_751_nl = (chn_inp_in_crt_sva_4_739_736_1[1]) | (cfg_precision_1_sva_st_81!=2'b10)
      | (~ IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_16);
  assign or_737_nl = (chn_inp_in_crt_sva_3_739_736_1[1]) | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_403_nl = MUX_s_1_2_2(or_tmp_52, or_tmp_736, main_stage_v_2);
  assign mux_404_nl = MUX_s_1_2_2((mux_403_nl), (or_737_nl), main_stage_v_3);
  assign mux_409_nl = MUX_s_1_2_2((mux_404_nl), (or_751_nl), main_stage_v_4);
  assign mux_410_nl = MUX_s_1_2_2((mux_409_nl), (mux_408_nl), or_11_cse);
  assign nor_1612_nl = ~((~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | and_tmp_56);
  assign or_756_nl = (~ IsNaN_6U_10U_5_land_2_lpi_1_dfm_5) | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_15;
  assign mux_411_nl = MUX_s_1_2_2((nor_1612_nl), or_tmp_756, or_756_nl);
  assign mux_412_nl = MUX_s_1_2_2(nand_tmp_37, (~ (mux_411_nl)), cfg_precision_1_sva_st_80[1]);
  assign or_752_nl = (chn_inp_in_crt_sva_3_739_736_1[1]) | (cfg_precision_1_sva_st_80[0]);
  assign mux_413_nl = MUX_s_1_2_2((mux_412_nl), nand_tmp_37, or_752_nl);
  assign mux_414_nl = MUX_s_1_2_2(nand_tmp_37, (~ or_tmp_756), cfg_precision_1_sva_st_91[1]);
  assign mux_415_nl = MUX_s_1_2_2((mux_414_nl), nand_tmp_37, or_523_cse);
  assign mux_416_nl = MUX_s_1_2_2((~ or_tmp_756), nand_tmp_37, or_740_cse);
  assign nor_1613_nl = ~((~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (main_stage_v_4 & (~ or_tmp_753)));
  assign mux_417_nl = MUX_s_1_2_2((nor_1613_nl), nand_tmp_37, or_763_cse);
  assign mux_418_nl = MUX_s_1_2_2((mux_417_nl), (mux_416_nl), main_stage_v_1);
  assign mux_419_nl = MUX_s_1_2_2((mux_418_nl), (mux_415_nl), main_stage_v_2);
  assign mux_420_nl = MUX_s_1_2_2((mux_419_nl), (mux_413_nl), main_stage_v_3);
  assign and_3332_nl = main_stage_v_3 & (~((~((chn_inp_in_crt_sva_3_739_736_1[2])
      | (~ FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_3))) | (cfg_precision_1_sva_st_80!=2'b10)));
  assign and_3333_nl = main_stage_v_4 & (~((~((chn_inp_in_crt_sva_4_739_736_1[2])
      | (~ FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_4))) | (cfg_precision_1_sva_st_81!=2'b10)));
  assign mux_422_nl = MUX_s_1_2_2((and_3333_nl), (and_3332_nl), or_11_cse);
  assign FpMul_6U_10U_1_FpMul_6U_10U_1_and_17_nl = (inp_lookup_3_FpMul_6U_10U_1_else_2_else_if_if_acc_1_itm_5_1
      | (~ FpMul_6U_10U_1_p_mant_p1_3_sva_mx2_21)) & inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4;
  assign mux_440_nl = MUX_s_1_2_2(not_tmp_346, IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_15,
      or_11_cse);
  assign mux_441_nl = MUX_s_1_2_2(or_tmp_792, (~ (mux_440_nl)), cfg_precision_1_sva_st_80[1]);
  assign mux_442_nl = MUX_s_1_2_2((mux_441_nl), or_tmp_792, or_792_cse);
  assign mux_443_nl = MUX_s_1_2_2(or_tmp_792, (~ or_tmp_798), cfg_precision_1_sva_st_91[1]);
  assign mux_444_nl = MUX_s_1_2_2((mux_443_nl), or_tmp_792, or_597_cse);
  assign mux_445_nl = MUX_s_1_2_2((~ or_tmp_798), or_tmp_792, or_801_cse);
  assign nor_1606_nl = ~((~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~((~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[2]) | (cfg_precision_1_sva_st_81[0])
      | not_tmp_345)));
  assign mux_446_nl = MUX_s_1_2_2((nor_1606_nl), or_tmp_792, or_802_cse);
  assign mux_447_nl = MUX_s_1_2_2((mux_446_nl), (mux_445_nl), main_stage_v_1);
  assign mux_448_nl = MUX_s_1_2_2((mux_447_nl), (mux_444_nl), main_stage_v_2);
  assign mux_449_nl = MUX_s_1_2_2((mux_448_nl), (mux_442_nl), main_stage_v_3);
  assign nor_1603_nl = ~((~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | and_tmp_59);
  assign or_811_nl = (~ IsNaN_6U_10U_5_land_3_lpi_1_dfm_5) | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_15;
  assign mux_450_nl = MUX_s_1_2_2((nor_1603_nl), or_tmp_811, or_811_nl);
  assign mux_451_nl = MUX_s_1_2_2(nand_tmp_45, (~ (mux_450_nl)), cfg_precision_1_sva_st_80[1]);
  assign mux_452_nl = MUX_s_1_2_2((mux_451_nl), nand_tmp_45, or_792_cse);
  assign mux_453_nl = MUX_s_1_2_2(nand_tmp_45, (~ or_tmp_811), cfg_precision_1_sva_st_91[1]);
  assign mux_454_nl = MUX_s_1_2_2((mux_453_nl), nand_tmp_45, or_597_cse);
  assign mux_455_nl = MUX_s_1_2_2((~ or_tmp_811), nand_tmp_45, or_801_cse);
  assign nor_1604_nl = ~((~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (main_stage_v_4 & (~ or_tmp_808)));
  assign mux_456_nl = MUX_s_1_2_2((nor_1604_nl), nand_tmp_45, or_802_cse);
  assign mux_457_nl = MUX_s_1_2_2((mux_456_nl), (mux_455_nl), main_stage_v_1);
  assign mux_458_nl = MUX_s_1_2_2((mux_457_nl), (mux_454_nl), main_stage_v_2);
  assign mux_459_nl = MUX_s_1_2_2((mux_458_nl), (mux_452_nl), main_stage_v_3);
  assign mux_462_nl = MUX_s_1_2_2(nand_tmp_47, nand_661_cse, or_11_cse);
  assign mux_463_nl = MUX_s_1_2_2(nand_tmp_47, or_2282_cse, or_11_cse);
  assign mux_464_nl = MUX_s_1_2_2((mux_463_nl), (mux_462_nl), FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_3);
  assign FpMul_6U_10U_1_FpMul_6U_10U_1_and_18_nl = (inp_lookup_4_FpMul_6U_10U_1_else_2_else_if_if_acc_1_itm_5_1
      | (~ FpMul_6U_10U_1_p_mant_p1_sva_mx2_21)) & inp_lookup_4_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs_2;
  assign and_3325_nl = main_stage_v_4 & (~((~((chn_inp_in_crt_sva_4_739_736_1[0])
      | (~ FpAdd_6U_10U_1_is_a_greater_acc_itm_6))) | (cfg_precision_1_sva_st_81!=2'b10)));
  assign nor_1595_nl = ~((~((chn_inp_in_crt_sva_5_739_736_1[0]) | (~ chn_inp_in_crt_sva_5_411_1)))
      | (cfg_precision_1_sva_st_82[0]) | not_tmp_374);
  assign mux_471_nl = MUX_s_1_2_2((nor_1595_nl), (and_3325_nl), or_11_cse);
  assign nl_inp_lookup_1_FpAdd_8U_23U_1_if_2_acc_nl = conv_u2u_49_50(FpAdd_8U_23U_1_addend_larger_qr_1_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_1_addend_smaller_qr_1_lpi_1_dfm_mx0);
  assign inp_lookup_1_FpAdd_8U_23U_1_if_2_acc_nl = nl_inp_lookup_1_FpAdd_8U_23U_1_if_2_acc_nl[49:0];
  assign nl_inp_lookup_1_FpAdd_8U_23U_1_else_2_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_1_addend_smaller_qr_1_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_1_addend_larger_qr_1_lpi_1_dfm_mx0) + 50'b1;
  assign inp_lookup_1_FpAdd_8U_23U_1_else_2_acc_nl = nl_inp_lookup_1_FpAdd_8U_23U_1_else_2_acc_nl[49:0];
  assign nand_585_nl = ~(main_stage_v_4 & (chn_inp_in_crt_sva_4_739_736_1[0]) & (cfg_precision_1_sva_st_81==2'b10));
  assign mux_474_nl = MUX_s_1_2_2(or_tmp_850, (nand_585_nl), or_11_cse);
  assign and_4166_nl = ((FpMul_6U_10U_1_o_expo_1_lpi_1_dfm[5:4]!=2'b11) | FpMul_6U_10U_1_lor_6_lpi_1_dfm_6)
      & or_tmp_4675;
  assign mux_2070_nl = MUX_s_1_2_2((and_4166_nl), and_4165_cse, IsNaN_6U_10U_5_land_1_lpi_1_dfm_6);
  assign mux_2071_nl = MUX_s_1_2_2((mux_2070_nl), and_4164_cse, IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_16);
  assign mux_2072_nl = MUX_s_1_2_2(or_tmp_4675, (mux_2071_nl), or_5950_cse);
  assign mux_2073_nl = MUX_s_1_2_2(or_tmp_4675, (mux_2072_nl), and_4141_cse);
  assign and_4138_nl = (~((FpMul_6U_10U_1_o_expo_1_lpi_1_dfm[5:4]==2'b11))) & or_tmp_4675;
  assign mux_2074_nl = MUX_s_1_2_2((and_4138_nl), or_tmp_4675, FpMul_6U_10U_1_lor_6_lpi_1_dfm_6);
  assign mux_2075_nl = MUX_s_1_2_2((mux_2074_nl), and_4165_cse, IsNaN_6U_10U_5_land_1_lpi_1_dfm_6);
  assign mux_2076_nl = MUX_s_1_2_2((mux_2075_nl), and_4164_cse, IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_16);
  assign mux_2077_nl = MUX_s_1_2_2(or_tmp_4675, (mux_2076_nl), or_5950_cse);
  assign mux_2078_nl = MUX_s_1_2_2(or_tmp_4675, (mux_2077_nl), and_4141_cse);
  assign and_3323_nl = main_stage_v_4 & (~((~((chn_inp_in_crt_sva_4_739_736_1[1])
      | (~ FpAdd_6U_10U_1_is_a_greater_acc_1_itm_6))) | (cfg_precision_1_sva_st_81!=2'b10)));
  assign nor_1589_nl = ~((~((~ chn_inp_in_crt_sva_5_427_1) | (chn_inp_in_crt_sva_5_739_736_1[1])))
      | (cfg_precision_1_sva_st_82!=2'b10) | (~ main_stage_v_5));
  assign mux_481_nl = MUX_s_1_2_2((nor_1589_nl), (and_3323_nl), or_11_cse);
  assign nl_inp_lookup_2_FpAdd_8U_23U_1_if_2_acc_nl = conv_u2u_49_50(FpAdd_8U_23U_1_addend_larger_qr_2_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_1_addend_smaller_qr_2_lpi_1_dfm_mx0);
  assign inp_lookup_2_FpAdd_8U_23U_1_if_2_acc_nl = nl_inp_lookup_2_FpAdd_8U_23U_1_if_2_acc_nl[49:0];
  assign nl_inp_lookup_2_FpAdd_8U_23U_1_else_2_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_1_addend_smaller_qr_2_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_1_addend_larger_qr_2_lpi_1_dfm_mx0) + 50'b1;
  assign inp_lookup_2_FpAdd_8U_23U_1_else_2_acc_nl = nl_inp_lookup_2_FpAdd_8U_23U_1_else_2_acc_nl[49:0];
  assign nand_582_nl = ~(main_stage_v_4 & (chn_inp_in_crt_sva_4_739_736_1[1]) & (cfg_precision_1_sva_st_81==2'b10));
  assign mux_484_nl = MUX_s_1_2_2(or_tmp_880, (nand_582_nl), or_11_cse);
  assign and_4161_nl = ((FpMul_6U_10U_1_o_expo_2_lpi_1_dfm[5:4]!=2'b11) | FpMul_6U_10U_1_lor_7_lpi_1_dfm_6)
      & or_tmp_4685;
  assign mux_2079_nl = MUX_s_1_2_2((and_4161_nl), and_4160_cse, IsNaN_6U_10U_5_land_2_lpi_1_dfm_6);
  assign mux_2080_nl = MUX_s_1_2_2((mux_2079_nl), and_4159_cse, IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_16);
  assign mux_2081_nl = MUX_s_1_2_2(or_tmp_4685, (mux_2080_nl), or_5967_cse);
  assign mux_2082_nl = MUX_s_1_2_2(or_tmp_4685, (mux_2081_nl), and_4136_cse);
  assign and_4133_nl = (~((FpMul_6U_10U_1_o_expo_2_lpi_1_dfm[5:4]==2'b11))) & or_tmp_4685;
  assign mux_2083_nl = MUX_s_1_2_2((and_4133_nl), or_tmp_4685, FpMul_6U_10U_1_lor_7_lpi_1_dfm_6);
  assign mux_2084_nl = MUX_s_1_2_2((mux_2083_nl), and_4160_cse, IsNaN_6U_10U_5_land_2_lpi_1_dfm_6);
  assign mux_2085_nl = MUX_s_1_2_2((mux_2084_nl), and_4159_cse, IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_16);
  assign mux_2086_nl = MUX_s_1_2_2(or_tmp_4685, (mux_2085_nl), or_5967_cse);
  assign mux_2087_nl = MUX_s_1_2_2(or_tmp_4685, (mux_2086_nl), and_4136_cse);
  assign mux_490_nl = MUX_s_1_2_2(or_tmp_899, nand_tmp_53, or_11_cse);
  assign mux_491_nl = MUX_s_1_2_2(or_3167_cse, nand_tmp_53, or_11_cse);
  assign mux_492_nl = MUX_s_1_2_2((mux_491_nl), (mux_490_nl), chn_inp_in_crt_sva_5_443_1);
  assign nl_inp_lookup_3_FpAdd_8U_23U_1_if_2_acc_nl = conv_u2u_49_50(FpAdd_8U_23U_1_addend_larger_qr_3_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_1_addend_smaller_qr_3_lpi_1_dfm_mx0);
  assign inp_lookup_3_FpAdd_8U_23U_1_if_2_acc_nl = nl_inp_lookup_3_FpAdd_8U_23U_1_if_2_acc_nl[49:0];
  assign nl_inp_lookup_3_FpAdd_8U_23U_1_else_2_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_1_addend_smaller_qr_3_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_1_addend_larger_qr_3_lpi_1_dfm_mx0) + 50'b1;
  assign inp_lookup_3_FpAdd_8U_23U_1_else_2_acc_nl = nl_inp_lookup_3_FpAdd_8U_23U_1_else_2_acc_nl[49:0];
  assign nand_581_nl = ~(main_stage_v_4 & (chn_inp_in_crt_sva_4_739_736_1[2]) & (cfg_precision_1_sva_st_81==2'b10));
  assign mux_499_nl = MUX_s_1_2_2(or_tmp_899, (nand_581_nl), or_11_cse);
  assign and_4130_nl = inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_8_5_1 & (inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_8_4_0_1[4]);
  assign and_4131_nl = FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_9_1
      & FpAdd_8U_23U_o_sign_3_lpi_1_dfm_9;
  assign nor_1876_nl = ~((FpMul_6U_10U_1_o_expo_3_lpi_1_dfm[5:4]!=2'b11) | FpMul_6U_10U_1_lor_8_lpi_1_dfm_6);
  assign mux_2088_nl = MUX_s_1_2_2((nor_1876_nl), (and_4131_nl), IsNaN_6U_10U_5_land_3_lpi_1_dfm_6);
  assign mux_2089_nl = MUX_s_1_2_2((mux_2088_nl), (and_4130_nl), IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_16);
  assign nor_1875_nl = ~((~ FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_4) | IsNaN_6U_10U_5_land_3_lpi_1_dfm_6);
  assign or_5992_nl = (inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_8_5_1 & (inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_8_4_0_1[4])
      & (FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_3_0_mx1w1==4'b1111)) | or_tmp_4698;
  assign or_5993_nl = (FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_9_1
      & FpAdd_8U_23U_o_sign_3_lpi_1_dfm_9 & (FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_3_0_mx1w1==4'b1111))
      | or_tmp_4698;
  assign or_5994_nl = ((FpMul_6U_10U_1_o_expo_3_lpi_1_dfm[5:4]==2'b11) & (~ FpMul_6U_10U_1_lor_8_lpi_1_dfm_6)
      & (FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_3_0_mx1w1==4'b1111)) | or_tmp_4698;
  assign mux_2091_nl = MUX_s_1_2_2((or_5994_nl), (or_5993_nl), IsNaN_6U_10U_5_land_3_lpi_1_dfm_6);
  assign mux_2092_nl = MUX_s_1_2_2((mux_2091_nl), (or_5992_nl), IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_16);
  assign mux_2093_nl = MUX_s_1_2_2(or_tmp_4698, (mux_2092_nl), or_5985_cse);
  assign mux_2094_nl = MUX_s_1_2_2((mux_2093_nl), (nor_1875_nl), chn_inp_in_crt_sva_4_739_736_1[2]);
  assign and_4156_nl = ((FpMul_6U_10U_1_o_expo_3_lpi_1_dfm[5:4]!=2'b11) | FpMul_6U_10U_1_lor_8_lpi_1_dfm_6)
      & or_tmp_4703;
  assign mux_2095_nl = MUX_s_1_2_2((and_4156_nl), and_4155_cse, IsNaN_6U_10U_5_land_3_lpi_1_dfm_6);
  assign mux_2096_nl = MUX_s_1_2_2((mux_2095_nl), and_4154_cse, IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_16);
  assign mux_2097_nl = MUX_s_1_2_2(or_tmp_4703, (mux_2096_nl), or_5985_cse);
  assign mux_2098_nl = MUX_s_1_2_2(or_tmp_4703, (mux_2097_nl), and_4126_cse);
  assign and_4123_nl = (~((FpMul_6U_10U_1_o_expo_3_lpi_1_dfm[5:4]==2'b11))) & or_tmp_4703;
  assign mux_2099_nl = MUX_s_1_2_2((and_4123_nl), or_tmp_4703, FpMul_6U_10U_1_lor_8_lpi_1_dfm_6);
  assign mux_2100_nl = MUX_s_1_2_2((mux_2099_nl), and_4155_cse, IsNaN_6U_10U_5_land_3_lpi_1_dfm_6);
  assign mux_2101_nl = MUX_s_1_2_2((mux_2100_nl), and_4154_cse, IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_16);
  assign mux_2102_nl = MUX_s_1_2_2(or_tmp_4703, (mux_2101_nl), or_5985_cse);
  assign mux_2103_nl = MUX_s_1_2_2(or_tmp_4703, (mux_2102_nl), and_4126_cse);
  assign and_3319_nl = main_stage_v_4 & (~((~((chn_inp_in_crt_sva_4_739_736_1[3])
      | (~ FpAdd_6U_10U_1_is_a_greater_acc_3_itm_6_1))) | (cfg_precision_1_sva_st_81!=2'b10)));
  assign nor_1578_nl = ~((~((chn_inp_in_crt_sva_5_739_736_1[3]) | (~ chn_inp_in_crt_sva_5_459_1)))
      | (cfg_precision_1_sva_st_82[0]) | not_tmp_374);
  assign mux_510_nl = MUX_s_1_2_2((nor_1578_nl), (and_3319_nl), or_11_cse);
  assign nl_inp_lookup_4_FpAdd_8U_23U_1_if_2_acc_nl = conv_u2u_49_50(FpAdd_8U_23U_1_addend_larger_qr_lpi_1_dfm_mx0)
      + conv_u2u_49_50(FpAdd_8U_23U_1_addend_smaller_qr_lpi_1_dfm_mx0);
  assign inp_lookup_4_FpAdd_8U_23U_1_if_2_acc_nl = nl_inp_lookup_4_FpAdd_8U_23U_1_if_2_acc_nl[49:0];
  assign nl_inp_lookup_4_FpAdd_8U_23U_1_else_2_acc_nl = ({1'b1 , (~ FpAdd_8U_23U_1_addend_smaller_qr_lpi_1_dfm_mx0)})
      + conv_u2u_49_50(FpAdd_8U_23U_1_addend_larger_qr_lpi_1_dfm_mx0) + 50'b1;
  assign inp_lookup_4_FpAdd_8U_23U_1_else_2_acc_nl = nl_inp_lookup_4_FpAdd_8U_23U_1_else_2_acc_nl[49:0];
  assign mux_513_nl = MUX_s_1_2_2(or_tmp_945, nand_579_cse, or_11_cse);
  assign or_6170_nl = (IsNaN_8U_23U_3_land_1_lpi_1_dfm_6 & (chn_inp_in_crt_sva_5_739_736_1[0])
      & or_11_cse) | mux_1901_tmp;
  assign and_1172_nl = (~ IsNaN_8U_23U_3_land_1_lpi_1_dfm_6) & (chn_inp_in_crt_sva_5_739_736_1[0])
      & or_11_cse & (~ mux_1901_tmp);
  assign or_6171_nl = (IsNaN_8U_23U_3_land_2_lpi_1_dfm_6 & (chn_inp_in_crt_sva_5_739_736_1[1])
      & or_11_cse) | mux_1902_tmp;
  assign and_1183_nl = (~ IsNaN_8U_23U_3_land_2_lpi_1_dfm_6) & (chn_inp_in_crt_sva_5_739_736_1[1])
      & or_11_cse & (~ mux_1902_tmp);
  assign nor_1910_nl = ~(and_dcpl_712 | mux_1903_tmp);
  assign and_4169_nl = and_dcpl_712 & (~ mux_1903_tmp);
  assign or_6172_nl = (IsNaN_8U_23U_3_land_lpi_1_dfm_5 & (chn_inp_in_crt_sva_5_739_736_1[3])
      & or_11_cse) | mux_1904_tmp;
  assign and_1201_nl = (~ IsNaN_8U_23U_3_land_lpi_1_dfm_5) & (chn_inp_in_crt_sva_5_739_736_1[3])
      & or_11_cse & (~ mux_1904_tmp);
  assign nor_1572_nl = ~(IsNaN_6U_10U_8_land_1_lpi_1_dfm_st_3 | (cfg_precision_1_sva_st_83!=2'b10)
      | (~((chn_inp_in_crt_sva_6_739_736_1[0]) & main_stage_v_6 & (IsNaN_8U_23U_3_land_1_lpi_1_dfm_7
      | (~(FpAdd_6U_10U_1_is_a_greater_lor_1_lpi_1_dfm_5 | (inp_lookup_1_FpMantRNE_49U_24U_1_else_and_svs_2
      & (~(FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_7_4_1 & FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_7_5_1)))))))));
  assign nor_1574_nl = ~((~ (chn_inp_in_crt_sva_5_739_736_1[0])) | IsNaN_8U_23U_2_land_1_lpi_1_dfm_9
      | (cfg_precision_1_sva_st_82[0]) | not_tmp_374);
  assign nor_1575_nl = ~(nor_126_cse | (~((~ inp_lookup_1_FpMantRNE_49U_24U_1_else_and_tmp)
      | inp_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_1_itm_7_1)) | (~ (chn_inp_in_crt_sva_5_739_736_1[0]))
      | IsNaN_8U_23U_2_land_1_lpi_1_dfm_9 | (cfg_precision_1_sva_st_82[0]) | not_tmp_374);
  assign mux_514_nl = MUX_s_1_2_2((nor_1575_nl), (nor_1574_nl), IsNaN_8U_23U_3_land_1_lpi_1_dfm_6);
  assign mux_515_nl = MUX_s_1_2_2((mux_514_nl), (nor_1572_nl), nor_1896_cse);
  assign nor_1568_nl = ~((chn_inp_in_crt_sva_5_739_736_1[0]) | mux_tmp_441);
  assign nor_1569_nl = ~((~ IsNaN_8U_23U_3_land_1_lpi_1_dfm_7) | (cfg_precision_1_sva_st_83!=2'b10)
      | (chn_inp_in_crt_sva_6_739_736_1[0]) | (~ main_stage_v_6));
  assign nor_1570_nl = ~(IsNaN_8U_23U_3_land_1_lpi_1_dfm_7 | (cfg_precision_1_sva_st_83!=2'b10)
      | (chn_inp_in_crt_sva_6_739_736_1[0]) | (~ main_stage_v_6));
  assign mux_520_nl = MUX_s_1_2_2((nor_1570_nl), (nor_1569_nl), IsZero_6U_10U_1_IsZero_6U_10U_1_and_itm_11);
  assign mux_521_nl = MUX_s_1_2_2((mux_520_nl), (nor_1568_nl), or_11_cse);
  assign mux_523_nl = MUX_s_1_2_2(or_tmp_962, or_tmp_959, IsNaN_8U_23U_3_land_1_lpi_1_dfm_7);
  assign mux_524_nl = MUX_s_1_2_2(or_tmp_959, or_tmp_962, IsNaN_8U_23U_3_land_1_lpi_1_dfm_7);
  assign mux_525_nl = MUX_s_1_2_2((mux_524_nl), (mux_523_nl), IsZero_6U_10U_1_IsZero_6U_10U_1_and_itm_11);
  assign mux_526_nl = MUX_s_1_2_2((mux_525_nl), mux_tmp_444, or_11_cse);
  assign nor_1562_nl = ~((~((FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_7_4_1 & FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_7_5_1
      & (~ FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_5)) | IsNaN_8U_23U_3_land_2_lpi_1_dfm_7))
      | IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_4 | (cfg_precision_1_sva_st_83[0]) | not_tmp_428);
  assign nor_1564_nl = ~((~((~ FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_5) | IsNaN_8U_23U_3_land_2_lpi_1_dfm_7))
      | IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_4 | (cfg_precision_1_sva_st_83[0]) | not_tmp_428);
  assign mux_527_nl = MUX_s_1_2_2((nor_1564_nl), (nor_1562_nl), inp_lookup_2_FpMantRNE_49U_24U_1_else_and_svs_2);
  assign nor_1567_nl = ~((FpAdd_8U_23U_1_int_mant_p1_2_sva_3[49]) | (~ or_2663_cse));
  assign mux_528_nl = MUX_s_1_2_2((nor_1567_nl), or_2663_cse, inp_lookup_2_FpAdd_8U_23U_1_if_3_if_acc_1_itm_7_1);
  assign nor_1566_nl = ~((~ (chn_inp_in_crt_sva_5_739_736_1[1])) | IsNaN_8U_23U_2_land_2_lpi_1_dfm_9
      | (cfg_precision_1_sva_st_82!=2'b10) | (~(main_stage_v_5 & (IsNaN_8U_23U_3_land_2_lpi_1_dfm_6
      | (mux_528_nl)))));
  assign mux_529_nl = MUX_s_1_2_2((nor_1566_nl), (mux_527_nl), nor_1896_cse);
  assign nor_1559_nl = ~((chn_inp_in_crt_sva_5_739_736_1[1]) | mux_tmp_454);
  assign nor_1560_nl = ~((~ IsNaN_8U_23U_3_land_2_lpi_1_dfm_7) | (cfg_precision_1_sva_st_83!=2'b10)
      | (chn_inp_in_crt_sva_6_739_736_1[1]) | (~ main_stage_v_6));
  assign nor_1561_nl = ~(IsNaN_8U_23U_3_land_2_lpi_1_dfm_7 | (cfg_precision_1_sva_st_83!=2'b10)
      | (chn_inp_in_crt_sva_6_739_736_1[1]) | (~ main_stage_v_6));
  assign mux_533_nl = MUX_s_1_2_2((nor_1561_nl), (nor_1560_nl), IsZero_6U_10U_1_IsZero_6U_10U_1_and_1_itm_9);
  assign mux_534_nl = MUX_s_1_2_2((mux_533_nl), (nor_1559_nl), or_11_cse);
  assign mux_536_nl = MUX_s_1_2_2(or_tmp_992, or_tmp_990, IsNaN_8U_23U_3_land_2_lpi_1_dfm_7);
  assign mux_537_nl = MUX_s_1_2_2(or_tmp_990, or_tmp_992, IsNaN_8U_23U_3_land_2_lpi_1_dfm_7);
  assign mux_538_nl = MUX_s_1_2_2((mux_537_nl), (mux_536_nl), IsZero_6U_10U_1_IsZero_6U_10U_1_and_1_itm_9);
  assign mux_539_nl = MUX_s_1_2_2((mux_538_nl), mux_tmp_457, or_11_cse);
  assign nor_1557_nl = ~((chn_inp_in_crt_sva_5_739_736_1[2]) | (cfg_precision_1_sva_st_82!=2'b10)
      | not_tmp_442);
  assign nor_1558_nl = ~((chn_inp_in_crt_sva_6_739_736_1[2]) | mux_tmp_465);
  assign mux_544_nl = MUX_s_1_2_2((nor_1558_nl), (nor_1557_nl), or_11_cse);
  assign mux_546_nl = MUX_s_1_2_2(mux_tmp_465, or_tmp_959, chn_inp_in_crt_sva_6_739_736_1[2]);
  assign mux_547_nl = MUX_s_1_2_2((mux_546_nl), mux_tmp_467, or_11_cse);
  assign nor_1552_nl = ~(IsNaN_6U_10U_8_land_lpi_1_dfm_st_4 | (~ (chn_inp_in_crt_sva_6_739_736_1[3]))
      | (cfg_precision_1_sva_st_83!=2'b10) | (~ main_stage_v_6));
  assign nor_1553_nl = ~(FpAdd_6U_10U_1_is_a_greater_lor_lpi_1_dfm_5 | ((~(FpMul_6U_10U_1_o_expo_lpi_1_dfm_7_4_1
      & FpMul_6U_10U_1_o_expo_lpi_1_dfm_7_5_1)) & inp_lookup_4_FpMantRNE_49U_24U_1_else_and_svs_2)
      | IsNaN_6U_10U_8_land_lpi_1_dfm_st_4 | (~ (chn_inp_in_crt_sva_6_739_736_1[3]))
      | (cfg_precision_1_sva_st_83!=2'b10) | (~ main_stage_v_6));
  assign mux_548_nl = MUX_s_1_2_2((nor_1553_nl), (nor_1552_nl), IsNaN_8U_23U_3_land_lpi_1_dfm_6);
  assign nor_1554_nl = ~((~ (chn_inp_in_crt_sva_5_739_736_1[3])) | IsNaN_8U_23U_2_land_lpi_1_dfm_9
      | (cfg_precision_1_sva_st_82[0]) | not_tmp_374);
  assign nor_1555_nl = ~(nor_136_cse | (~((~ inp_lookup_4_FpMantRNE_49U_24U_1_else_and_tmp)
      | inp_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_1_itm_7_1)) | (~ (chn_inp_in_crt_sva_5_739_736_1[3]))
      | IsNaN_8U_23U_2_land_lpi_1_dfm_9 | (cfg_precision_1_sva_st_82[0]) | not_tmp_374);
  assign mux_549_nl = MUX_s_1_2_2((nor_1555_nl), (nor_1554_nl), IsNaN_8U_23U_3_land_lpi_1_dfm_5);
  assign mux_550_nl = MUX_s_1_2_2((mux_549_nl), (mux_548_nl), nor_1896_cse);
  assign nor_1549_nl = ~((chn_inp_in_crt_sva_5_739_736_1[3]) | mux_tmp_475);
  assign nor_1550_nl = ~((~ IsNaN_8U_23U_3_land_lpi_1_dfm_6) | (chn_inp_in_crt_sva_6_739_736_1[3])
      | (cfg_precision_1_sva_st_83!=2'b10) | (~ main_stage_v_6));
  assign nor_1551_nl = ~(IsNaN_8U_23U_3_land_lpi_1_dfm_6 | (chn_inp_in_crt_sva_6_739_736_1[3])
      | (cfg_precision_1_sva_st_83!=2'b10) | (~ main_stage_v_6));
  assign mux_554_nl = MUX_s_1_2_2((nor_1551_nl), (nor_1550_nl), IsZero_6U_10U_1_IsZero_6U_10U_1_and_3_itm_9);
  assign mux_555_nl = MUX_s_1_2_2((mux_554_nl), (nor_1549_nl), or_11_cse);
  assign or_1054_nl = (~(IsNaN_8U_23U_3_land_lpi_1_dfm_6 | (chn_inp_in_crt_sva_6_739_736_1[3])))
      | (cfg_precision_1_sva_st_83!=2'b10) | (~ main_stage_v_6);
  assign or_1057_nl = (~((~ IsNaN_8U_23U_3_land_lpi_1_dfm_6) | (chn_inp_in_crt_sva_6_739_736_1[3])))
      | (cfg_precision_1_sva_st_83!=2'b10) | (~ main_stage_v_6);
  assign mux_557_nl = MUX_s_1_2_2((or_1057_nl), (or_1054_nl), IsZero_6U_10U_1_IsZero_6U_10U_1_and_3_itm_9);
  assign mux_558_nl = MUX_s_1_2_2((mux_557_nl), mux_tmp_478, or_11_cse);
  assign and_4221_nl = (~ IsNaN_8U_23U_3_land_1_lpi_1_dfm_7) & and_1211_rgt;
  assign and_3314_nl = (cfg_precision_1_sva_st_83==2'b10) & (chn_inp_in_crt_sva_6_739_736_1[0])
      & main_stage_v_6 & (~(or_tmp_1060 & (inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7
      | (~ inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8))));
  assign nor_1545_nl = ~(inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2
      | (~ inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2)
      | (~ inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_2)
      | inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
      | (~ (chn_inp_in_crt_sva_7_739_736_1[0])) | (cfg_precision_1_sva_st_84!=2'b10)
      | (~ main_stage_v_7));
  assign mux_560_nl = MUX_s_1_2_2(nor_1546_cse, (nor_1545_nl), inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2);
  assign and_3315_nl = (chn_inp_in_crt_sva_7_739_736_1[0]) & (cfg_precision_1_sva_st_84==2'b10)
      & main_stage_v_7;
  assign mux_561_nl = MUX_s_1_2_2((and_3315_nl), (mux_560_nl), FpAdd_6U_10U_1_or_12_cse);
  assign mux_562_nl = MUX_s_1_2_2((mux_561_nl), (and_3314_nl), or_11_cse);
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_1_sva_2 = conv_u2u_4_5({FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_2_sva_mx0w0
      , (~ (FpAdd_8U_23U_1_o_expo_1_lpi_1_dfm_7_mx0w0[0]))}) + 5'b1101;
  assign nor_1543_nl = ~(inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8
      | inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7 | (~ inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8)
      | (cfg_precision_1_sva_st_83!=2'b10) | not_tmp_424);
  assign nor_1544_nl = ~((~ (chn_inp_in_crt_sva_7_739_736_1[0])) | inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2
      | (~ inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2)
      | inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
      | (cfg_precision_1_sva_st_84!=2'b10) | (~ main_stage_v_7));
  assign mux_563_nl = MUX_s_1_2_2((nor_1544_nl), (nor_1543_nl), or_11_cse);
  assign nor_1540_nl = ~(inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7
      | (~ inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8) | (cfg_precision_1_sva_st_83!=2'b10)
      | not_tmp_424);
  assign mux_565_nl = MUX_s_1_2_2(nor_1546_cse, (nor_1540_nl), or_11_cse);
  assign nor_1536_nl = ~(inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8 |
      (~ nor_tmp_139));
  assign mux_568_nl = MUX_s_1_2_2((nor_1536_nl), nor_tmp_139, inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7);
  assign nor_1535_nl = ~((~ main_stage_v_6) | (cfg_precision_1_sva_st_83!=2'b10)
      | (mux_568_nl));
  assign nor_1537_nl = ~((((~((~ inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2)
      | inp_lookup_1_FpMantRNE_24U_11U_else_and_svs)) | (~ inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2)
      | inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs)
      & (chn_inp_in_crt_sva_7_739_736_1[0]) & inp_lookup_1_FpMantRNE_24U_11U_else_and_svs_2)
      | (~ main_stage_v_7) | (cfg_precision_1_sva_st_84!=2'b10));
  assign mux_569_nl = MUX_s_1_2_2((nor_1537_nl), (nor_1535_nl), or_11_cse);
  assign or_1102_nl = (chn_inp_in_crt_sva_7_739_736_1[0]) | (cfg_precision_1_sva_st_84!=2'b10)
      | (~ main_stage_v_7);
  assign mux_570_nl = MUX_s_1_2_2((or_1102_nl), or_tmp_1098, or_11_cse);
  assign FpNormalize_6U_23U_1_if_or_nl = (FpAdd_6U_10U_1_int_mant_p1_1_lpi_1_dfm_mx0[22:0]!=23'b00000000000000000000000);
  assign FpAdd_6U_10U_1_mux_2_nl = MUX_s_1_2_2((FpAdd_6U_10U_1_int_mant_p1_1_sva_1[23]),
      (FpAdd_6U_10U_1_int_mant_p1_1_sva[23]), IsNaN_8U_23U_3_land_1_lpi_1_dfm_7);
  assign mux_571_nl = MUX_s_1_2_2(or_tmp_959, or_tmp_962, FpAdd_6U_10U_1_mux_2_nl);
  assign or_1106_nl = (~((~ chn_inp_in_crt_sva_7_411_1) | (chn_inp_in_crt_sva_7_739_736_1[0])))
      | (cfg_precision_1_sva_st_84!=2'b10) | (~ main_stage_v_7);
  assign mux_572_nl = MUX_s_1_2_2((or_1106_nl), (mux_571_nl), or_11_cse);
  assign and_4220_nl = (~ IsNaN_8U_23U_3_land_2_lpi_1_dfm_7) & and_1223_rgt;
  assign nor_1530_nl = ~((cfg_precision_1_sva_st_83[0]) | (~((cfg_precision_1_sva_st_83[1])
      & (chn_inp_in_crt_sva_6_739_736_1[1]) & main_stage_v_6 & (IsNaN_8U_23U_4_IsNaN_8U_23U_4_nor_1_tmp
      | (~(inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7 | (~ inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8)))))));
  assign and_3387_nl = (chn_inp_in_crt_sva_7_739_736_1[1]) & main_stage_v_7 & (cfg_precision_1_sva_st_84==2'b10);
  assign and_3309_nl = (~(inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
      | (~ inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2)))
      & (~((inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2
      | (~ inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2)
      | (~ IsNaN_6U_10U_9_land_2_lpi_1_dfm_8)) & inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2))
      & (chn_inp_in_crt_sva_7_739_736_1[1]) & main_stage_v_7 & (cfg_precision_1_sva_st_84==2'b10);
  assign mux_574_nl = MUX_s_1_2_2((and_3309_nl), (and_3387_nl), IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_5);
  assign mux_575_nl = MUX_s_1_2_2((mux_574_nl), (nor_1530_nl), or_11_cse);
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_2_sva_2 = conv_u2u_4_5({FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_3_sva_mx0w0
      , (~ (FpAdd_8U_23U_1_o_expo_2_lpi_1_dfm_7[0]))}) + 5'b1101;
  assign nor_1528_nl = ~(inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8
      | inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7 | (~ inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8)
      | (cfg_precision_1_sva_st_83[0]) | not_tmp_428);
  assign nor_1529_nl = ~(inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2
      | inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
      | (~ inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2)
      | (cfg_precision_1_sva_st_84[0]) | (~ and_dcpl_21));
  assign mux_576_nl = MUX_s_1_2_2((nor_1529_nl), (nor_1528_nl), or_11_cse);
  assign nor_1524_nl = ~(inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7
      | (~ inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8) | (cfg_precision_1_sva_st_83[0])
      | not_tmp_428);
  assign nor_1525_nl = ~(inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
      | (~ inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2)
      | (cfg_precision_1_sva_st_84[0]) | (~ and_dcpl_21));
  assign mux_578_nl = MUX_s_1_2_2((nor_1525_nl), (nor_1524_nl), or_11_cse);
  assign nor_1519_nl = ~(inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8 |
      (~ nor_tmp_146));
  assign mux_580_nl = MUX_s_1_2_2((nor_1519_nl), nor_tmp_146, inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7);
  assign nor_1518_nl = ~((~ main_stage_v_6) | (cfg_precision_1_sva_st_83!=2'b10)
      | (mux_580_nl));
  assign nor_1520_nl = ~((((~((~ inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2)
      | inp_lookup_2_FpMantRNE_24U_11U_else_and_svs)) | (~ inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2)
      | inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs)
      & (chn_inp_in_crt_sva_7_739_736_1[1]) & inp_lookup_2_FpMantRNE_24U_11U_else_and_svs_2)
      | (~ main_stage_v_7) | (cfg_precision_1_sva_st_84!=2'b10));
  assign mux_581_nl = MUX_s_1_2_2((nor_1520_nl), (nor_1518_nl), or_11_cse);
  assign or_1147_nl = (cfg_precision_1_sva_st_84!=2'b10) | (chn_inp_in_crt_sva_7_739_736_1[1])
      | (~ main_stage_v_7);
  assign mux_582_nl = MUX_s_1_2_2((or_1147_nl), or_tmp_1143, or_11_cse);
  assign FpNormalize_6U_23U_1_if_or_1_nl = (FpAdd_6U_10U_1_int_mant_p1_2_lpi_1_dfm_mx0[22:0]!=23'b00000000000000000000000);
  assign FpAdd_6U_10U_1_mux_18_nl = MUX_s_1_2_2((FpAdd_6U_10U_1_int_mant_p1_2_sva_1[23]),
      (FpAdd_6U_10U_1_int_mant_p1_2_sva[23]), IsNaN_8U_23U_3_land_2_lpi_1_dfm_7);
  assign mux_583_nl = MUX_s_1_2_2(or_tmp_990, or_tmp_992, FpAdd_6U_10U_1_mux_18_nl);
  assign mux_584_nl = MUX_s_1_2_2(or_tmp_1147, or_tmp_1106, chn_inp_in_crt_sva_7_427_1);
  assign mux_585_nl = MUX_s_1_2_2((mux_584_nl), (mux_583_nl), or_11_cse);
  assign nor_1514_nl = ~((~ (chn_inp_in_crt_sva_6_739_736_1[2])) | (cfg_precision_1_sva_st_83!=2'b10)
      | (~(main_stage_v_6 & (IsNaN_8U_23U_4_IsNaN_8U_23U_4_nor_2_tmp | (~(inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7
      | (~ inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8)))))));
  assign and_3307_nl = main_stage_v_7 & (chn_inp_in_crt_sva_7_739_736_1[2]) & (cfg_precision_1_sva_st_84==2'b10);
  assign nor_1516_nl = ~((~ inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2)
      | inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2
      | (~ IsNaN_6U_10U_9_land_3_lpi_1_dfm_8) | inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
      | (~ main_stage_v_7) | (~ (chn_inp_in_crt_sva_7_739_736_1[2])) | (cfg_precision_1_sva_st_84!=2'b10));
  assign mux_588_nl = MUX_s_1_2_2(nor_1517_cse, (nor_1516_nl), inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2);
  assign mux_589_nl = MUX_s_1_2_2((mux_588_nl), (and_3307_nl), IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_5);
  assign mux_590_nl = MUX_s_1_2_2((mux_589_nl), (nor_1514_nl), or_11_cse);
  assign nor_1512_nl = ~(inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7
      | (~ inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8) | (~ (chn_inp_in_crt_sva_6_739_736_1[2]))
      | (cfg_precision_1_sva_st_83!=2'b10) | (~ main_stage_v_6));
  assign mux_592_nl = MUX_s_1_2_2(nor_1517_cse, (nor_1512_nl), or_11_cse);
  assign or_1179_nl = ((inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7
      | (~ inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8)) & inp_lookup_3_FpMantRNE_24U_11U_else_and_svs
      & (chn_inp_in_crt_sva_6_739_736_1[2])) | (cfg_precision_1_sva_st_83!=2'b10)
      | (~ main_stage_v_6);
  assign or_1182_nl = (((~((~ inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2)
      | inp_lookup_3_FpMantRNE_24U_11U_else_and_svs)) | inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
      | (~ inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2))
      & (chn_inp_in_crt_sva_7_739_736_1[2])) | (cfg_precision_1_sva_st_84!=2'b10)
      | (~ main_stage_v_7);
  assign mux_594_nl = MUX_s_1_2_2(or_tmp_1182, (or_1182_nl), inp_lookup_3_FpMantRNE_24U_11U_else_and_svs_2);
  assign mux_595_nl = MUX_s_1_2_2((mux_594_nl), (or_1179_nl), or_11_cse);
  assign or_1189_nl = (chn_inp_in_crt_sva_7_739_736_1[2]) | (cfg_precision_1_sva_st_84!=2'b10)
      | (~ main_stage_v_7);
  assign mux_596_nl = MUX_s_1_2_2((or_1189_nl), or_tmp_1185, or_11_cse);
  assign FpNormalize_6U_23U_1_if_or_2_nl = (FpAdd_6U_10U_1_int_mant_p1_3_lpi_1_dfm_mx0[22:0]!=23'b00000000000000000000000);
  assign FpAdd_6U_10U_1_mux_34_nl = MUX_s_1_2_2((FpAdd_6U_10U_1_int_mant_p1_3_sva_1[23]),
      (FpAdd_6U_10U_1_int_mant_p1_3_sva[23]), IsNaN_8U_23U_3_land_3_lpi_1_dfm_7);
  assign nor_1507_nl = ~((~((~ (FpAdd_6U_10U_1_mux_34_nl)) | (chn_inp_in_crt_sva_6_739_736_1[2])))
      | (cfg_precision_1_sva_st_83!=2'b10) | (~ main_stage_v_6));
  assign nor_1509_nl = ~((~((~ chn_inp_in_crt_sva_7_443_1) | (chn_inp_in_crt_sva_7_739_736_1[2])))
      | (cfg_precision_1_sva_st_84!=2'b10) | (~ main_stage_v_7));
  assign mux_597_nl = MUX_s_1_2_2((nor_1509_nl), (nor_1507_nl), or_11_cse);
  assign and_4219_nl = (~ IsNaN_8U_23U_3_land_lpi_1_dfm_6) & and_1247_rgt;
  assign nor_1504_nl = ~((~ (chn_inp_in_crt_sva_6_739_736_1[3])) | (cfg_precision_1_sva_st_83!=2'b10)
      | (~(main_stage_v_6 & (IsNaN_8U_23U_4_IsNaN_8U_23U_4_nor_3_tmp | (~(inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7
      | (~ inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8)))))));
  assign and_3386_nl = (chn_inp_in_crt_sva_7_739_736_1[3]) & (cfg_precision_1_sva_st_84==2'b10)
      & main_stage_v_7;
  assign and_3300_nl = (~(inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
      | (~ inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2)))
      & (~((inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2
      | (~ inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2)
      | (~ IsNaN_6U_10U_9_land_lpi_1_dfm_8)) & inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2))
      & (chn_inp_in_crt_sva_7_739_736_1[3]) & (cfg_precision_1_sva_st_84==2'b10)
      & main_stage_v_7;
  assign mux_600_nl = MUX_s_1_2_2((and_3300_nl), (and_3386_nl), IsNaN_6U_10U_8_land_lpi_1_dfm_st_5);
  assign mux_601_nl = MUX_s_1_2_2((mux_600_nl), (nor_1504_nl), or_11_cse);
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva_2 = conv_u2u_4_5({FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_1_sva_mx0w0
      , (~ (FpAdd_8U_23U_1_o_expo_lpi_1_dfm_7[0]))}) + 5'b1101;
  assign nor_1502_nl = ~(inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8
      | inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7 | (~ inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8)
      | (~ (chn_inp_in_crt_sva_6_739_736_1[3])) | (cfg_precision_1_sva_st_83!=2'b10)
      | (~ main_stage_v_6));
  assign nor_1503_nl = ~(inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2
      | (~ (chn_inp_in_crt_sva_7_739_736_1[3])) | inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
      | (~ inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2)
      | (cfg_precision_1_sva_st_84!=2'b10) | (~ main_stage_v_7));
  assign mux_602_nl = MUX_s_1_2_2((nor_1503_nl), (nor_1502_nl), or_11_cse);
  assign nor_1500_nl = ~(inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7
      | (~ inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8) | (~ (chn_inp_in_crt_sva_6_739_736_1[3]))
      | (cfg_precision_1_sva_st_83!=2'b10) | (~ main_stage_v_6));
  assign nor_1501_nl = ~((~ (chn_inp_in_crt_sva_7_739_736_1[3])) | inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
      | (~ inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2)
      | (cfg_precision_1_sva_st_84!=2'b10) | (~ main_stage_v_7));
  assign mux_604_nl = MUX_s_1_2_2((nor_1501_nl), (nor_1500_nl), or_11_cse);
  assign or_1232_nl = ((inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7
      | (~ inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8)) & inp_lookup_4_FpMantRNE_24U_11U_else_and_svs
      & (chn_inp_in_crt_sva_6_739_736_1[3])) | (cfg_precision_1_sva_st_83!=2'b10)
      | (~ main_stage_v_6);
  assign or_1236_nl = inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
      | (~ inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2)
      | (cfg_precision_1_sva_st_84!=2'b10) | (~ main_stage_v_7);
  assign mux_606_nl = MUX_s_1_2_2(or_tmp_1182, (or_1236_nl), chn_inp_in_crt_sva_7_739_736_1[3]);
  assign nor_158_nl = ~(inp_lookup_4_FpMantRNE_24U_11U_else_and_svs | (~ inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2));
  assign mux_607_nl = MUX_s_1_2_2((mux_606_nl), or_tmp_1232, nor_158_nl);
  assign mux_608_nl = MUX_s_1_2_2(or_tmp_1182, (mux_607_nl), inp_lookup_4_FpMantRNE_24U_11U_else_and_svs_2);
  assign mux_609_nl = MUX_s_1_2_2((mux_608_nl), (or_1232_nl), or_11_cse);
  assign mux_610_nl = MUX_s_1_2_2(or_tmp_1232, or_tmp_1239, or_11_cse);
  assign FpNormalize_6U_23U_1_if_or_3_nl = (FpAdd_6U_10U_1_int_mant_p1_lpi_1_dfm_mx0[22:0]!=23'b00000000000000000000000);
  assign FpAdd_6U_10U_1_mux_50_nl = MUX_s_1_2_2((FpAdd_6U_10U_1_int_mant_p1_sva_1[23]),
      (FpAdd_6U_10U_1_int_mant_p1_sva[23]), IsNaN_8U_23U_3_land_lpi_1_dfm_6);
  assign nor_1496_nl = ~((~((~ (FpAdd_6U_10U_1_mux_50_nl)) | (chn_inp_in_crt_sva_6_739_736_1[3])))
      | (cfg_precision_1_sva_st_83!=2'b10) | (~ main_stage_v_6));
  assign nor_1498_nl = ~((~((~ chn_inp_in_crt_sva_7_459_1) | (chn_inp_in_crt_sva_7_739_736_1[3])))
      | (cfg_precision_1_sva_st_84!=2'b10) | (~ main_stage_v_7));
  assign mux_611_nl = MUX_s_1_2_2((nor_1498_nl), (nor_1496_nl), or_11_cse);
  assign inp_lookup_1_IsInf_6U_23U_1_IsInf_6U_23U_1_and_nl = FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_5_mx0w0
      & FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_4_mx0w0 & (FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_3_0_mx0w0==4'b1111);
  assign nor_1489_nl = ~((~ (chn_inp_in_crt_sva_7_739_736_1[0])) | FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_tmp
      | (cfg_precision_1_sva_st_84!=2'b10) | (~ main_stage_v_7));
  assign mux_620_nl = MUX_s_1_2_2(nor_1490_cse, (nor_1489_nl), or_11_cse);
  assign inp_lookup_1_FpMul_6U_10U_xor_1_nl = FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_8_4_1
      ^ chn_inp_in_crt_sva_7_411_1;
  assign inp_lookup_2_IsInf_6U_23U_1_IsInf_6U_23U_1_and_nl = FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_5_mx0w0
      & FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_4_mx0w0 & (FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_3_0_mx0w0==4'b1111);
  assign nor_1480_nl = ~(FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_2_tmp | (cfg_precision_1_sva_st_84[0])
      | (~ and_dcpl_21));
  assign nor_1481_nl = ~(reg_FpMul_6U_10U_lor_4_lpi_1_dfm_3_cse | (cfg_precision_1_sva_st_85[0])
      | not_tmp_537);
  assign mux_630_nl = MUX_s_1_2_2((nor_1481_nl), (nor_1480_nl), or_11_cse);
  assign inp_lookup_2_FpMul_6U_10U_xor_1_nl = FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_8_4_1
      ^ chn_inp_in_crt_sva_7_427_1;
  assign inp_lookup_3_IsInf_6U_23U_1_IsInf_6U_23U_1_and_nl = FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_5_mx0w0
      & FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_4_mx0w0 & (FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_3_0_mx0w0==4'b1111);
  assign nor_1474_nl = ~(FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_4_tmp | (~ (chn_inp_in_crt_sva_7_739_736_1[2]))
      | (cfg_precision_1_sva_st_84!=2'b10) | (~ main_stage_v_7));
  assign nor_1475_nl = ~(reg_FpMul_6U_10U_lor_5_lpi_1_dfm_3_cse | (~ (chn_inp_in_crt_sva_8_739_736_1[2]))
      | (cfg_precision_1_sva_st_85!=2'b10) | (~ main_stage_v_8));
  assign mux_640_nl = MUX_s_1_2_2((nor_1475_nl), (nor_1474_nl), or_11_cse);
  assign inp_lookup_3_FpMul_6U_10U_xor_1_nl = FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_8_4_1
      ^ chn_inp_in_crt_sva_7_443_1;
  assign inp_lookup_4_IsInf_6U_23U_1_IsInf_6U_23U_1_and_nl = FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_5_mx0w0
      & FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_4_mx0w0 & (FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_3_0_mx0w0==4'b1111);
  assign nor_1468_nl = ~(FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_6_tmp | (~ (chn_inp_in_crt_sva_7_739_736_1[3]))
      | (cfg_precision_1_sva_st_84!=2'b10) | (~ main_stage_v_7));
  assign mux_650_nl = MUX_s_1_2_2(nor_1469_cse, (nor_1468_nl), or_11_cse);
  assign inp_lookup_4_FpMul_6U_10U_xor_1_nl = FpMul_6U_10U_1_o_expo_lpi_1_dfm_8_4_1
      ^ chn_inp_in_crt_sva_7_459_1;
  assign nl_FpMul_6U_10U_else_2_else_acc_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_13_1_1
      , FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_5_1 , FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_3_0_1})
      + 6'b100001;
  assign FpMul_6U_10U_else_2_else_acc_nl = nl_FpMul_6U_10U_else_2_else_acc_nl[5:0];
  assign nl_FpMul_6U_10U_else_2_else_ac_int_cctor_1_sva_2 = (FpMul_6U_10U_else_2_else_acc_nl)
      + ({FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_10_5_1 , FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_1_lpi_1_dfm_10_4_0_1});
  assign nor_1464_nl = ~((~ main_stage_v_8) | (~ (chn_inp_in_crt_sva_8_739_736_1[0]))
      | (cfg_precision_1_sva_st_85!=2'b10) | (~ inp_lookup_1_FpMul_6U_10U_else_2_if_acc_itm_6_1)
      | reg_FpMul_6U_10U_lor_3_lpi_1_dfm_3_cse | inp_lookup_1_FpMul_6U_10U_oelse_1_acc_itm_7_1
      | (~((~ or_tmp_1363) | (inp_lookup_1_FpMul_6U_10U_p_mant_p1_mul_tmp[21]))));
  assign nor_1465_nl = ~((~ main_stage_v_9) | (~ (chn_inp_in_crt_sva_9_739_736_1[0]))
      | (cfg_precision_1_sva_st_86!=2'b10) | FpMul_6U_10U_lor_6_lpi_1_dfm_st_2 |
      (~(inp_lookup_1_FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs
      & (inp_lookup_1_FpMul_6U_10U_else_2_else_slc_FpMul_6U_10U_p_mant_p1_21_itm_2
      | (~(or_tmp_1369 | (FpMul_6U_10U_p_mant_p1_1_sva_2[21])))))));
  assign mux_654_nl = MUX_s_1_2_2((nor_1465_nl), (nor_1464_nl), or_11_cse);
  assign nor_1912_nl = ~(inp_lookup_1_FpMul_6U_10U_oelse_1_acc_itm_7_1 | (~ inp_lookup_1_FpMul_6U_10U_else_2_if_acc_itm_6_1)
      | (~ (chn_inp_in_crt_sva_8_739_736_1[0])) | (cfg_precision_1_sva_st_85!=2'b10)
      | (~ main_stage_v_8) | reg_FpMul_6U_10U_lor_3_lpi_1_dfm_3_cse);
  assign nor_1463_nl = ~((~ (chn_inp_in_crt_sva_9_739_736_1[0])) | FpMul_6U_10U_lor_6_lpi_1_dfm_st_2
      | (~ inp_lookup_1_FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs)
      | (~ main_stage_v_9) | (cfg_precision_1_sva_st_86!=2'b10));
  assign mux_656_nl = MUX_s_1_2_2((nor_1463_nl), (nor_1912_nl), or_11_cse);
  assign nl_FpMul_6U_10U_else_2_else_acc_2_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_13_1_1
      , FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_5_1 , FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_3_0_1})
      + 6'b100001;
  assign FpMul_6U_10U_else_2_else_acc_2_nl = nl_FpMul_6U_10U_else_2_else_acc_2_nl[5:0];
  assign nl_FpMul_6U_10U_else_2_else_ac_int_cctor_2_sva_2 = (FpMul_6U_10U_else_2_else_acc_2_nl)
      + ({FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_10_5_1 , FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_2_lpi_1_dfm_10_4_0_1});
  assign nor_1454_nl = ~((~ main_stage_v_8) | (~ (chn_inp_in_crt_sva_8_739_736_1[1]))
      | (cfg_precision_1_sva_st_85!=2'b10) | (~ inp_lookup_2_FpMul_6U_10U_else_2_if_acc_itm_6_1)
      | reg_FpMul_6U_10U_lor_4_lpi_1_dfm_3_cse | inp_lookup_2_FpMul_6U_10U_oelse_1_acc_itm_7_1
      | (~((~ or_tmp_1393) | (inp_lookup_2_FpMul_6U_10U_p_mant_p1_mul_tmp[21]))));
  assign nor_1455_nl = ~((~ main_stage_v_9) | (~ (chn_inp_in_crt_sva_9_739_736_1[1]))
      | (cfg_precision_1_sva_st_100!=2'b10) | FpMul_6U_10U_lor_7_lpi_1_dfm_st_2 |
      (~(inp_lookup_2_FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs
      & (inp_lookup_2_FpMul_6U_10U_else_2_else_slc_FpMul_6U_10U_p_mant_p1_21_itm_2
      | (~(or_tmp_1399 | (FpMul_6U_10U_p_mant_p1_2_sva_2[21])))))));
  assign mux_662_nl = MUX_s_1_2_2((nor_1455_nl), (nor_1454_nl), or_11_cse);
  assign nor_1452_nl = ~((~ inp_lookup_2_FpMul_6U_10U_else_2_if_acc_itm_6_1) | reg_FpMul_6U_10U_lor_4_lpi_1_dfm_3_cse
      | inp_lookup_2_FpMul_6U_10U_oelse_1_acc_itm_7_1 | (cfg_precision_1_sva_st_85[0])
      | not_tmp_537);
  assign nor_1453_nl = ~((~ (chn_inp_in_crt_sva_9_739_736_1[1])) | (~ inp_lookup_2_FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs)
      | FpMul_6U_10U_lor_7_lpi_1_dfm_st_2 | (~ main_stage_v_9) | (cfg_precision_1_sva_st_100!=2'b10));
  assign mux_664_nl = MUX_s_1_2_2((nor_1453_nl), (nor_1452_nl), or_11_cse);
  assign nl_FpMul_6U_10U_else_2_else_acc_3_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_13_1_1
      , FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_5_1 , FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_3_0_1})
      + 6'b100001;
  assign FpMul_6U_10U_else_2_else_acc_3_nl = nl_FpMul_6U_10U_else_2_else_acc_3_nl[5:0];
  assign nl_FpMul_6U_10U_else_2_else_ac_int_cctor_3_sva_2 = (FpMul_6U_10U_else_2_else_acc_3_nl)
      + ({FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_10_5_1 , FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_3_lpi_1_dfm_10_4_0_1});
  assign nor_1446_nl = ~((~ main_stage_v_8) | (~ (chn_inp_in_crt_sva_8_739_736_1[2]))
      | (cfg_precision_1_sva_st_85!=2'b10) | (~ inp_lookup_3_FpMul_6U_10U_else_2_if_acc_itm_6_1)
      | reg_FpMul_6U_10U_lor_5_lpi_1_dfm_3_cse | inp_lookup_3_FpMul_6U_10U_oelse_1_acc_itm_7_1
      | (~((~ or_tmp_1422) | (inp_lookup_3_FpMul_6U_10U_p_mant_p1_mul_tmp[21]))));
  assign nor_1447_nl = ~((~ main_stage_v_9) | (~ (chn_inp_in_crt_sva_9_739_736_1[2]))
      | (cfg_precision_1_sva_st_112!=2'b10) | FpMul_6U_10U_lor_8_lpi_1_dfm_st_2 |
      (~(inp_lookup_3_FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs
      & (inp_lookup_3_FpMul_6U_10U_else_2_else_slc_FpMul_6U_10U_p_mant_p1_21_itm_2
      | (~(or_tmp_1428 | (FpMul_6U_10U_p_mant_p1_3_sva_2[21])))))));
  assign mux_669_nl = MUX_s_1_2_2((nor_1447_nl), (nor_1446_nl), or_11_cse);
  assign and_3284_nl = inp_lookup_3_FpMul_6U_10U_else_2_if_acc_itm_6_1 & (~(inp_lookup_3_FpMul_6U_10U_oelse_1_acc_itm_7_1
      | (~ (chn_inp_in_crt_sva_8_739_736_1[2])) | (cfg_precision_1_sva_st_85!=2'b10)
      | (~ main_stage_v_8) | reg_FpMul_6U_10U_lor_5_lpi_1_dfm_3_cse));
  assign nor_1445_nl = ~((~ (chn_inp_in_crt_sva_9_739_736_1[2])) | (~ inp_lookup_3_FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs)
      | FpMul_6U_10U_lor_8_lpi_1_dfm_st_2 | (~ main_stage_v_9) | (cfg_precision_1_sva_st_112!=2'b10));
  assign mux_671_nl = MUX_s_1_2_2((nor_1445_nl), (and_3284_nl), or_11_cse);
  assign nl_FpMul_6U_10U_else_2_else_acc_4_nl = ({FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_13_1_1
      , FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_5_1 , FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_3_0_1})
      + 6'b100001;
  assign FpMul_6U_10U_else_2_else_acc_4_nl = nl_FpMul_6U_10U_else_2_else_acc_4_nl[5:0];
  assign nl_FpMul_6U_10U_else_2_else_ac_int_cctor_sva_2 = (FpMul_6U_10U_else_2_else_acc_4_nl)
      + ({FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_10_5_1 , FpWidthDec_8U_23U_6U_10U_0U_1U_o_expo_lpi_1_dfm_10_4_0_1});
  assign nor_1441_nl = ~((~ main_stage_v_8) | (~ (chn_inp_in_crt_sva_8_739_736_1[3]))
      | (cfg_precision_1_sva_st_85!=2'b10) | (~ inp_lookup_4_FpMul_6U_10U_else_2_if_acc_itm_6_1)
      | reg_FpMul_6U_10U_lor_lpi_1_dfm_3_cse | inp_lookup_4_FpMul_6U_10U_oelse_1_acc_itm_7_1
      | (~((~ or_tmp_1448) | (inp_lookup_4_FpMul_6U_10U_p_mant_p1_mul_tmp[21]))));
  assign nor_1442_nl = ~((~ main_stage_v_9) | (~ (chn_inp_in_crt_sva_9_739_736_1[3]))
      | (cfg_precision_1_sva_st_124!=2'b10) | FpMul_6U_10U_lor_1_lpi_1_dfm_st_2 |
      (~(inp_lookup_4_FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs
      & (inp_lookup_4_FpMul_6U_10U_else_2_else_slc_FpMul_6U_10U_p_mant_p1_21_itm_2
      | (~(or_tmp_1454 | (FpMul_6U_10U_p_mant_p1_sva_2[21])))))));
  assign mux_676_nl = MUX_s_1_2_2((nor_1442_nl), (nor_1441_nl), or_11_cse);
  assign and_3282_nl = inp_lookup_4_FpMul_6U_10U_else_2_if_acc_itm_6_1 & (~(inp_lookup_4_FpMul_6U_10U_oelse_1_acc_itm_7_1
      | (~ (chn_inp_in_crt_sva_8_739_736_1[3])) | (cfg_precision_1_sva_st_85!=2'b10)
      | (~ main_stage_v_8) | reg_FpMul_6U_10U_lor_lpi_1_dfm_3_cse));
  assign nor_1440_nl = ~((~ inp_lookup_4_FpMul_6U_10U_else_2_if_slc_FpMul_6U_10U_else_2_if_acc_6_svs)
      | (~ (chn_inp_in_crt_sva_9_739_736_1[3])) | FpMul_6U_10U_lor_1_lpi_1_dfm_st_2
      | (~ main_stage_v_9) | (cfg_precision_1_sva_st_124!=2'b10));
  assign mux_678_nl = MUX_s_1_2_2((nor_1440_nl), (and_3282_nl), or_11_cse);
  assign mux_700_nl = MUX_s_1_2_2(nor_tmp_199, and_3113_cse, or_11_cse);
  assign mux_718_nl = MUX_s_1_2_2(nor_tmp_208, and_3111_cse, or_11_cse);
  assign mux_736_nl = MUX_s_1_2_2(nor_tmp_216, and_3110_cse, or_11_cse);
  assign mux_754_nl = MUX_s_1_2_2(nor_tmp_224, and_3112_cse, or_11_cse);
  assign mux_760_nl = MUX_s_1_2_2(nor_tmp_227, nor_tmp_199, or_11_cse);
  assign mux_765_nl = MUX_s_1_2_2(nor_tmp_230, nor_tmp_208, or_11_cse);
  assign mux_770_nl = MUX_s_1_2_2(nor_tmp_232, nor_tmp_216, or_11_cse);
  assign mux_775_nl = MUX_s_1_2_2(nor_tmp_234, nor_tmp_224, or_11_cse);
  assign nor_1418_nl = ~((~ FpAdd_6U_10U_mux_2_tmp_23) | (~ (chn_inp_in_crt_sva_11_739_736_1[0]))
      | (cfg_precision_1_sva_st_88[0]) | not_tmp_698);
  assign and_3276_nl = inp_lookup_1_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2
      & main_stage_v_12 & (chn_inp_in_crt_sva_12_739_736_1[0]) & (cfg_precision_1_sva_st_89==2'b10);
  assign mux_781_nl = MUX_s_1_2_2((and_3276_nl), (nor_1418_nl), or_11_cse);
  assign or_1676_nl = nor_1896_cse | FpAdd_6U_10U_mux_2_tmp_23 | FpNormalize_6U_23U_if_FpNormalize_6U_23U_if_nand_tmp
      | (~ (chn_inp_in_crt_sva_11_739_736_1[0])) | (cfg_precision_1_sva_st_88[0])
      | not_tmp_698;
  assign or_1679_nl = FpAdd_6U_10U_mux_2_tmp_23 | FpNormalize_6U_23U_if_FpNormalize_6U_23U_if_nand_tmp
      | (~ (chn_inp_in_crt_sva_11_739_736_1[0])) | (cfg_precision_1_sva_st_88[0])
      | not_tmp_698;
  assign mux_783_nl = MUX_s_1_2_2(or_tmp_1665, (or_1679_nl), or_11_cse);
  assign mux_784_nl = MUX_s_1_2_2((mux_783_nl), (or_1676_nl), reg_FpNormalize_6U_23U_lor_1_lpi_1_dfm_4_cse);
  assign nor_1415_nl = ~(FpAdd_6U_10U_mux_2_tmp_23 | (~ (chn_inp_in_crt_sva_11_739_736_1[0]))
      | (cfg_precision_1_sva_st_88[0]) | not_tmp_698);
  assign nor_1416_nl = ~(inp_lookup_1_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2
      | (~ main_stage_v_12) | (~ (chn_inp_in_crt_sva_12_739_736_1[0])) | (cfg_precision_1_sva_st_89!=2'b10));
  assign mux_785_nl = MUX_s_1_2_2((nor_1416_nl), (nor_1415_nl), or_11_cse);
  assign nand_87_nl = ~(main_stage_v_12 & (~((~((~ IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_24)
      | IsNaN_6U_10U_2_land_1_lpi_1_dfm_26)) | (~ (chn_inp_in_crt_sva_12_739_736_1[0]))
      | (cfg_precision_1_sva_st_89!=2'b10))));
  assign mux_787_nl = MUX_s_1_2_2(or_tmp_1690, (nand_87_nl), IsNaN_6U_10U_3_land_1_lpi_1_dfm_8);
  assign mux_788_nl = MUX_s_1_2_2((mux_787_nl), mux_tmp_708, or_11_cse);
  assign and_3275_nl = main_stage_v_12 & (chn_inp_in_crt_sva_12_739_736_1[0]);
  assign mux_791_nl = MUX_s_1_2_2((and_3275_nl), nor_tmp_227, or_11_cse);
  assign or_1708_nl = (~ FpAdd_6U_10U_mux_18_tmp_23) | (~ (chn_inp_in_crt_sva_11_739_736_1[1]))
      | (cfg_precision_1_sva_st_102[0]) | not_tmp_703;
  assign mux_798_nl = MUX_s_1_2_2(or_tmp_1697, (or_1708_nl), or_11_cse);
  assign or_1712_nl = FpAdd_6U_10U_mux_18_tmp_23 | FpNormalize_6U_23U_if_FpNormalize_6U_23U_if_nand_1_tmp
      | (~ (chn_inp_in_crt_sva_11_739_736_1[1])) | (cfg_precision_1_sva_st_102[0])
      | not_tmp_703;
  assign mux_800_nl = MUX_s_1_2_2(or_tmp_1699, (or_1712_nl), or_11_cse);
  assign nor_1410_nl = ~(FpAdd_6U_10U_mux_18_tmp_23 | (~ (chn_inp_in_crt_sva_11_739_736_1[1]))
      | (cfg_precision_1_sva_st_102[0]) | not_tmp_703);
  assign nor_1411_nl = ~(inp_lookup_2_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2
      | (~ main_stage_v_12) | (~ (chn_inp_in_crt_sva_12_739_736_1[1])) | (cfg_precision_1_sva_st_103!=2'b10));
  assign mux_801_nl = MUX_s_1_2_2((nor_1411_nl), (nor_1410_nl), or_11_cse);
  assign nor_1408_nl = ~((~ main_stage_v_12) | (~ (chn_inp_in_crt_sva_12_739_736_1[1]))
      | (cfg_precision_1_sva_st_103[0]) | (~((cfg_precision_1_sva_st_103[1]) & ((~((~
      IsNaN_6U_10U_3_land_2_lpi_1_dfm_8) | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_24))
      | IsNaN_6U_10U_2_land_2_lpi_1_dfm_26))));
  assign mux_802_nl = MUX_s_1_2_2((nor_1408_nl), nor_1407_cse, or_11_cse);
  assign and_3274_nl = main_stage_v_12 & (chn_inp_in_crt_sva_12_739_736_1[1]);
  assign mux_805_nl = MUX_s_1_2_2((and_3274_nl), nor_tmp_230, or_11_cse);
  assign nor_1404_nl = ~((~ FpAdd_6U_10U_mux_34_tmp_23) | (~ (chn_inp_in_crt_sva_11_739_736_1[2]))
      | (cfg_precision_1_sva_st_114[0]) | not_tmp_708);
  assign nor_1405_nl = ~((~ inp_lookup_3_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2)
      | (cfg_precision_1_sva_st_115[0]) | not_tmp_733);
  assign mux_815_nl = MUX_s_1_2_2((nor_1405_nl), (nor_1404_nl), or_11_cse);
  assign nor_1400_nl = ~(nor_1896_cse | FpAdd_6U_10U_mux_34_tmp_23 | FpNormalize_6U_23U_if_FpNormalize_6U_23U_if_nand_2_tmp
      | (~ (chn_inp_in_crt_sva_11_739_736_1[2])) | (cfg_precision_1_sva_st_114[0])
      | not_tmp_708);
  assign nor_1402_nl = ~(FpAdd_6U_10U_mux_34_tmp_23 | FpNormalize_6U_23U_if_FpNormalize_6U_23U_if_nand_2_tmp
      | (~ (chn_inp_in_crt_sva_11_739_736_1[2])) | (cfg_precision_1_sva_st_114[0])
      | not_tmp_708);
  assign nor_1403_nl = ~(inp_lookup_3_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2
      | (cfg_precision_1_sva_st_115[0]) | not_tmp_733);
  assign mux_817_nl = MUX_s_1_2_2((nor_1403_nl), (nor_1402_nl), or_11_cse);
  assign mux_818_nl = MUX_s_1_2_2((mux_817_nl), (nor_1400_nl), FpNormalize_6U_23U_lor_3_lpi_1_dfm_5);
  assign or_1763_nl = FpAdd_6U_10U_mux_34_tmp_23 | (~ (chn_inp_in_crt_sva_11_739_736_1[2]))
      | (cfg_precision_1_sva_st_114[0]) | not_tmp_708;
  assign mux_819_nl = MUX_s_1_2_2(or_tmp_1741, (or_1763_nl), or_11_cse);
  assign nor_1398_nl = ~((~ main_stage_v_12) | (~ (chn_inp_in_crt_sva_12_739_736_1[2]))
      | (cfg_precision_1_sva_st_115[0]) | (~((cfg_precision_1_sva_st_115[1]) & ((~((~
      IsNaN_6U_10U_3_land_3_lpi_1_dfm_8) | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_24))
      | IsNaN_6U_10U_2_land_3_lpi_1_dfm_26))));
  assign mux_820_nl = MUX_s_1_2_2((nor_1398_nl), nor_1397_cse, or_11_cse);
  assign and_3273_nl = (chn_inp_in_crt_sva_12_739_736_1[2]) & main_stage_v_12;
  assign mux_823_nl = MUX_s_1_2_2((and_3273_nl), nor_tmp_232, or_11_cse);
  assign nor_1394_nl = ~((~ FpAdd_6U_10U_mux_50_tmp_23) | (~ (chn_inp_in_crt_sva_11_739_736_1[3]))
      | (cfg_precision_1_sva_st_126[0]) | not_tmp_711);
  assign and_3384_nl = inp_lookup_4_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2
      & main_stage_v_12 & (chn_inp_in_crt_sva_12_739_736_1[3]) & (cfg_precision_1_sva_st_127==2'b10);
  assign mux_828_nl = MUX_s_1_2_2((and_3384_nl), (nor_1394_nl), or_11_cse);
  assign or_1797_nl = FpAdd_6U_10U_mux_50_tmp_23 | FpNormalize_6U_23U_if_FpNormalize_6U_23U_if_nand_3_tmp
      | (~ (chn_inp_in_crt_sva_11_739_736_1[3])) | (cfg_precision_1_sva_st_126[0])
      | not_tmp_711;
  assign mux_830_nl = MUX_s_1_2_2(or_tmp_1784, (or_1797_nl), or_11_cse);
  assign nor_1392_nl = ~(FpAdd_6U_10U_mux_50_tmp_23 | (~ (chn_inp_in_crt_sva_11_739_736_1[3]))
      | (cfg_precision_1_sva_st_126[0]) | not_tmp_711);
  assign nor_1393_nl = ~(inp_lookup_4_FpAdd_6U_10U_slc_FpAdd_6U_10U_int_mant_p1_23_itm_2
      | (~ main_stage_v_12) | (~ (chn_inp_in_crt_sva_12_739_736_1[3])) | (cfg_precision_1_sva_st_127!=2'b10));
  assign mux_831_nl = MUX_s_1_2_2((nor_1393_nl), (nor_1392_nl), or_11_cse);
  assign nand_665_nl = ~(((~((~ IsNaN_6U_10U_3_land_lpi_1_dfm_8) | IsNaN_6U_10U_2_land_lpi_1_dfm_st_23))
      | IsNaN_6U_10U_2_land_lpi_1_dfm_26) & main_stage_v_12 & (chn_inp_in_crt_sva_12_739_736_1[3])
      & (cfg_precision_1_sva_st_127==2'b10));
  assign mux_833_nl = MUX_s_1_2_2((nand_665_nl), mux_tmp_754, or_11_cse);
  assign and_3272_nl = main_stage_v_12 & (chn_inp_in_crt_sva_12_739_736_1[3]);
  assign mux_835_nl = MUX_s_1_2_2((and_3272_nl), nor_tmp_234, or_11_cse);
  assign or_1821_nl = (chn_inp_in_crt_sva_12_739_736_1[0]) | (~ main_stage_v_12);
  assign mux_837_nl = MUX_s_1_2_2((or_1821_nl), or_tmp_1818, or_11_cse);
  assign mux_838_nl = MUX_s_1_2_2(nor_tmp_250, nor_tmp_227, or_11_cse);
  assign nor_1387_nl = ~((~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ nor_tmp_250));
  assign mux_839_nl = MUX_s_1_2_2((nor_1387_nl), (mux_838_nl), inp_lookup_if_unequal_tmp_12);
  assign mux_843_nl = MUX_s_1_2_2(nor_tmp_252, nor_tmp_234, or_11_cse);
  assign nor_1386_nl = ~((~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ nor_tmp_252));
  assign mux_844_nl = MUX_s_1_2_2((nor_1386_nl), (mux_843_nl), inp_lookup_if_unequal_tmp_12);
  assign or_1832_nl = (chn_inp_in_crt_sva_12_739_736_1[3]) | (~ main_stage_v_12);
  assign mux_842_nl = MUX_s_1_2_2((or_1832_nl), or_tmp_1826, or_11_cse);
  assign or_1843_nl = (chn_inp_in_crt_sva_12_739_736_1[1]) | (~ main_stage_v_12);
  assign mux_847_nl = MUX_s_1_2_2((or_1843_nl), or_tmp_1840, or_11_cse);
  assign and_3266_nl = inp_lookup_if_unequal_tmp_19 & (chn_inp_in_crt_sva_12_739_736_1[1])
      & main_stage_v_12;
  assign mux_848_nl = MUX_s_1_2_2((and_3266_nl), nor_tmp_253, or_11_cse);
  assign mux_851_nl = MUX_s_1_2_2(nor_tmp_256, nor_tmp_232, or_11_cse);
  assign nor_1385_nl = ~((~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ nor_tmp_256));
  assign mux_852_nl = MUX_s_1_2_2((nor_1385_nl), (mux_851_nl), inp_lookup_if_unequal_tmp_12);
  assign or_1852_nl = (chn_inp_in_crt_sva_12_739_736_1[2]) | (~ main_stage_v_12);
  assign mux_850_nl = MUX_s_1_2_2((or_1852_nl), or_tmp_1849, or_11_cse);
  assign nor_732_nl = ~((cfg_precision_1_sva_st_80[1]) | (~ or_dcpl_159));
  assign or_4349_nl = (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[0]) |
      (cfg_precision_1_sva_st_80[0]);
  assign mux_1872_nl = MUX_s_1_2_2((nor_732_nl), or_dcpl_159, or_4349_nl);
  assign or_4671_nl = main_stage_v_3 | (~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[0])
      | (cfg_precision_1_sva_st_91!=2'b10);
  assign mux_1919_nl = MUX_s_1_2_2((or_4671_nl), (mux_1872_nl), or_11_cse);
  assign nor_1375_nl = ~((~((~ (inp_lookup_1_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21]))
      | inp_lookup_1_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1)) | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_14);
  assign nor_1377_nl = ~((FpMul_6U_10U_2_p_mant_p1_1_sva[21]) | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_14);
  assign mux_855_nl = MUX_s_1_2_2((nor_1377_nl), (nor_1375_nl), nor_44_cse);
  assign nand_89_nl = ~((~(FpMul_6U_10U_2_lor_6_lpi_1_dfm_5 | (~ inp_lookup_1_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2)))
      & (mux_855_nl));
  assign mux_856_nl = MUX_s_1_2_2((nand_89_nl), IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_14,
      IsNaN_6U_10U_7_land_1_lpi_1_dfm_5);
  assign mux_858_nl = MUX_s_1_2_2(nand_tmp_90, (mux_856_nl), or_11_cse);
  assign mux_861_nl = MUX_s_1_2_2(not_tmp_776, (mux_858_nl), nor_257_cse);
  assign nor_1378_nl = ~((cfg_precision_1_sva_st_90!=2'b10) | (chn_inp_in_crt_sva_1_739_395_1[341]));
  assign nor_1379_nl = ~((~ chn_inp_in_rsci_bawt) | (cfg_precision_rsci_d!=2'b10)
      | (chn_inp_in_rsci_d_mxwt[736]));
  assign mux_862_nl = MUX_s_1_2_2((nor_1379_nl), (nor_1378_nl), main_stage_v_1);
  assign mux_863_nl = MUX_s_1_2_2(not_tmp_776, nand_tmp_90, nor_1380_cse);
  assign mux_864_nl = MUX_s_1_2_2((mux_863_nl), (mux_862_nl), or_11_cse);
  assign mux_865_nl = MUX_s_1_2_2((mux_864_nl), (mux_861_nl), main_stage_v_2);
  assign nor_1349_nl = ~((~((~ (inp_lookup_3_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21]))
      | inp_lookup_3_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1)) | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_14);
  assign nor_1351_nl = ~((FpMul_6U_10U_2_p_mant_p1_3_sva[21]) | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_14);
  assign mux_889_nl = MUX_s_1_2_2((nor_1351_nl), (nor_1349_nl), nor_67_cse);
  assign nand_97_nl = ~((~(FpMul_6U_10U_2_lor_8_lpi_1_dfm_5 | (~ inp_lookup_3_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2)))
      & (mux_889_nl));
  assign mux_890_nl = MUX_s_1_2_2((nand_97_nl), IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_14,
      IsNaN_6U_10U_7_land_3_lpi_1_dfm_5);
  assign mux_892_nl = MUX_s_1_2_2(nand_tmp_98, (mux_890_nl), or_11_cse);
  assign mux_895_nl = MUX_s_1_2_2(not_tmp_810, (mux_892_nl), nor_275_cse);
  assign nor_1352_nl = ~((cfg_precision_1_sva_st_90!=2'b10) | (chn_inp_in_crt_sva_1_739_395_1[343]));
  assign nor_1353_nl = ~((~ chn_inp_in_rsci_bawt) | (cfg_precision_rsci_d!=2'b10)
      | (chn_inp_in_rsci_d_mxwt[738]));
  assign mux_896_nl = MUX_s_1_2_2((nor_1353_nl), (nor_1352_nl), main_stage_v_1);
  assign mux_897_nl = MUX_s_1_2_2(not_tmp_810, nand_tmp_98, nor_1354_cse);
  assign mux_898_nl = MUX_s_1_2_2((mux_897_nl), (mux_896_nl), or_11_cse);
  assign mux_899_nl = MUX_s_1_2_2((mux_898_nl), (mux_895_nl), main_stage_v_2);
  assign mux_922_nl = MUX_s_1_2_2(nand_tmp_5, nand_728_cse_1, or_11_cse);
  assign mux_924_nl = MUX_s_1_2_2(nand_tmp_12, or_tmp_621, or_11_cse);
  assign mux_2105_nl = MUX_s_1_2_2(or_tmp_4714, nor_1336_cse_1, or_2010_cse);
  assign mux_2106_nl = MUX_s_1_2_2((mux_2105_nl), or_tmp_4714, chn_inp_in_crt_sva_1_739_395_1[344]);
  assign and_4209_nl = or_tmp_4721 & (~ or_2010_cse);
  assign mux_2109_nl = MUX_s_1_2_2((and_4209_nl), or_tmp_4721, chn_inp_in_crt_sva_1_739_395_1[343]);
  assign mux_2112_nl = MUX_s_1_2_2(or_tmp_4726, and_4210_cse, or_2010_cse);
  assign mux_2113_nl = MUX_s_1_2_2((mux_2112_nl), or_tmp_4726, chn_inp_in_crt_sva_1_739_395_1[341]);
  assign mux_2115_nl = MUX_s_1_2_2(or_tmp_4730, nor_1336_cse_1, or_2010_cse);
  assign mux_2116_nl = MUX_s_1_2_2((mux_2115_nl), or_tmp_4730, chn_inp_in_crt_sva_1_739_395_1[342]);
  assign and_227_nl = main_stage_v_1 & (chn_inp_in_crt_sva_1_739_395_1[341]) & or_2010_cse;
  assign mux_939_nl = MUX_s_1_2_2(and_tmp_29, (and_227_nl), or_11_cse);
  assign or_171_nl = (~ main_stage_v_1) | (chn_inp_in_crt_sva_1_739_395_1[341]) |
      (~ inp_lookup_1_FpMul_6U_10U_2_else_2_if_acc_itm_6) | or_5873_cse | (cfg_precision_1_sva_st_90!=2'b10);
  assign mux_117_nl = MUX_s_1_2_2(or_5800_cse, (or_171_nl), or_11_cse);
  assign or_174_nl = nor_1896_cse | (~ main_stage_v_1) | (chn_inp_in_crt_sva_1_739_395_1[341])
      | (~ inp_lookup_1_FpMul_6U_10U_2_else_2_if_acc_itm_6) | or_5873_cse | (cfg_precision_1_sva_st_90!=2'b10);
  assign mux_118_nl = MUX_s_1_2_2((or_174_nl), (mux_117_nl), nor_44_cse);
  assign nor_1695_nl = ~(((FpFractionToFloat_35U_6U_10U_1_mux_tmp[4:3]==2'b11) &
      (IntLeadZero_35U_1_leading_sign_35_0_rtn_1_sva_2[5]) & inp_lookup_1_FpMantRNE_36U_11U_1_else_and_svs_2
      & (~ IsNaN_6U_10U_6_nor_tmp) & FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_st_2
      & (FpFractionToFloat_35U_6U_10U_1_mux_tmp[2:0]==3'b111) & (~ (chn_inp_in_crt_sva_1_739_395_1[341])))
      | (~ main_stage_v_1) | (cfg_precision_1_sva_st_90!=2'b10));
  assign and_3392_nl = (chn_inp_in_crt_sva_1_739_395_1[341]) & main_stage_v_1 & (cfg_precision_1_sva_st_90==2'b10);
  assign mux_120_nl = MUX_s_1_2_2((and_3392_nl), (nor_1695_nl), and_3149_cse);
  assign mux_121_nl = MUX_s_1_2_2((mux_120_nl), nor_1318_cse, nor_5_cse);
  assign nor_1698_nl = ~(FpMul_6U_10U_2_lor_6_lpi_1_dfm_st_3 | (~ inp_lookup_1_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs)
      | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10));
  assign or_192_nl = (~((~ IsNaN_6U_10U_7_land_1_lpi_1_dfm_5) | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_14))
      | (chn_inp_in_crt_sva_2_739_736_1[0]);
  assign mux_122_nl = MUX_s_1_2_2((nor_1698_nl), nor_1697_cse, or_192_nl);
  assign mux_123_nl = MUX_s_1_2_2((mux_122_nl), (mux_121_nl), or_11_cse);
  assign and_231_nl = main_stage_v_1 & (chn_inp_in_crt_sva_1_739_395_1[342]) & or_2010_cse;
  assign mux_941_nl = MUX_s_1_2_2(and_tmp_35, (and_231_nl), or_11_cse);
  assign or_239_nl = (~ main_stage_v_1) | (chn_inp_in_crt_sva_1_739_395_1[342]) |
      (~ inp_lookup_2_FpMul_6U_10U_2_else_2_if_acc_itm_6) | or_5890_cse | (cfg_precision_1_sva_st_90!=2'b10);
  assign mux_140_nl = MUX_s_1_2_2(or_tmp_238, (or_239_nl), or_11_cse);
  assign nor_1677_nl = ~(((FpFractionToFloat_35U_6U_10U_1_mux_40_tmp==5'b11111) &
      (IntLeadZero_35U_1_leading_sign_35_0_rtn_2_sva_2[5]) & inp_lookup_2_FpMantRNE_36U_11U_1_else_and_svs_2
      & (~ IsNaN_6U_10U_6_nor_1_tmp) & FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_st_2
      & (~ (chn_inp_in_crt_sva_1_739_395_1[342]))) | (~ main_stage_v_1) | (cfg_precision_1_sva_st_90!=2'b10));
  assign and_3390_nl = (chn_inp_in_crt_sva_1_739_395_1[342]) & main_stage_v_1 & (cfg_precision_1_sva_st_90==2'b10);
  assign mux_143_nl = MUX_s_1_2_2((and_3390_nl), (nor_1677_nl), and_4145_cse);
  assign mux_144_nl = MUX_s_1_2_2((mux_143_nl), nor_1318_cse, nor_13_cse);
  assign nor_1680_nl = ~(FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_3 | (~ inp_lookup_2_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs)
      | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10));
  assign or_258_nl = (~((~ IsNaN_6U_10U_7_land_2_lpi_1_dfm_5) | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_14))
      | (chn_inp_in_crt_sva_2_739_736_1[1]);
  assign mux_145_nl = MUX_s_1_2_2((nor_1680_nl), nor_1697_cse, or_258_nl);
  assign mux_146_nl = MUX_s_1_2_2((mux_145_nl), (mux_144_nl), or_11_cse);
  assign and_235_nl = (chn_inp_in_crt_sva_1_739_395_1[343]) & main_stage_v_1 & or_2010_cse;
  assign mux_943_nl = MUX_s_1_2_2(and_tmp_42, (and_235_nl), or_11_cse);
  assign or_311_nl = (chn_inp_in_crt_sva_1_739_395_1[343]) | (~ main_stage_v_1) |
      (~ inp_lookup_3_FpMul_6U_10U_2_else_2_if_acc_itm_6_1) | FpMul_6U_10U_2_if_2_FpMul_6U_10U_2_if_2_or_5_tmp
      | (cfg_precision_1_sva_st_90!=2'b10);
  assign mux_162_nl = MUX_s_1_2_2(or_tmp_306, (or_311_nl), or_11_cse);
  assign or_314_nl = nor_1896_cse | (chn_inp_in_crt_sva_1_739_395_1[343]) | (~ main_stage_v_1)
      | (~ inp_lookup_3_FpMul_6U_10U_2_else_2_if_acc_itm_6_1) | FpMul_6U_10U_2_if_2_FpMul_6U_10U_2_if_2_or_5_tmp
      | (cfg_precision_1_sva_st_90!=2'b10);
  assign mux_163_nl = MUX_s_1_2_2((or_314_nl), (mux_162_nl), nor_67_cse);
  assign nand_458_nl = ~((FpFractionToFloat_35U_6U_10U_1_mux_41_tmp==5'b11111) &
      (IntLeadZero_35U_1_leading_sign_35_0_rtn_3_sva_2[5]) & inp_lookup_3_FpMantRNE_36U_11U_1_else_and_svs_2
      & (~ IsNaN_6U_10U_6_nor_2_tmp) & FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_st_2
      & (~ (chn_inp_in_crt_sva_1_739_395_1[343])));
  assign mux_944_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_1_739_395_1[343]), (nand_458_nl),
      and_3249_cse);
  assign nor_1305_nl = ~((~ main_stage_v_1) | (cfg_precision_1_sva_st_90[0]) | (~((cfg_precision_1_sva_st_90[1])
      & (nor_301_cse | (mux_944_nl)))));
  assign nor_1307_nl = ~(FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_3 | (~ inp_lookup_3_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs)
      | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10));
  assign or_2090_nl = (~((~ IsNaN_6U_10U_7_land_3_lpi_1_dfm_5) | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_14))
      | (chn_inp_in_crt_sva_2_739_736_1[2]);
  assign mux_945_nl = MUX_s_1_2_2((nor_1307_nl), nor_1697_cse, or_2090_nl);
  assign mux_946_nl = MUX_s_1_2_2((mux_945_nl), (nor_1305_nl), or_11_cse);
  assign and_237_nl = (chn_inp_in_crt_sva_1_739_395_1[344]) & main_stage_v_1 & or_2010_cse;
  assign mux_947_nl = MUX_s_1_2_2(and_tmp_50, (and_237_nl), or_11_cse);
  assign or_374_nl = (chn_inp_in_crt_sva_1_739_395_1[344]) | (~ main_stage_v_1) |
      (~ inp_lookup_4_FpMul_6U_10U_2_else_2_if_acc_itm_6) | FpMul_6U_10U_2_if_2_FpMul_6U_10U_2_if_2_or_7_tmp
      | (cfg_precision_1_sva_st_90!=2'b10);
  assign mux_180_nl = MUX_s_1_2_2(or_tmp_374, (or_374_nl), or_11_cse);
  assign nor_1300_nl = ~((z_out[49]) | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10));
  assign nor_1301_nl = ~(and_3246_cse | and_3358_cse | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10));
  assign mux_949_nl = MUX_s_1_2_2((nor_1301_nl), (nor_1300_nl), chn_inp_in_crt_sva_2_739_736_1[0]);
  assign nor_1302_nl = ~((FpAdd_8U_23U_int_mant_p1_1_lpi_1_dfm_3_49_1_1[48]) | inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4
      | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10));
  assign nor_1303_nl = ~(IsNaN_6U_10U_5_land_1_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_15
      | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10));
  assign mux_950_nl = MUX_s_1_2_2((nor_1303_nl), (nor_1302_nl), chn_inp_in_crt_sva_3_739_736_1[0]);
  assign mux_951_nl = MUX_s_1_2_2((mux_950_nl), (mux_949_nl), or_11_cse);
  assign nor_1296_nl = ~((z_out_1[49]) | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10));
  assign nor_1297_nl = ~(and_3244_cse | and_3355_cse | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10));
  assign mux_952_nl = MUX_s_1_2_2((nor_1297_nl), (nor_1296_nl), chn_inp_in_crt_sva_2_739_736_1[1]);
  assign nor_1298_nl = ~((FpAdd_8U_23U_int_mant_p1_2_lpi_1_dfm_3_49_1_1[48]) | inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4
      | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10));
  assign nor_1299_nl = ~(IsNaN_6U_10U_5_land_2_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_15
      | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10));
  assign mux_953_nl = MUX_s_1_2_2((nor_1299_nl), (nor_1298_nl), chn_inp_in_crt_sva_3_739_736_1[1]);
  assign mux_954_nl = MUX_s_1_2_2((mux_953_nl), (mux_952_nl), or_11_cse);
  assign nor_1292_nl = ~((z_out_2[49]) | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10));
  assign nor_1293_nl = ~(and_3242_cse | and_3351_cse | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10));
  assign mux_955_nl = MUX_s_1_2_2((nor_1293_nl), (nor_1292_nl), chn_inp_in_crt_sva_2_739_736_1[2]);
  assign nor_1294_nl = ~((FpAdd_8U_23U_int_mant_p1_3_lpi_1_dfm_3_49_1_1[48]) | inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4
      | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10));
  assign nor_1295_nl = ~(IsNaN_6U_10U_5_land_3_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_15
      | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10));
  assign mux_956_nl = MUX_s_1_2_2((nor_1295_nl), (nor_1294_nl), chn_inp_in_crt_sva_3_739_736_1[2]);
  assign mux_957_nl = MUX_s_1_2_2((mux_956_nl), (mux_955_nl), or_11_cse);
  assign nor_1288_nl = ~((z_out_3[49]) | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10));
  assign nor_1289_nl = ~(and_3240_cse | and_3345_cse | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10));
  assign mux_958_nl = MUX_s_1_2_2((nor_1289_nl), (nor_1288_nl), chn_inp_in_crt_sva_2_739_736_1[3]);
  assign nor_1290_nl = ~((FpAdd_8U_23U_int_mant_p1_lpi_1_dfm_3_49_1_1[48]) | inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4
      | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10));
  assign nor_1291_nl = ~(IsNaN_6U_10U_5_land_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_lpi_1_dfm_st_15
      | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10));
  assign mux_959_nl = MUX_s_1_2_2((nor_1291_nl), (nor_1290_nl), chn_inp_in_crt_sva_3_739_736_1[3]);
  assign mux_960_nl = MUX_s_1_2_2((mux_959_nl), (mux_958_nl), or_11_cse);
  assign nor_1284_nl = ~(((~ IsNaN_6U_10U_4_nor_tmp) & inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_5_1
      & (inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_4_0_1==5'b11111) & IsNaN_8U_23U_land_1_lpi_1_dfm_st_4
      & (~ (chn_inp_in_crt_sva_2_739_736_1[0]))) | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10));
  assign mux_961_nl = MUX_s_1_2_2((nor_1284_nl), and_3393_cse, and_3246_cse);
  assign nor_1285_nl = ~((~((~(IsNaN_6U_10U_5_land_1_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_15))
      | (chn_inp_in_crt_sva_3_739_736_1[0]))) | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10));
  assign mux_962_nl = MUX_s_1_2_2((nor_1285_nl), (mux_961_nl), or_11_cse);
  assign nor_1279_nl = ~(((~ IsNaN_6U_10U_4_nor_1_tmp) & inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_6_5_1
      & (inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_6_4_0_1==5'b11111) & IsNaN_8U_23U_land_2_lpi_1_dfm_st_4
      & (~ (chn_inp_in_crt_sva_2_739_736_1[1]))) | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10));
  assign mux_963_nl = MUX_s_1_2_2((nor_1279_nl), and_3391_cse, and_3244_cse);
  assign nor_1280_nl = ~((~((~(IsNaN_6U_10U_5_land_2_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_15))
      | (chn_inp_in_crt_sva_3_739_736_1[1]))) | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10));
  assign mux_964_nl = MUX_s_1_2_2((nor_1280_nl), (mux_963_nl), or_11_cse);
  assign nor_1275_nl = ~(((~ IsNaN_6U_10U_4_nor_2_tmp) & inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_6_5_1
      & (inp_lookup_else_if_a0_15_10_3_lpi_1_dfm_6_4_0_1==5'b11111) & IsNaN_8U_23U_land_3_lpi_1_dfm_st_4
      & (~ (chn_inp_in_crt_sva_2_739_736_1[2]))) | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10));
  assign mux_965_nl = MUX_s_1_2_2((nor_1275_nl), and_3401_cse, and_3242_cse);
  assign nor_1276_nl = ~((~((~(IsNaN_6U_10U_5_land_3_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_15))
      | (chn_inp_in_crt_sva_3_739_736_1[2]))) | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10));
  assign mux_966_nl = MUX_s_1_2_2((nor_1276_nl), (mux_965_nl), or_11_cse);
  assign or_460_nl = (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[0]) | (cfg_precision_1_sva_st_80!=2'b10)
      | FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_3;
  assign mux_214_nl = MUX_s_1_2_2((or_460_nl), or_5800_cse, or_11_cse);
  assign or_458_nl = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[0]) | (cfg_precision_1_sva_st_80!=2'b10)
      | FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_3;
  assign mux_210_nl = MUX_s_1_2_2((or_458_nl), (mux_214_nl), nor_35_cse);
  assign FpMul_6U_10U_2_else_2_else_and_nl = inp_lookup_1_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1
      & (inp_lookup_1_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21]);
  assign or_2179_nl = (~((~ (inp_lookup_1_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21]))
      | inp_lookup_1_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1 | (chn_inp_in_crt_sva_2_739_736_1[0])))
      | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10);
  assign mux_967_nl = MUX_s_1_2_2(nand_772_cse, (or_2179_nl), inp_lookup_1_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2);
  assign or_2174_nl = inp_lookup_1_FpMantRNE_22U_11U_2_else_and_tmp | FpMul_6U_10U_2_lor_6_lpi_1_dfm_5;
  assign mux_968_nl = MUX_s_1_2_2((mux_967_nl), or_2176_cse, or_2174_nl);
  assign or_2171_nl = FpMul_6U_10U_2_lor_6_lpi_1_dfm_st_3 | (~ inp_lookup_1_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs)
      | IsNaN_6U_10U_7_land_1_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_14;
  assign mux_969_nl = MUX_s_1_2_2((mux_968_nl), nand_772_cse, or_2171_nl);
  assign or_2185_nl = (~((~((~(nor_1273_cse | inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4))
      | FpMul_6U_10U_2_lor_6_lpi_1_dfm_st_4 | (~ inp_lookup_1_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4)
      | IsNaN_6U_10U_6_land_1_lpi_1_dfm_5 | IsNaN_6U_10U_7_land_1_lpi_1_dfm_6)) |
      (chn_inp_in_crt_sva_3_739_736_1[0]))) | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_970_nl = MUX_s_1_2_2((or_2185_nl), (mux_969_nl), or_11_cse);
  assign nor_1267_nl = ~((~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[0])
      | (~ IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_14) | (cfg_precision_1_sva_st_91!=2'b10));
  assign nor_1268_nl = ~((~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[0])
      | (cfg_precision_1_sva_st_80[0]) | (~((cfg_precision_1_sva_st_80[1]) & IsNaN_6U_10U_6_land_1_lpi_1_dfm_5)));
  assign mux_971_nl = MUX_s_1_2_2((nor_1268_nl), (nor_1267_nl), or_11_cse);
  assign nor_1265_nl = ~((~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[0])
      | (~ IsNaN_6U_10U_7_land_1_lpi_1_dfm_5) | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_14
      | (cfg_precision_1_sva_st_91!=2'b10));
  assign nor_1266_nl = ~((~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[0])
      | (cfg_precision_1_sva_st_80!=2'b10) | (~ IsNaN_6U_10U_7_land_1_lpi_1_dfm_6)
      | IsNaN_6U_10U_6_land_1_lpi_1_dfm_5);
  assign mux_972_nl = MUX_s_1_2_2((nor_1266_nl), (nor_1265_nl), or_11_cse);
  assign FpMul_6U_10U_2_FpMul_6U_10U_2_and_nl = (inp_lookup_1_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1
      | (~ FpMul_6U_10U_2_p_mant_p1_1_sva_mx2_21)) & inp_lookup_1_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2;
  assign or_520_nl = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[1]) | FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_3
      | (cfg_precision_1_sva_st_80!=2'b10);
  assign or_522_nl = (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[1]) | FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_3
      | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_252_nl = MUX_s_1_2_2((or_522_nl), or_tmp_234, or_11_cse);
  assign mux_248_nl = MUX_s_1_2_2((mux_252_nl), (or_520_nl), or_507_cse);
  assign nor_1261_nl = ~((~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[1])
      | (cfg_precision_1_sva_st_91!=2'b10) | FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_3
      | (~ inp_lookup_2_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs)
      | IsNaN_6U_10U_7_land_2_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_14
      | (~(or_tmp_2199 | (inp_lookup_2_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2
      & ((~ (inp_lookup_2_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21])) | inp_lookup_2_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1)))));
  assign nor_1263_nl = ~((~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[1])
      | (cfg_precision_1_sva_st_80!=2'b10) | FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_4
      | (~ inp_lookup_2_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4)
      | IsNaN_6U_10U_6_land_2_lpi_1_dfm_5 | IsNaN_6U_10U_7_land_2_lpi_1_dfm_6 | (~((nor_1264_cse
      | inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4)
      & (~(FpMul_6U_10U_2_else_2_else_and_1_itm_2 & (~(inp_lookup_2_FpMul_6U_10U_2_else_2_else_slc_FpMul_6U_10U_2_p_mant_p1_21_itm_2
      & FpMul_6U_10U_2_else_2_else_if_if_slc_FpMul_6U_10U_2_else_2_else_if_if_acc_1_5_mdf_2_sva_st_1)))))));
  assign mux_976_nl = MUX_s_1_2_2((nor_1263_nl), (nor_1261_nl), or_11_cse);
  assign FpMul_6U_10U_2_else_2_else_and_1_nl = inp_lookup_2_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1
      & (inp_lookup_2_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21]);
  assign or_2216_nl = (~((~ (inp_lookup_2_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21]))
      | inp_lookup_2_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1 | (chn_inp_in_crt_sva_2_739_736_1[1])))
      | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10);
  assign mux_977_nl = MUX_s_1_2_2(nand_358_cse, (or_2216_nl), inp_lookup_2_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2);
  assign mux_978_nl = MUX_s_1_2_2((mux_977_nl), or_2176_cse, or_tmp_2199);
  assign or_2211_nl = FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_3 | (~ inp_lookup_2_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs)
      | IsNaN_6U_10U_7_land_2_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_14;
  assign mux_979_nl = MUX_s_1_2_2((mux_978_nl), nand_358_cse, or_2211_nl);
  assign or_2223_nl = (~((~((~(nor_1264_cse | inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4))
      | FpMul_6U_10U_2_lor_7_lpi_1_dfm_st_4 | (~ inp_lookup_2_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4)
      | IsNaN_6U_10U_6_land_2_lpi_1_dfm_5 | IsNaN_6U_10U_7_land_2_lpi_1_dfm_6)) |
      (chn_inp_in_crt_sva_3_739_736_1[1]))) | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_980_nl = MUX_s_1_2_2((or_2223_nl), (mux_979_nl), or_11_cse);
  assign nor_1254_nl = ~((~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[1])
      | (cfg_precision_1_sva_st_91!=2'b10) | (~ IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_14));
  assign nor_1255_nl = ~((~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[1])
      | (~ IsNaN_6U_10U_6_land_2_lpi_1_dfm_5) | (cfg_precision_1_sva_st_80!=2'b10));
  assign mux_981_nl = MUX_s_1_2_2((nor_1255_nl), (nor_1254_nl), or_11_cse);
  assign nor_1252_nl = ~((~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[1])
      | (cfg_precision_1_sva_st_91!=2'b10) | (~ IsNaN_6U_10U_7_land_2_lpi_1_dfm_5)
      | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_14);
  assign nor_1253_nl = ~((~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[1])
      | IsNaN_6U_10U_6_land_2_lpi_1_dfm_5 | (~ IsNaN_6U_10U_7_land_2_lpi_1_dfm_6)
      | (cfg_precision_1_sva_st_80!=2'b10));
  assign mux_982_nl = MUX_s_1_2_2((nor_1253_nl), (nor_1252_nl), or_11_cse);
  assign FpMul_6U_10U_2_FpMul_6U_10U_2_and_16_nl = (inp_lookup_2_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1
      | (~ FpMul_6U_10U_2_p_mant_p1_2_sva_mx2_21)) & inp_lookup_2_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2;
  assign or_596_nl = (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[2]) | FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_3
      | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_297_nl = MUX_s_1_2_2((or_596_nl), or_tmp_306, or_11_cse);
  assign or_594_nl = (~ reg_chn_inp_out_rsci_ld_core_psct_cse) | chn_inp_out_rsci_bawt
      | (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[2]) | FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_3
      | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_286_nl = MUX_s_1_2_2((or_594_nl), (mux_297_nl), nor_55_cse);
  assign nor_1248_nl = ~((~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[2])
      | (cfg_precision_1_sva_st_91!=2'b10) | FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_3
      | (~ inp_lookup_3_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs)
      | IsNaN_6U_10U_7_land_3_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_14
      | (~(or_tmp_2234 | (inp_lookup_3_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2
      & ((~ (inp_lookup_3_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21])) | inp_lookup_3_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1)))));
  assign nor_1250_nl = ~((~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[2])
      | (cfg_precision_1_sva_st_80!=2'b10) | FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_4
      | (~ inp_lookup_3_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4)
      | IsNaN_6U_10U_6_land_3_lpi_1_dfm_5 | IsNaN_6U_10U_7_land_3_lpi_1_dfm_6 | (~((nor_1251_cse
      | inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4)
      & (~(FpMul_6U_10U_2_else_2_else_and_2_itm_2 & (~(inp_lookup_3_FpMul_6U_10U_2_else_2_else_slc_FpMul_6U_10U_2_p_mant_p1_21_itm_2
      & FpMul_6U_10U_2_else_2_else_if_if_slc_FpMul_6U_10U_2_else_2_else_if_if_acc_1_5_mdf_3_sva_st_1)))))));
  assign mux_986_nl = MUX_s_1_2_2((nor_1250_nl), (nor_1248_nl), or_11_cse);
  assign FpMul_6U_10U_2_else_2_else_and_2_nl = inp_lookup_3_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1
      & (inp_lookup_3_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21]);
  assign or_2254_nl = (~((~ (inp_lookup_3_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21]))
      | inp_lookup_3_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1 | (chn_inp_in_crt_sva_2_739_736_1[2])))
      | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10);
  assign mux_987_nl = MUX_s_1_2_2(or_tmp_277, (or_2254_nl), inp_lookup_3_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2);
  assign mux_988_nl = MUX_s_1_2_2((mux_987_nl), or_2176_cse, or_tmp_2234);
  assign or_2246_nl = FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_3 | (~ inp_lookup_3_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs)
      | IsNaN_6U_10U_7_land_3_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_14;
  assign mux_989_nl = MUX_s_1_2_2((mux_988_nl), or_tmp_277, or_2246_nl);
  assign or_2260_nl = (~((~((~(nor_1251_cse | inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4))
      | FpMul_6U_10U_2_lor_8_lpi_1_dfm_st_4 | (~ inp_lookup_3_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4)
      | IsNaN_6U_10U_6_land_3_lpi_1_dfm_5 | IsNaN_6U_10U_7_land_3_lpi_1_dfm_6)) |
      (chn_inp_in_crt_sva_3_739_736_1[2]))) | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_990_nl = MUX_s_1_2_2((or_2260_nl), (mux_989_nl), or_11_cse);
  assign nor_1241_nl = ~((chn_inp_in_crt_sva_2_739_736_1[2]) | (~ main_stage_v_2)
      | (cfg_precision_1_sva_st_91[0]) | (~((cfg_precision_1_sva_st_91[1]) & IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_14)));
  assign nor_1242_nl = ~((~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[2])
      | (~ IsNaN_6U_10U_6_land_3_lpi_1_dfm_5) | (cfg_precision_1_sva_st_80!=2'b10));
  assign mux_991_nl = MUX_s_1_2_2((nor_1242_nl), (nor_1241_nl), or_11_cse);
  assign nor_1239_nl = ~((chn_inp_in_crt_sva_2_739_736_1[2]) | (~ main_stage_v_2)
      | (cfg_precision_1_sva_st_91!=2'b10) | (~ IsNaN_6U_10U_7_land_3_lpi_1_dfm_5)
      | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_14);
  assign nor_1240_nl = ~((~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[2])
      | (~ IsNaN_6U_10U_7_land_3_lpi_1_dfm_6) | IsNaN_6U_10U_6_land_3_lpi_1_dfm_5
      | (cfg_precision_1_sva_st_80!=2'b10));
  assign mux_992_nl = MUX_s_1_2_2((nor_1240_nl), (nor_1239_nl), or_11_cse);
  assign FpMul_6U_10U_2_FpMul_6U_10U_2_and_17_nl = (inp_lookup_3_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1
      | (~ FpMul_6U_10U_2_p_mant_p1_3_sva_mx2_21)) & inp_lookup_3_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2;
  assign or_640_nl = (~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[3]) | (cfg_precision_1_sva_st_91!=2'b10)
      | inp_lookup_4_FpMul_6U_10U_1_oelse_1_acc_itm_7_1 | FpMul_6U_10U_1_if_2_FpMul_6U_10U_1_if_2_or_6_tmp
      | (~ inp_lookup_4_FpMul_6U_10U_1_else_2_if_acc_itm_6_1);
  assign or_642_nl = (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[3]) | (cfg_precision_1_sva_st_80!=2'b10)
      | FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_3;
  assign mux_336_nl = MUX_s_1_2_2((or_642_nl), (or_640_nl), or_11_cse);
  assign FpMul_6U_10U_2_else_2_else_and_3_nl = inp_lookup_4_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1
      & (inp_lookup_4_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21]);
  assign or_2277_nl = (~((~ (inp_lookup_4_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21]))
      | inp_lookup_4_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1 | (chn_inp_in_crt_sva_2_739_736_1[3])))
      | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10);
  assign mux_996_nl = MUX_s_1_2_2(nand_701_cse, (or_2277_nl), inp_lookup_4_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2);
  assign or_2274_nl = inp_lookup_4_FpMantRNE_22U_11U_2_else_and_tmp | FpMul_6U_10U_2_lor_1_lpi_1_dfm_5;
  assign mux_997_nl = MUX_s_1_2_2((mux_996_nl), or_2176_cse, or_2274_nl);
  assign or_2272_nl = FpMul_6U_10U_2_lor_1_lpi_1_dfm_st_3 | (~ inp_lookup_4_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs)
      | IsNaN_6U_10U_7_land_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_lpi_1_dfm_st_14;
  assign mux_998_nl = MUX_s_1_2_2((mux_997_nl), nand_701_cse, or_2272_nl);
  assign or_2287_nl = (~(nor_1237_cse | (chn_inp_in_crt_sva_3_739_736_1[3]))) | (~
      main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_999_nl = MUX_s_1_2_2((or_2287_nl), or_2282_cse, inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4);
  assign or_2278_nl = FpMul_6U_10U_2_lor_1_lpi_1_dfm_st_4 | (~ inp_lookup_4_FpMul_6U_10U_2_else_2_if_slc_FpMul_6U_10U_2_else_2_if_acc_6_svs_st_4)
      | IsNaN_6U_10U_6_land_lpi_1_dfm_5 | IsNaN_6U_10U_7_land_lpi_1_dfm_6;
  assign mux_1000_nl = MUX_s_1_2_2((mux_999_nl), nand_661_cse, or_2278_nl);
  assign mux_1001_nl = MUX_s_1_2_2((mux_1000_nl), (mux_998_nl), or_11_cse);
  assign nor_1233_nl = ~((~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[3])
      | (cfg_precision_1_sva_st_91[0]) | (~((cfg_precision_1_sva_st_91[1]) & IsNaN_6U_10U_2_land_lpi_1_dfm_st_14)));
  assign nor_1234_nl = ~((~ main_stage_v_3) | (~ IsNaN_6U_10U_6_land_lpi_1_dfm_5)
      | (chn_inp_in_crt_sva_3_739_736_1[3]) | (cfg_precision_1_sva_st_80!=2'b10));
  assign mux_1002_nl = MUX_s_1_2_2((nor_1234_nl), (nor_1233_nl), or_11_cse);
  assign nor_1231_nl = ~((~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[3])
      | (cfg_precision_1_sva_st_91!=2'b10) | (~ IsNaN_6U_10U_7_land_lpi_1_dfm_5)
      | IsNaN_6U_10U_2_land_lpi_1_dfm_st_14);
  assign nor_1232_nl = ~((~ main_stage_v_3) | (~ IsNaN_6U_10U_7_land_lpi_1_dfm_6)
      | IsNaN_6U_10U_6_land_lpi_1_dfm_5 | (chn_inp_in_crt_sva_3_739_736_1[3]) | (cfg_precision_1_sva_st_80!=2'b10));
  assign mux_1003_nl = MUX_s_1_2_2((nor_1232_nl), (nor_1231_nl), or_11_cse);
  assign FpMul_6U_10U_2_FpMul_6U_10U_2_and_18_nl = (inp_lookup_4_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1
      | (~ FpMul_6U_10U_2_p_mant_p1_sva_mx2_21)) & inp_lookup_4_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2;
  assign nor_1226_nl = ~(and_3240_cse | and_3345_cse | (~ main_stage_v_2) | (chn_inp_in_crt_sva_2_739_736_1[3])
      | (cfg_precision_1_sva_st_91!=2'b10));
  assign nor_1227_nl = ~((~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[3])
      | (cfg_precision_1_sva_st_80!=2'b10) | IsNaN_6U_10U_5_land_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_lpi_1_dfm_st_15);
  assign mux_1006_nl = MUX_s_1_2_2((nor_1227_nl), (nor_1226_nl), or_11_cse);
  assign FpMul_6U_10U_1_else_2_else_and_nl = inp_lookup_1_FpMul_6U_10U_1_else_2_else_if_if_acc_1_itm_5_1
      & (inp_lookup_1_FpMul_6U_10U_1_p_mant_p1_mul_tmp[21]);
  assign and_3222_nl = (chn_inp_in_crt_sva_3_739_736_1[0]) & main_stage_v_3 & (cfg_precision_1_sva_st_80==2'b10);
  assign nor_1218_nl = ~((~((((~ (inp_lookup_1_FpMul_6U_10U_1_p_mant_p1_mul_tmp[21]))
      | inp_lookup_1_FpMul_6U_10U_1_else_2_else_if_if_acc_1_itm_5_1) & inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4)
      | (chn_inp_in_crt_sva_3_739_736_1[0]))) | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10));
  assign or_2308_nl = FpMul_6U_10U_1_lor_6_lpi_1_dfm_5 | inp_lookup_1_FpMantRNE_22U_11U_1_else_and_tmp;
  assign mux_1007_nl = MUX_s_1_2_2((nor_1218_nl), nor_1217_cse, or_2308_nl);
  assign or_2306_nl = FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_3 | (~ inp_lookup_1_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs)
      | IsNaN_6U_10U_5_land_1_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_15;
  assign mux_1008_nl = MUX_s_1_2_2((mux_1007_nl), (and_3222_nl), or_2306_nl);
  assign and_3397_nl = (chn_inp_in_crt_sva_4_739_736_1[0]) & main_stage_v_4 & (cfg_precision_1_sva_st_81==2'b10);
  assign nor_1222_nl = ~((~(nor_1224_cse | (chn_inp_in_crt_sva_4_739_736_1[0])))
      | (~ main_stage_v_4) | (cfg_precision_1_sva_st_81!=2'b10));
  assign mux_1009_nl = MUX_s_1_2_2((nor_1222_nl), nor_1221_cse, inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5);
  assign or_2313_nl = (~ inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5)
      | IsNaN_6U_10U_5_land_1_lpi_1_dfm_6 | FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_4 |
      IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_16;
  assign mux_1010_nl = MUX_s_1_2_2((mux_1009_nl), (and_3397_nl), or_2313_nl);
  assign mux_1011_nl = MUX_s_1_2_2((mux_1010_nl), (mux_1008_nl), or_11_cse);
  assign nor_1215_nl = ~((~ main_stage_v_3) | (~ (chn_inp_in_crt_sva_3_739_736_1[0]))
      | (cfg_precision_1_sva_st_80[0]) | not_tmp_940);
  assign and_3221_nl = inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5
      & (chn_inp_in_crt_sva_4_739_736_1[0]) & (cfg_precision_1_sva_st_81==2'b10);
  assign nor_1216_nl = ~(inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5
      | (~ (chn_inp_in_crt_sva_4_739_736_1[0])) | (cfg_precision_1_sva_st_81!=2'b10));
  assign mux_1013_nl = MUX_s_1_2_2((nor_1216_nl), (and_3221_nl), inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5);
  assign and_3220_nl = main_stage_v_4 & (mux_1013_nl);
  assign mux_1014_nl = MUX_s_1_2_2((and_3220_nl), (nor_1215_nl), or_11_cse);
  assign and_4218_nl = (~ IsNaN_6U_10U_7_land_1_lpi_1_dfm_6) & and_1768_rgt;
  assign nor_1213_nl = ~((~ main_stage_v_3) | (~ (chn_inp_in_crt_sva_3_739_736_1[0]))
      | (cfg_precision_1_sva_st_80[0]) | (~((cfg_precision_1_sva_st_80[1]) & ((~(FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_3
      | IsNaN_6U_10U_5_land_1_lpi_1_dfm_5 | (~ IsNaN_8U_23U_3_IsNaN_8U_23U_3_nor_tmp)))
      | mux_1015_cse))));
  assign mux_1016_nl = MUX_s_1_2_2((~ inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5),
      inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5,
      inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5);
  assign nor_1214_nl = ~((~ main_stage_v_4) | (~ (chn_inp_in_crt_sva_4_739_736_1[0]))
      | (cfg_precision_1_sva_st_81[0]) | (~((cfg_precision_1_sva_st_81[1]) & ((~(IsNaN_6U_10U_5_land_1_lpi_1_dfm_6
      | FpMul_6U_10U_1_lor_6_lpi_1_dfm_6 | (~ FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_4)))
      | (mux_1016_nl)))));
  assign mux_1017_nl = MUX_s_1_2_2((nor_1214_nl), (nor_1213_nl), or_11_cse);
  assign mux_1019_nl = MUX_s_1_2_2(nor_1210_cse, mux_1015_cse, chn_inp_in_crt_sva_3_739_736_1[0]);
  assign nor_1209_nl = ~((~ main_stage_v_3) | (cfg_precision_1_sva_st_80[0]) | (~((cfg_precision_1_sva_st_80[1])
      & (mux_1019_nl))));
  assign mux_1020_nl = MUX_s_1_2_2((~ inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5),
      inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5,
      inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5);
  assign nor_1212_nl = ~(FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_4 | (~ inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5));
  assign mux_1021_nl = MUX_s_1_2_2((nor_1212_nl), (mux_1020_nl), chn_inp_in_crt_sva_4_739_736_1[0]);
  assign nor_1211_nl = ~((~ main_stage_v_4) | (cfg_precision_1_sva_st_81[0]) | (~((cfg_precision_1_sva_st_81[1])
      & (mux_1021_nl))));
  assign mux_1022_nl = MUX_s_1_2_2((nor_1211_nl), (nor_1209_nl), or_11_cse);
  assign FpMul_6U_10U_1_else_2_else_and_1_nl = inp_lookup_2_FpMul_6U_10U_1_else_2_else_if_if_acc_1_itm_5_1
      & (inp_lookup_2_FpMul_6U_10U_1_p_mant_p1_mul_tmp[21]);
  assign and_3218_nl = (chn_inp_in_crt_sva_3_739_736_1[1]) & main_stage_v_3 & (cfg_precision_1_sva_st_80==2'b10);
  assign nor_1201_nl = ~((~((((~ (inp_lookup_2_FpMul_6U_10U_1_p_mant_p1_mul_tmp[21]))
      | inp_lookup_2_FpMul_6U_10U_1_else_2_else_if_if_acc_1_itm_5_1) & inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4)
      | (chn_inp_in_crt_sva_3_739_736_1[1]))) | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10));
  assign or_2345_nl = FpMul_6U_10U_1_lor_7_lpi_1_dfm_5 | inp_lookup_2_FpMantRNE_22U_11U_1_else_and_tmp;
  assign mux_1023_nl = MUX_s_1_2_2((nor_1201_nl), nor_1217_cse, or_2345_nl);
  assign or_2343_nl = FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_3 | (~ inp_lookup_2_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs)
      | IsNaN_6U_10U_5_land_2_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_15;
  assign mux_1024_nl = MUX_s_1_2_2((mux_1023_nl), (and_3218_nl), or_2343_nl);
  assign and_3396_nl = (chn_inp_in_crt_sva_4_739_736_1[1]) & main_stage_v_4 & (cfg_precision_1_sva_st_81==2'b10);
  assign nor_1205_nl = ~((~(nor_1207_cse | (chn_inp_in_crt_sva_4_739_736_1[1])))
      | (~ main_stage_v_4) | (cfg_precision_1_sva_st_81!=2'b10));
  assign mux_1025_nl = MUX_s_1_2_2((nor_1205_nl), nor_1221_cse, inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5);
  assign or_2350_nl = (~ inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5)
      | IsNaN_6U_10U_5_land_2_lpi_1_dfm_6 | FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_4 |
      IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_16;
  assign mux_1026_nl = MUX_s_1_2_2((mux_1025_nl), (and_3396_nl), or_2350_nl);
  assign mux_1027_nl = MUX_s_1_2_2((mux_1026_nl), (mux_1024_nl), or_11_cse);
  assign and_3216_nl = main_stage_v_3 & (chn_inp_in_crt_sva_3_739_736_1[1]) & (~
      mux_tmp_950);
  assign nor_1198_nl = ~((~ inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5)
      | (cfg_precision_1_sva_st_81!=2'b10));
  assign nor_1199_nl = ~(inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5
      | (cfg_precision_1_sva_st_81!=2'b10));
  assign mux_1029_nl = MUX_s_1_2_2((nor_1199_nl), (nor_1198_nl), inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5);
  assign and_3217_nl = main_stage_v_4 & (chn_inp_in_crt_sva_4_739_736_1[1]) & (mux_1029_nl);
  assign mux_1030_nl = MUX_s_1_2_2((and_3217_nl), (and_3216_nl), or_11_cse);
  assign and_4217_nl = (~ IsNaN_6U_10U_7_land_2_lpi_1_dfm_6) & and_1772_rgt;
  assign nor_1196_nl = ~((~ main_stage_v_3) | (~ (chn_inp_in_crt_sva_3_739_736_1[1]))
      | (cfg_precision_1_sva_st_80[0]) | (~((cfg_precision_1_sva_st_80[1]) & ((~(FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_3
      | IsNaN_6U_10U_5_land_2_lpi_1_dfm_5 | (~ IsNaN_8U_23U_3_IsNaN_8U_23U_3_nor_1_tmp)))
      | mux_1031_cse))));
  assign mux_1032_nl = MUX_s_1_2_2((~ inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5),
      inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5,
      inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5);
  assign nor_1197_nl = ~((~ main_stage_v_4) | (~ (chn_inp_in_crt_sva_4_739_736_1[1]))
      | (cfg_precision_1_sva_st_81[0]) | (~((cfg_precision_1_sva_st_81[1]) & ((~(IsNaN_6U_10U_5_land_2_lpi_1_dfm_6
      | FpMul_6U_10U_1_lor_7_lpi_1_dfm_6 | (~ FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_4)))
      | (mux_1032_nl)))));
  assign mux_1033_nl = MUX_s_1_2_2((nor_1197_nl), (nor_1196_nl), or_11_cse);
  assign mux_1035_nl = MUX_s_1_2_2(nor_1193_cse, mux_1031_cse, chn_inp_in_crt_sva_3_739_736_1[1]);
  assign nor_1192_nl = ~((~ main_stage_v_3) | (cfg_precision_1_sva_st_80[0]) | (~((cfg_precision_1_sva_st_80[1])
      & (mux_1035_nl))));
  assign mux_1036_nl = MUX_s_1_2_2((~ inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5),
      inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5,
      inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5);
  assign nor_1195_nl = ~(FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_4 | (~ inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5));
  assign mux_1037_nl = MUX_s_1_2_2((nor_1195_nl), (mux_1036_nl), chn_inp_in_crt_sva_4_739_736_1[1]);
  assign nor_1194_nl = ~((~ main_stage_v_4) | (cfg_precision_1_sva_st_81[0]) | (~((cfg_precision_1_sva_st_81[1])
      & (mux_1037_nl))));
  assign mux_1038_nl = MUX_s_1_2_2((nor_1194_nl), (nor_1192_nl), or_11_cse);
  assign FpMul_6U_10U_1_else_2_else_and_2_nl = inp_lookup_3_FpMul_6U_10U_1_else_2_else_if_if_acc_1_itm_5_1
      & (inp_lookup_3_FpMul_6U_10U_1_p_mant_p1_mul_tmp[21]);
  assign and_3214_nl = (chn_inp_in_crt_sva_3_739_736_1[2]) & main_stage_v_3 & (cfg_precision_1_sva_st_80==2'b10);
  assign nor_1184_nl = ~((~((((~ (inp_lookup_3_FpMul_6U_10U_1_p_mant_p1_mul_tmp[21]))
      | inp_lookup_3_FpMul_6U_10U_1_else_2_else_if_if_acc_1_itm_5_1) & inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4)
      | (chn_inp_in_crt_sva_3_739_736_1[2]))) | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10));
  assign or_2382_nl = FpMul_6U_10U_1_lor_8_lpi_1_dfm_5 | inp_lookup_3_FpMantRNE_22U_11U_1_else_and_tmp;
  assign mux_1039_nl = MUX_s_1_2_2((nor_1184_nl), nor_1217_cse, or_2382_nl);
  assign or_2380_nl = FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_3 | (~ inp_lookup_3_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs)
      | IsNaN_6U_10U_5_land_3_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_15;
  assign mux_1040_nl = MUX_s_1_2_2((mux_1039_nl), (and_3214_nl), or_2380_nl);
  assign and_3395_nl = (chn_inp_in_crt_sva_4_739_736_1[2]) & main_stage_v_4 & (cfg_precision_1_sva_st_81==2'b10);
  assign nor_1188_nl = ~((~(nor_1190_cse | (chn_inp_in_crt_sva_4_739_736_1[2])))
      | (~ main_stage_v_4) | (cfg_precision_1_sva_st_81!=2'b10));
  assign mux_1041_nl = MUX_s_1_2_2((nor_1188_nl), nor_1221_cse, inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5);
  assign or_2387_nl = (~ inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5)
      | IsNaN_6U_10U_5_land_3_lpi_1_dfm_6 | FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_4 |
      IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_16;
  assign mux_1042_nl = MUX_s_1_2_2((mux_1041_nl), (and_3395_nl), or_2387_nl);
  assign mux_1043_nl = MUX_s_1_2_2((mux_1042_nl), (mux_1040_nl), or_11_cse);
  assign and_3212_nl = main_stage_v_3 & (chn_inp_in_crt_sva_3_739_736_1[2]) & (~
      mux_tmp_966);
  assign and_3213_nl = main_stage_v_4 & (chn_inp_in_crt_sva_4_739_736_1[2]) & (~
      mux_tmp_967);
  assign mux_1046_nl = MUX_s_1_2_2((and_3213_nl), (and_3212_nl), or_11_cse);
  assign and_4216_nl = (~ IsNaN_6U_10U_7_land_3_lpi_1_dfm_6) & and_1776_rgt;
  assign mux_1047_nl = MUX_s_1_2_2((~ inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4),
      inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4,
      inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4);
  assign nor_1181_nl = ~((~ main_stage_v_3) | (~ (chn_inp_in_crt_sva_3_739_736_1[2]))
      | (cfg_precision_1_sva_st_80[0]) | (~((cfg_precision_1_sva_st_80[1]) & ((~(FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_3
      | IsNaN_6U_10U_5_land_3_lpi_1_dfm_5 | (~ IsNaN_8U_23U_3_IsNaN_8U_23U_3_nor_2_tmp)))
      | (mux_1047_nl)))));
  assign mux_1048_nl = MUX_s_1_2_2((~ inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5),
      inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5,
      inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5);
  assign nor_1182_nl = ~((~ main_stage_v_4) | (~ (chn_inp_in_crt_sva_4_739_736_1[2]))
      | (cfg_precision_1_sva_st_81[0]) | (~((cfg_precision_1_sva_st_81[1]) & ((~(IsNaN_6U_10U_5_land_3_lpi_1_dfm_6
      | FpMul_6U_10U_1_lor_8_lpi_1_dfm_6 | (~ FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_4)))
      | (mux_1048_nl)))));
  assign mux_1049_nl = MUX_s_1_2_2((nor_1182_nl), (nor_1181_nl), or_11_cse);
  assign or_2410_nl = (~ inp_lookup_3_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs)
      | FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_3 | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_1050_nl = MUX_s_1_2_2((or_2410_nl), mux_tmp_966, chn_inp_in_crt_sva_3_739_736_1[2]);
  assign and_3210_nl = main_stage_v_3 & (~ (mux_1050_nl));
  assign or_2411_nl = FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_4 | (~ inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5)
      | (cfg_precision_1_sva_st_81!=2'b10);
  assign mux_1051_nl = MUX_s_1_2_2((or_2411_nl), mux_tmp_967, chn_inp_in_crt_sva_4_739_736_1[2]);
  assign and_3211_nl = main_stage_v_4 & (~ (mux_1051_nl));
  assign mux_1052_nl = MUX_s_1_2_2((and_3211_nl), (and_3210_nl), or_11_cse);
  assign FpMul_6U_10U_1_else_2_else_and_3_nl = inp_lookup_4_FpMul_6U_10U_1_else_2_else_if_if_acc_1_itm_5_1
      & (inp_lookup_4_FpMul_6U_10U_1_p_mant_p1_mul_tmp[21]);
  assign nand_433_nl = ~(or_5689_cse & inp_lookup_4_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs_2
      & main_stage_v_3 & (cfg_precision_1_sva_st_80==2'b10));
  assign or_2415_nl = FpMul_6U_10U_1_lor_1_lpi_1_dfm_5 | inp_lookup_4_FpMantRNE_22U_11U_1_else_and_tmp;
  assign mux_1053_nl = MUX_s_1_2_2((nand_433_nl), or_2282_cse, or_2415_nl);
  assign or_2418_nl = FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_3 | (~ inp_lookup_4_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs)
      | IsNaN_6U_10U_5_land_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_lpi_1_dfm_st_15 | (mux_1053_nl);
  assign mux_1054_nl = MUX_s_1_2_2((or_2418_nl), or_2282_cse, chn_inp_in_crt_sva_3_739_736_1[3]);
  assign nor_1178_nl = ~(IsNaN_6U_10U_5_land_lpi_1_dfm_6 | FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_4
      | IsNaN_6U_10U_4_land_lpi_1_dfm_5 | (~ inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5));
  assign nor_1179_nl = ~(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_9_1
      | nor_1180_cse | IsNaN_6U_10U_5_land_lpi_1_dfm_6 | FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_4
      | IsNaN_6U_10U_4_land_lpi_1_dfm_5 | (~ inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5));
  assign mux_1055_nl = MUX_s_1_2_2((nor_1179_nl), (nor_1178_nl), inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4);
  assign or_2427_nl = (~ main_stage_v_4) | (cfg_precision_1_sva_st_81!=2'b10) | (~((chn_inp_in_crt_sva_4_739_736_1[3])
      | (mux_1055_nl)));
  assign mux_1056_nl = MUX_s_1_2_2((or_2427_nl), (mux_1054_nl), or_11_cse);
  assign and_4117_nl = (~ IsNaN_6U_10U_7_land_lpi_1_dfm_6) & and_1780_rgt;
  assign nor_1173_nl = ~(nand_661_cse | ((FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_3 | IsNaN_6U_10U_5_land_lpi_1_dfm_5
      | IsNaN_8U_23U_3_IsNaN_8U_23U_3_nand_3_tmp | IsNaN_8U_23U_3_nor_3_tmp) & mux_1061_cse));
  assign mux_1062_nl = MUX_s_1_2_2(inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4,
      (~ inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_4),
      inp_lookup_4_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_5);
  assign nor_1174_nl = ~(nand_579_cse | ((FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_4 | IsNaN_6U_10U_4_land_lpi_1_dfm_5
      | IsNaN_6U_10U_5_land_lpi_1_dfm_6 | IsNaN_8U_23U_2_land_lpi_1_dfm_st_7) & (mux_1062_nl)));
  assign mux_1063_nl = MUX_s_1_2_2((nor_1174_nl), (nor_1173_nl), or_11_cse);
  assign nor_1151_nl = ~((~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[0])
      | (cfg_precision_1_sva_st_81!=2'b10) | (~(IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_tmp
      | FpAdd_6U_10U_1_is_a_greater_acc_itm_6 | inp_lookup_1_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp
      | mux_476_cse)));
  assign or_2520_nl = inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
      | and_tmp_158;
  assign nand_136_nl = ~(inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
      & (~ and_tmp_158));
  assign mux_1090_nl = MUX_s_1_2_2((nand_136_nl), (or_2520_nl), inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6);
  assign nor_1153_nl = ~((chn_inp_in_crt_sva_5_739_736_1[0]) | (cfg_precision_1_sva_st_82[0])
      | (~((cfg_precision_1_sva_st_82[1]) & main_stage_v_5 & (IsNaN_8U_23U_3_land_1_lpi_1_dfm_6
      | IsNaN_6U_10U_8_land_1_lpi_1_dfm_6 | (mux_1090_nl)))));
  assign mux_1091_nl = MUX_s_1_2_2((nor_1153_nl), (nor_1151_nl), or_11_cse);
  assign inp_lookup_1_FpAdd_6U_10U_1_IsZero_6U_10U_8_or_nl = (FpMul_6U_10U_1_o_mant_1_lpi_1_dfm_3!=10'b0000000000)
      | FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_3_5_mx1w1 | FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_3_4_mx1w1
      | (FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_3_3_0_mx1w1!=4'b0000);
  assign nor_1143_nl = ~((~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[1])
      | (cfg_precision_1_sva_st_81!=2'b10) | (~(IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_1_tmp
      | FpAdd_6U_10U_1_is_a_greater_acc_1_itm_6 | inp_lookup_2_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp
      | mux_485_cse)));
  assign or_2557_nl = inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
      | and_tmp_162;
  assign nand_140_nl = ~(inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
      & (~ and_tmp_162));
  assign mux_1107_nl = MUX_s_1_2_2((nand_140_nl), (or_2557_nl), inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6);
  assign nor_1145_nl = ~((~ main_stage_v_5) | (chn_inp_in_crt_sva_5_739_736_1[1])
      | (cfg_precision_1_sva_st_82[0]) | (~((cfg_precision_1_sva_st_82[1]) & (IsNaN_8U_23U_3_land_2_lpi_1_dfm_6
      | IsNaN_6U_10U_8_land_2_lpi_1_dfm_4 | (mux_1107_nl)))));
  assign mux_1108_nl = MUX_s_1_2_2((nor_1145_nl), (nor_1143_nl), or_11_cse);
  assign inp_lookup_2_FpAdd_6U_10U_1_IsZero_6U_10U_8_or_nl = (FpMul_6U_10U_1_o_mant_2_lpi_1_dfm_3!=10'b0000000000)
      | FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_3_5_mx1w1 | FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_3_4_mx1w1
      | (FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_3_3_0_mx1w1!=4'b0000);
  assign nor_1135_nl = ~((~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[2])
      | (cfg_precision_1_sva_st_81!=2'b10) | (~(IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_2_tmp
      | FpAdd_6U_10U_1_is_a_greater_acc_2_itm_6 | inp_lookup_3_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp
      | mux_500_cse)));
  assign or_2594_nl = inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
      | and_tmp_166;
  assign nand_144_nl = ~(inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
      & (~ and_tmp_166));
  assign mux_1124_nl = MUX_s_1_2_2((nand_144_nl), (or_2594_nl), inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6);
  assign nor_1137_nl = ~((~ main_stage_v_5) | (chn_inp_in_crt_sva_5_739_736_1[2])
      | (cfg_precision_1_sva_st_82[0]) | (~((cfg_precision_1_sva_st_82[1]) & (IsNaN_8U_23U_3_land_3_lpi_1_dfm_6
      | IsNaN_6U_10U_8_land_3_lpi_1_dfm_4 | (mux_1124_nl)))));
  assign mux_1125_nl = MUX_s_1_2_2((nor_1137_nl), (nor_1135_nl), or_11_cse);
  assign inp_lookup_3_FpAdd_6U_10U_1_IsZero_6U_10U_8_or_nl = (FpMul_6U_10U_1_o_mant_3_lpi_1_dfm_3_mx0w1!=10'b0000000000)
      | FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_5_mx1w1 | FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_4_mx1w1
      | (FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_3_3_0_mx1w1!=4'b0000);
  assign nor_1127_nl = ~((~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[3])
      | (cfg_precision_1_sva_st_81!=2'b10) | (~(IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_3_tmp
      | FpAdd_6U_10U_1_is_a_greater_acc_3_itm_6_1 | inp_lookup_4_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp
      | mux_1140_cse)));
  assign or_2632_nl = nor_1130_cse | mux_tmp_1059;
  assign mux_1142_nl = MUX_s_1_2_2(mux_tmp_1059, (or_2632_nl), IsNaN_8U_23U_2_land_lpi_1_dfm_9);
  assign nor_1129_nl = ~((~ main_stage_v_5) | (chn_inp_in_crt_sva_5_739_736_1[3])
      | (cfg_precision_1_sva_st_82[0]) | (~((cfg_precision_1_sva_st_82[1]) & (IsNaN_8U_23U_3_land_lpi_1_dfm_5
      | IsNaN_6U_10U_8_land_lpi_1_dfm_4 | (mux_1142_nl)))));
  assign mux_1143_nl = MUX_s_1_2_2((nor_1129_nl), (nor_1127_nl), or_11_cse);
  assign inp_lookup_4_FpAdd_6U_10U_1_IsZero_6U_10U_8_or_nl = (FpMul_6U_10U_1_o_mant_lpi_1_dfm_3_mx0w0!=10'b0000000000)
      | FpMul_6U_10U_1_o_expo_lpi_1_dfm_3_5_mx0w1 | FpMul_6U_10U_1_o_expo_lpi_1_dfm_3_4_mx0w1
      | (FpMul_6U_10U_1_o_expo_lpi_1_dfm_3_3_0_mx0w1!=4'b0000);
  assign nor_1123_nl = ~(((nor_126_cse | IsNaN_8U_23U_2_land_1_lpi_1_dfm_9 | IsNaN_8U_23U_2_land_1_lpi_1_dfm_st_7
      | IsNaN_8U_23U_3_land_1_lpi_1_dfm_6) & (chn_inp_in_crt_sva_5_739_736_1[0]))
      | (cfg_precision_1_sva_st_82[0]) | not_tmp_374);
  assign or_2650_nl = (~ inp_lookup_1_FpMantRNE_49U_24U_1_else_and_tmp) | inp_lookup_1_FpAdd_8U_23U_1_if_4_if_acc_1_itm_7_1;
  assign mux_1154_nl = MUX_s_1_2_2(nor_1124_cse, (nor_1123_nl), or_2650_nl);
  assign nor_1125_nl = ~((chn_inp_in_crt_sva_6_739_736_1[0]) | (cfg_precision_1_sva_st_83!=2'b10)
      | (~ main_stage_v_6));
  assign nor_1126_nl = ~((~(FpMul_6U_10U_1_o_expo_1_lpi_1_dfm_7_4_1 | (~ inp_lookup_1_FpMantRNE_49U_24U_1_else_and_svs_2)
      | (~ (chn_inp_in_crt_sva_6_739_736_1[0])))) | (cfg_precision_1_sva_st_83!=2'b10)
      | (~ main_stage_v_6));
  assign or_2656_nl = IsNaN_8U_23U_3_land_1_lpi_1_dfm_7 | FpAdd_6U_10U_1_is_a_greater_lor_1_lpi_1_dfm_5
      | IsNaN_6U_10U_8_land_1_lpi_1_dfm_st_3 | IsNaN_6U_10U_9_land_1_lpi_1_dfm_7;
  assign mux_1155_nl = MUX_s_1_2_2((nor_1126_nl), (nor_1125_nl), or_2656_nl);
  assign mux_1156_nl = MUX_s_1_2_2((mux_1155_nl), (mux_1154_nl), or_11_cse);
  assign mux_1157_nl = MUX_s_1_2_2(or_tmp_1098, or_tmp_2486, or_11_cse);
  assign nor_1119_nl = ~(((FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_1_cse | IsNaN_8U_23U_3_land_2_lpi_1_dfm_6
      | IsNaN_8U_23U_2_land_2_lpi_1_dfm_st_7 | IsNaN_8U_23U_2_land_2_lpi_1_dfm_9)
      & (chn_inp_in_crt_sva_5_739_736_1[1])) | (cfg_precision_1_sva_st_82!=2'b10)
      | (~ main_stage_v_5));
  assign nor_1120_nl = ~((chn_inp_in_crt_sva_5_739_736_1[1]) | (cfg_precision_1_sva_st_82!=2'b10)
      | (~ main_stage_v_5));
  assign mux_1158_nl = MUX_s_1_2_2((nor_1120_nl), (nor_1119_nl), or_2663_cse);
  assign nor_1121_nl = ~((chn_inp_in_crt_sva_6_739_736_1[1]) | (cfg_precision_1_sva_st_83[0])
      | nand_570_cse);
  assign nor_1122_nl = ~((~(FpMul_6U_10U_1_o_expo_2_lpi_1_dfm_7_4_1 | (~ inp_lookup_2_FpMantRNE_49U_24U_1_else_and_svs_2)
      | (~ (chn_inp_in_crt_sva_6_739_736_1[1])))) | (cfg_precision_1_sva_st_83[0])
      | nand_570_cse);
  assign or_2669_nl = IsNaN_8U_23U_3_land_2_lpi_1_dfm_7 | FpAdd_6U_10U_1_is_a_greater_lor_2_lpi_1_dfm_5
      | IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_4 | IsNaN_6U_10U_9_land_2_lpi_1_dfm_7;
  assign mux_1159_nl = MUX_s_1_2_2((nor_1122_nl), (nor_1121_nl), or_2669_nl);
  assign mux_1160_nl = MUX_s_1_2_2((mux_1159_nl), (mux_1158_nl), or_11_cse);
  assign mux_1161_nl = MUX_s_1_2_2(or_tmp_1143, or_tmp_2490, or_11_cse);
  assign and_3198_nl = (FpAdd_8U_23U_1_FpAdd_8U_23U_1_nor_2_cse | IsNaN_8U_23U_2_land_3_lpi_1_dfm_st_7
      | IsNaN_8U_23U_2_land_3_lpi_1_dfm_9 | IsNaN_8U_23U_3_land_3_lpi_1_dfm_6) &
      (chn_inp_in_crt_sva_5_739_736_1[2]);
  assign mux_1162_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_5_739_736_1[2]), (and_3198_nl),
      or_2676_cse);
  assign nor_1116_nl = ~((cfg_precision_1_sva_st_82!=2'b10) | (~ main_stage_v_5)
      | (mux_1162_nl));
  assign nor_1117_nl = ~((chn_inp_in_crt_sva_6_739_736_1[2]) | (cfg_precision_1_sva_st_83!=2'b10)
      | (~ main_stage_v_6));
  assign nor_1118_nl = ~((~(FpMul_6U_10U_1_o_expo_3_lpi_1_dfm_7_4_1 | (~ reg_inp_lookup_3_FpMantRNE_49U_24U_1_else_and_svs_1_cse)
      | (~ (chn_inp_in_crt_sva_6_739_736_1[2])))) | (cfg_precision_1_sva_st_83!=2'b10)
      | (~ main_stage_v_6));
  assign or_2678_nl = IsNaN_8U_23U_3_land_3_lpi_1_dfm_7 | FpAdd_6U_10U_1_is_a_greater_lor_3_lpi_1_dfm_5
      | IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_4 | IsNaN_6U_10U_9_land_3_lpi_1_dfm_7;
  assign mux_1163_nl = MUX_s_1_2_2((nor_1118_nl), (nor_1117_nl), or_2678_nl);
  assign mux_1164_nl = MUX_s_1_2_2((mux_1163_nl), (nor_1116_nl), or_11_cse);
  assign mux_1165_nl = MUX_s_1_2_2(or_tmp_1185, or_tmp_2494, or_11_cse);
  assign nor_1112_nl = ~(((nor_136_cse | IsNaN_8U_23U_2_land_lpi_1_dfm_9 | IsNaN_8U_23U_2_land_lpi_1_dfm_st_8
      | IsNaN_8U_23U_3_land_lpi_1_dfm_5) & (chn_inp_in_crt_sva_5_739_736_1[3])) |
      (cfg_precision_1_sva_st_82[0]) | not_tmp_374);
  assign or_2685_nl = (~ inp_lookup_4_FpMantRNE_49U_24U_1_else_and_tmp) | inp_lookup_4_FpAdd_8U_23U_1_if_4_if_acc_1_itm_7_1;
  assign mux_1166_nl = MUX_s_1_2_2(nor_1113_cse, (nor_1112_nl), or_2685_nl);
  assign nor_1114_nl = ~((chn_inp_in_crt_sva_6_739_736_1[3]) | (~ (cfg_precision_1_sva_st_83[1]))
      | (~ main_stage_v_6) | (cfg_precision_1_sva_st_83[0]));
  assign nor_1115_nl = ~((~(FpMul_6U_10U_1_o_expo_lpi_1_dfm_7_4_1 | (~ inp_lookup_4_FpMantRNE_49U_24U_1_else_and_svs_2)
      | (~ (chn_inp_in_crt_sva_6_739_736_1[3])))) | (~ (cfg_precision_1_sva_st_83[1]))
      | (~ main_stage_v_6) | (cfg_precision_1_sva_st_83[0]));
  assign or_2691_nl = IsNaN_8U_23U_3_land_lpi_1_dfm_6 | FpAdd_6U_10U_1_is_a_greater_lor_lpi_1_dfm_5
      | IsNaN_6U_10U_8_land_lpi_1_dfm_st_4 | IsNaN_6U_10U_9_land_lpi_1_dfm_7;
  assign mux_1167_nl = MUX_s_1_2_2((nor_1115_nl), (nor_1114_nl), or_2691_nl);
  assign mux_1168_nl = MUX_s_1_2_2((mux_1167_nl), (mux_1166_nl), or_11_cse);
  assign mux_1169_nl = MUX_s_1_2_2(or_tmp_1239, or_tmp_2498, or_11_cse);
  assign nl_inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_nl = conv_u2u_4_5({FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_i_shift_acc_psp_4_sva_mx0w0
      , (~ (FpAdd_8U_23U_1_o_expo_3_lpi_1_dfm_7[0]))}) + 5'b1101;
  assign inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_nl = nl_inp_lookup_3_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_nl[4:0];
  assign and_3192_nl = or_tmp_1060 & inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8
      & (~ inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7) & inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8;
  assign mux_1183_nl = MUX_s_1_2_2(or_tmp_2723, (and_3192_nl), chn_inp_in_crt_sva_6_739_736_1[0]);
  assign and_3191_nl = (~((~ main_stage_v_6) | (cfg_precision_1_sva_st_83!=2'b10)))
      & (mux_1183_nl);
  assign and_3193_nl = FpAdd_6U_10U_1_or_12_cse & (~((((~ inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_2)
      | inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2
      | (~ inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2)
      | inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
      | (~ inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2))
      & (chn_inp_in_crt_sva_7_739_736_1[0])) | (~ main_stage_v_7) | (cfg_precision_1_sva_st_84!=2'b10)));
  assign mux_1184_nl = MUX_s_1_2_2((and_3193_nl), (and_3191_nl), or_11_cse);
  assign mux_2119_nl = MUX_s_1_2_2(or_tmp_4741, (~ or_5683_itm), inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8);
  assign or_6080_nl = inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8
      | inp_lookup_1_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7;
  assign mux_2120_nl = MUX_s_1_2_2((mux_2119_nl), or_tmp_4741, or_6080_nl);
  assign nor_1101_nl = ~((~ inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8)
      | inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7 | (~ inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8)
      | IsNaN_8U_23U_4_IsNaN_8U_23U_4_nor_1_tmp | (~ main_stage_v_6) | (cfg_precision_1_sva_st_83!=2'b10));
  assign and_3380_nl = or_tmp_2738 & main_stage_v_6 & (cfg_precision_1_sva_st_83==2'b10);
  assign mux_1188_nl = MUX_s_1_2_2((and_3380_nl), (nor_1101_nl), chn_inp_in_crt_sva_6_739_736_1[1]);
  assign nor_1103_nl = ~(((inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2
      | (~ inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2)
      | inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
      | (~ inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2)
      | IsNaN_6U_10U_8_land_2_lpi_1_dfm_st_5) & (chn_inp_in_crt_sva_7_739_736_1[1]))
      | (~ main_stage_v_7) | (cfg_precision_1_sva_st_84!=2'b10));
  assign nor_1104_nl = ~((~ IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_19) | (chn_inp_in_crt_sva_7_739_736_1[1])
      | (~ main_stage_v_7) | (cfg_precision_1_sva_st_84!=2'b10));
  assign mux_1189_nl = MUX_s_1_2_2((nor_1104_nl), (nor_1103_nl), IsNaN_6U_10U_9_land_2_lpi_1_dfm_8);
  assign mux_1190_nl = MUX_s_1_2_2((mux_1189_nl), (mux_1188_nl), or_11_cse);
  assign mux_2121_nl = MUX_s_1_2_2(or_tmp_4745, (~ or_5684_itm), inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8);
  assign or_6087_nl = inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8
      | inp_lookup_2_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7;
  assign mux_2122_nl = MUX_s_1_2_2((mux_2121_nl), or_tmp_4745, or_6087_nl);
  assign nor_1094_nl = ~((~ inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8)
      | inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7 | (~ inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8)
      | IsNaN_8U_23U_4_IsNaN_8U_23U_4_nor_2_tmp | (~ main_stage_v_6) | (cfg_precision_1_sva_st_83!=2'b10));
  assign and_3378_nl = or_tmp_2703 & main_stage_v_6 & (cfg_precision_1_sva_st_83==2'b10);
  assign mux_1194_nl = MUX_s_1_2_2((and_3378_nl), (nor_1094_nl), chn_inp_in_crt_sva_6_739_736_1[2]);
  assign nor_1096_nl = ~(((inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2
      | (~ inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2)
      | inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
      | (~ inp_lookup_3_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2)
      | IsNaN_6U_10U_8_land_3_lpi_1_dfm_st_5) & (chn_inp_in_crt_sva_7_739_736_1[2]))
      | (~ main_stage_v_7) | (cfg_precision_1_sva_st_84!=2'b10));
  assign nor_1097_nl = ~((~ IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_19) | (chn_inp_in_crt_sva_7_739_736_1[2])
      | (~ main_stage_v_7) | (cfg_precision_1_sva_st_84!=2'b10));
  assign mux_1195_nl = MUX_s_1_2_2((nor_1097_nl), (nor_1096_nl), IsNaN_6U_10U_9_land_3_lpi_1_dfm_8);
  assign mux_1196_nl = MUX_s_1_2_2((mux_1195_nl), (mux_1194_nl), or_11_cse);
  assign or_2773_nl = (cfg_precision_1_sva_st_84!=2'b10) | (~(IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_19
      & main_stage_v_7));
  assign or_2771_nl = IsNaN_6U_10U_9_land_3_lpi_1_dfm_8 | (chn_inp_in_crt_sva_7_739_736_1[2]);
  assign mux_1197_nl = MUX_s_1_2_2((or_2773_nl), or_tmp_1182, or_2771_nl);
  assign mux_1198_nl = MUX_s_1_2_2((mux_1197_nl), or_tmp_2768, or_11_cse);
  assign nor_1090_nl = ~((~ inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8)
      | inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7 | (~ inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8)
      | IsNaN_8U_23U_4_IsNaN_8U_23U_4_nor_3_tmp | (~ main_stage_v_6) | (cfg_precision_1_sva_st_83!=2'b10));
  assign and_3377_nl = or_tmp_2695 & main_stage_v_6 & (cfg_precision_1_sva_st_83==2'b10);
  assign mux_1199_nl = MUX_s_1_2_2((and_3377_nl), (nor_1090_nl), chn_inp_in_crt_sva_6_739_736_1[3]);
  assign nor_1092_nl = ~(((inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs_2
      | (~ inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_8_svs_2)
      | inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_7_svs
      | (~ inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_if_slc_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_8_svs_st_2)
      | IsNaN_6U_10U_8_land_lpi_1_dfm_st_5) & (chn_inp_in_crt_sva_7_739_736_1[3]))
      | (~ main_stage_v_7) | (cfg_precision_1_sva_st_84!=2'b10));
  assign nor_1093_nl = ~((~ IsNaN_6U_10U_2_land_lpi_1_dfm_st_18) | (chn_inp_in_crt_sva_7_739_736_1[3])
      | (~ main_stage_v_7) | (cfg_precision_1_sva_st_84!=2'b10));
  assign mux_1200_nl = MUX_s_1_2_2((nor_1093_nl), (nor_1092_nl), IsNaN_6U_10U_9_land_lpi_1_dfm_8);
  assign mux_1201_nl = MUX_s_1_2_2((mux_1200_nl), (mux_1199_nl), or_11_cse);
  assign nor_1866_nl = ~((chn_inp_in_crt_sva_6_739_736_1[3]) | IsNaN_6U_10U_9_land_lpi_1_dfm_7
      | IsNaN_6U_10U_2_land_lpi_1_dfm_st_17);
  assign mux_2125_nl = MUX_s_1_2_2(or_tmp_4753, (nor_1866_nl), inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_acc_itm_8);
  assign or_6101_nl = inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_else_acc_itm_8
      | inp_lookup_4_FpWidthDec_8U_23U_6U_10U_0U_1U_else_if_acc_itm_7;
  assign mux_2126_nl = MUX_s_1_2_2((mux_2125_nl), or_tmp_4753, or_6101_nl);
  assign IsNaN_6U_23U_2_IsNaN_6U_23U_2_nand_nl = ~(FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_5_mx0w0
      & FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_4_mx0w0 & (FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_7_3_0_mx0w0==4'b1111));
  assign IsNaN_6U_23U_2_IsNaN_6U_23U_2_nand_1_nl = ~(FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_5_mx0w0
      & FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_4_mx0w0 & (FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_7_3_0_mx0w0==4'b1111));
  assign IsNaN_6U_23U_2_IsNaN_6U_23U_2_nand_2_nl = ~(FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_5_mx0w0
      & FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_4_mx0w0 & (FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_7_3_0_mx0w0==4'b1111));
  assign IsNaN_6U_23U_2_IsNaN_6U_23U_2_nand_3_nl = ~(FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_5_mx0w0
      & FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_4_mx0w0 & (FpAdd_6U_10U_1_o_expo_lpi_1_dfm_7_3_0_mx0w0==4'b1111));
  assign and_3184_nl = (~((~((~ IsNaN_6U_10U_IsNaN_6U_10U_nor_tmp) & inp_lookup_1_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp
      & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_12_1_1 & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_12_0_1
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_21==4'b1111))) & FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_tmp))
      & (chn_inp_in_crt_sva_7_739_736_1[0]) & (cfg_precision_1_sva_st_84[1]) & main_stage_v_7
      & (~ (cfg_precision_1_sva_st_84[0]));
  assign and_3375_nl = main_stage_v_8 & (chn_inp_in_crt_sva_8_739_736_1[0]) & (cfg_precision_1_sva_st_85==2'b10);
  assign mux_1207_nl = MUX_s_1_2_2((and_3375_nl), nor_1490_cse, or_2797_cse);
  assign mux_1208_nl = MUX_s_1_2_2((mux_1207_nl), (and_3184_nl), or_11_cse);
  assign or_2805_nl = (~(IsNaN_6U_10U_IsNaN_6U_10U_nor_1_tmp | (~ FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_2_tmp)))
      | (cfg_precision_1_sva_st_84[0]) | (~ and_dcpl_21);
  assign mux_1210_nl = MUX_s_1_2_2(or_tmp_1302, or_tmp_2804, reg_FpMul_6U_10U_lor_4_lpi_1_dfm_3_cse);
  assign mux_1211_nl = MUX_s_1_2_2((mux_1210_nl), (or_2805_nl), or_11_cse);
  assign nor_1082_nl = ~(((~((~ IsNaN_6U_10U_IsNaN_6U_10U_nor_1_tmp) & inp_lookup_2_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp
      & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_12_1_1 & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_12_0_1
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_21==4'b1111))) & FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_2_tmp)
      | (cfg_precision_1_sva_st_84[0]) | (~((cfg_precision_1_sva_st_84[1]) & main_stage_v_7
      & (chn_inp_in_crt_sva_7_739_736_1[1]))));
  assign mux_1212_nl = MUX_s_1_2_2(and_3374_cse, nor_1488_cse, or_2810_cse);
  assign mux_1213_nl = MUX_s_1_2_2((mux_1212_nl), (nor_1082_nl), or_11_cse);
  assign and_3182_nl = (~((~((~ IsNaN_6U_10U_IsNaN_6U_10U_nor_3_tmp) & inp_lookup_4_IsNaN_6U_10U_1_aif_IsNaN_6U_10U_1_aelse_IsNaN_6U_10U_1_aelse_or_tmp
      & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_12_1_1 & FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_12_0_1
      & (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_21==4'b1111))) & FpMul_6U_10U_if_2_FpMul_6U_10U_if_2_or_6_tmp))
      & (chn_inp_in_crt_sva_7_739_736_1[3]) & (cfg_precision_1_sva_st_84[1]) & main_stage_v_7
      & (~ (cfg_precision_1_sva_st_84[0]));
  assign and_3373_nl = main_stage_v_8 & (chn_inp_in_crt_sva_8_739_736_1[3]) & (cfg_precision_1_sva_st_85==2'b10);
  assign mux_1218_nl = MUX_s_1_2_2((and_3373_nl), nor_1469_cse, or_2822_cse);
  assign mux_1219_nl = MUX_s_1_2_2((mux_1218_nl), (and_3182_nl), or_11_cse);
  assign nor_1078_nl = ~((~ (chn_inp_in_crt_sva_8_739_736_1[0])) | (cfg_precision_1_sva_st_85!=2'b10)
      | (~(or_tmp_1363 & main_stage_v_8)));
  assign and_3181_nl = (chn_inp_in_crt_sva_9_739_736_1[0]) & or_tmp_1369 & main_stage_v_9
      & (cfg_precision_1_sva_st_86==2'b10);
  assign mux_1220_nl = MUX_s_1_2_2((and_3181_nl), (nor_1078_nl), or_11_cse);
  assign nand_676_nl = ~((chn_inp_in_crt_sva_9_739_736_1[0]) & IsNaN_6U_10U_land_1_lpi_1_dfm_6
      & main_stage_v_9 & (cfg_precision_1_sva_st_86==2'b10));
  assign mux_1222_nl = MUX_s_1_2_2((nand_676_nl), or_tmp_1253, or_11_cse);
  assign nor_1074_nl = ~((~ (chn_inp_in_crt_sva_8_739_736_1[0])) | (cfg_precision_1_sva_st_85!=2'b10)
      | IsNaN_6U_10U_1_land_1_lpi_1_dfm_5 | IsNaN_6U_10U_land_1_lpi_1_dfm_5 | (~
      main_stage_v_8));
  assign nor_1075_nl = ~((~ (chn_inp_in_crt_sva_9_739_736_1[0])) | IsNaN_6U_10U_land_1_lpi_1_dfm_6
      | IsNaN_6U_10U_1_land_1_lpi_1_dfm_6 | (~ main_stage_v_9) | (cfg_precision_1_sva_st_86!=2'b10));
  assign mux_1223_nl = MUX_s_1_2_2((nor_1075_nl), (nor_1074_nl), or_11_cse);
  assign nor_1072_nl = ~((cfg_precision_1_sva_st_85[0]) | (~((cfg_precision_1_sva_st_85[1])
      & (chn_inp_in_crt_sva_8_739_736_1[1]) & or_tmp_1393 & main_stage_v_8)));
  assign and_3180_nl = (chn_inp_in_crt_sva_9_739_736_1[1]) & or_tmp_1399 & main_stage_v_9
      & (cfg_precision_1_sva_st_100==2'b10);
  assign mux_1224_nl = MUX_s_1_2_2((and_3180_nl), (nor_1072_nl), or_11_cse);
  assign nand_674_nl = ~((chn_inp_in_crt_sva_9_739_736_1[1]) & IsNaN_6U_10U_land_2_lpi_1_dfm_6
      & main_stage_v_9 & (cfg_precision_1_sva_st_100==2'b10));
  assign mux_1226_nl = MUX_s_1_2_2((nand_674_nl), or_tmp_2804, or_11_cse);
  assign nor_1068_nl = ~((cfg_precision_1_sva_st_85!=2'b10) | (~ (chn_inp_in_crt_sva_8_739_736_1[1]))
      | IsNaN_6U_10U_1_land_2_lpi_1_dfm_5 | IsNaN_6U_10U_land_2_lpi_1_dfm_5 | (~
      main_stage_v_8));
  assign nor_1069_nl = ~((~ (chn_inp_in_crt_sva_9_739_736_1[1])) | IsNaN_6U_10U_land_2_lpi_1_dfm_6
      | IsNaN_6U_10U_1_land_2_lpi_1_dfm_6 | (~ main_stage_v_9) | (cfg_precision_1_sva_st_100!=2'b10));
  assign mux_1227_nl = MUX_s_1_2_2((nor_1069_nl), (nor_1068_nl), or_11_cse);
  assign and_3178_nl = (chn_inp_in_crt_sva_8_739_736_1[2]) & or_tmp_1422 & (cfg_precision_1_sva_st_85==2'b10)
      & main_stage_v_8;
  assign and_3179_nl = (chn_inp_in_crt_sva_9_739_736_1[2]) & or_tmp_1428 & main_stage_v_9
      & (cfg_precision_1_sva_st_112==2'b10);
  assign mux_1228_nl = MUX_s_1_2_2((and_3179_nl), (and_3178_nl), or_11_cse);
  assign nand_672_nl = ~((chn_inp_in_crt_sva_9_739_736_1[2]) & IsNaN_6U_10U_land_3_lpi_1_dfm_6
      & main_stage_v_9 & (cfg_precision_1_sva_st_112==2'b10));
  assign mux_1230_nl = MUX_s_1_2_2((nand_672_nl), or_tmp_1310, or_11_cse);
  assign nor_1063_nl = ~((~ (chn_inp_in_crt_sva_8_739_736_1[2])) | IsNaN_6U_10U_1_land_3_lpi_1_dfm_5
      | IsNaN_6U_10U_land_3_lpi_1_dfm_5 | (cfg_precision_1_sva_st_85!=2'b10) | (~
      main_stage_v_8));
  assign nor_1064_nl = ~((~ (chn_inp_in_crt_sva_9_739_736_1[2])) | IsNaN_6U_10U_land_3_lpi_1_dfm_6
      | IsNaN_6U_10U_1_land_3_lpi_1_dfm_6 | (~ main_stage_v_9) | (cfg_precision_1_sva_st_112!=2'b10));
  assign mux_1231_nl = MUX_s_1_2_2((nor_1064_nl), (nor_1063_nl), or_11_cse);
  assign and_3176_nl = (chn_inp_in_crt_sva_8_739_736_1[3]) & or_tmp_1448 & (cfg_precision_1_sva_st_85==2'b10)
      & main_stage_v_8;
  assign and_3177_nl = (chn_inp_in_crt_sva_9_739_736_1[3]) & or_tmp_1454 & main_stage_v_9
      & (cfg_precision_1_sva_st_124==2'b10);
  assign mux_1232_nl = MUX_s_1_2_2((and_3177_nl), (and_3176_nl), or_11_cse);
  assign nand_390_nl = ~((chn_inp_in_crt_sva_9_739_736_1[3]) & IsNaN_6U_10U_land_lpi_1_dfm_6
      & main_stage_v_9 & (cfg_precision_1_sva_st_124==2'b10));
  assign mux_1234_nl = MUX_s_1_2_2((nand_390_nl), or_tmp_1338, or_11_cse);
  assign nor_1059_nl = ~((~ (chn_inp_in_crt_sva_8_739_736_1[3])) | IsNaN_6U_10U_1_land_lpi_1_dfm_5
      | IsNaN_6U_10U_land_lpi_1_dfm_5 | (cfg_precision_1_sva_st_85!=2'b10) | (~ main_stage_v_8));
  assign nor_1060_nl = ~((~ (chn_inp_in_crt_sva_9_739_736_1[3])) | IsNaN_6U_10U_land_lpi_1_dfm_6
      | IsNaN_6U_10U_1_land_lpi_1_dfm_6 | (~ main_stage_v_9) | (cfg_precision_1_sva_st_124!=2'b10));
  assign mux_1235_nl = MUX_s_1_2_2((nor_1060_nl), (nor_1059_nl), or_11_cse);
  assign or_2930_nl = (~ (chn_inp_in_crt_sva_10_739_736_1[3])) | (cfg_precision_1_sva_st_125!=2'b10)
      | (~(((~(IsNaN_6U_10U_2_land_lpi_1_dfm_st_21 | (~ IsNaN_6U_10U_3_land_lpi_1_dfm_6)))
      | IsNaN_6U_10U_2_land_lpi_1_dfm_24) & main_stage_v_10));
  assign mux_1246_nl = MUX_s_1_2_2(mux_tmp_754, (or_2930_nl), or_11_cse);
  assign nor_1049_nl = ~((~ main_stage_v_10) | (~ (chn_inp_in_crt_sva_10_739_736_1[2]))
      | (cfg_precision_1_sva_st_113[0]) | (~((cfg_precision_1_sva_st_113[1]) & ((~(IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_22
      | (~ IsNaN_6U_10U_3_land_3_lpi_1_dfm_6))) | IsNaN_6U_10U_2_land_3_lpi_1_dfm_24))));
  assign mux_1249_nl = MUX_s_1_2_2(nor_1397_cse, (nor_1049_nl), or_11_cse);
  assign nor_1046_nl = ~((~ main_stage_v_10) | (~ (chn_inp_in_crt_sva_10_739_736_1[1]))
      | (cfg_precision_1_sva_st_101[0]) | (~((cfg_precision_1_sva_st_101[1]) & ((~(IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_22
      | (~ IsNaN_6U_10U_3_land_2_lpi_1_dfm_6))) | IsNaN_6U_10U_2_land_2_lpi_1_dfm_24))));
  assign mux_1253_nl = MUX_s_1_2_2(nor_1407_cse, (nor_1046_nl), or_11_cse);
  assign nor_1042_nl = ~((cfg_precision_1_sva_st_87[0]) | (~((cfg_precision_1_sva_st_87[1])
      & IsNaN_6U_10U_2_land_1_lpi_1_dfm_24 & main_stage_v_10)));
  assign nor_1043_nl = ~((cfg_precision_1_sva_st_87[0]) | not_tmp_1212);
  assign mux_1258_nl = MUX_s_1_2_2((nor_1043_nl), (nor_1042_nl), IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_22);
  assign nand_166_nl = ~((chn_inp_in_crt_sva_10_739_736_1[0]) & (mux_1258_nl));
  assign mux_1259_nl = MUX_s_1_2_2(mux_tmp_708, (nand_166_nl), or_11_cse);
  assign mux_1262_nl = MUX_s_1_2_2(nor_tmp_234, and_tmp_182, or_11_cse);
  assign and_284_nl = or_11_cse & (chn_inp_in_crt_sva_10_739_736_1[3]) & mux_tmp_1183;
  assign mux_1263_nl = MUX_s_1_2_2((and_284_nl), (mux_1262_nl), inp_lookup_if_unequal_tmp_12);
  assign mux_1266_nl = MUX_s_1_2_2(nor_tmp_232, and_tmp_184, or_11_cse);
  assign and_286_nl = or_11_cse & (chn_inp_in_crt_sva_10_739_736_1[2]) & mux_tmp_1187;
  assign mux_1267_nl = MUX_s_1_2_2((and_286_nl), (mux_1266_nl), inp_lookup_if_unequal_tmp_12);
  assign mux_1271_nl = MUX_s_1_2_2(nor_tmp_253, and_tmp_187, or_11_cse);
  assign mux_1274_nl = MUX_s_1_2_2(nor_tmp_227, and_tmp_188, or_11_cse);
  assign and_290_nl = or_11_cse & (chn_inp_in_crt_sva_10_739_736_1[0]) & mux_tmp_1195;
  assign mux_1275_nl = MUX_s_1_2_2((and_290_nl), (mux_1274_nl), inp_lookup_if_unequal_tmp_12);
  assign mux_1264_nl = MUX_s_1_2_2(or_tmp_1826, or_tmp_2986, or_11_cse);
  assign mux_1268_nl = MUX_s_1_2_2(or_tmp_1849, or_tmp_2990, or_11_cse);
  assign mux_1272_nl = MUX_s_1_2_2(or_tmp_1840, or_tmp_2993, or_11_cse);
  assign mux_1276_nl = MUX_s_1_2_2(or_tmp_1818, or_tmp_2997, or_11_cse);
  assign nor_1040_nl = ~((cfg_precision_1_sva_st_86[1]) | (~ or_tmp_2999));
  assign mux_2192_nl = MUX_s_1_2_2((nor_1040_nl), or_tmp_2999, cfg_precision_1_sva_st_86[0]);
  assign and_3173_nl = main_stage_v_9 & (~((mux_2192_nl) | (~ (chn_inp_in_crt_sva_9_739_736_1[0]))));
  assign nor_1041_nl = ~((cfg_precision_1_sva_st_87[1]) | (~ or_tmp_3002));
  assign mux_2197_nl = MUX_s_1_2_2((nor_1041_nl), or_tmp_3002, cfg_precision_1_sva_st_87[0]);
  assign and_3174_nl = main_stage_v_10 & (~((mux_2197_nl) | (~ (chn_inp_in_crt_sva_10_739_736_1[0]))));
  assign mux_1281_nl = MUX_s_1_2_2((and_3174_nl), (and_3173_nl), or_11_cse);
  assign nor_1038_nl = ~((cfg_precision_1_sva_st_86[1]) | (~ or_tmp_3007));
  assign mux_1282_nl = MUX_s_1_2_2((nor_1038_nl), or_tmp_3007, cfg_precision_1_sva_st_86[0]);
  assign and_3171_nl = main_stage_v_9 & (~ (mux_1282_nl)) & (chn_inp_in_crt_sva_9_739_736_1[0]);
  assign nor_1039_nl = ~((cfg_precision_1_sva_st_87[1]) | (~ or_tmp_3011));
  assign mux_1284_nl = MUX_s_1_2_2((nor_1039_nl), or_tmp_3011, cfg_precision_1_sva_st_87[0]);
  assign and_3172_nl = main_stage_v_10 & (~ (mux_1284_nl)) & (chn_inp_in_crt_sva_10_739_736_1[0]);
  assign mux_1286_nl = MUX_s_1_2_2((and_3172_nl), (and_3171_nl), or_11_cse);
  assign mux_1288_nl = MUX_s_1_2_2(and_tmp_188, mux_tmp_1209, or_11_cse);
  assign nor_1036_nl = ~((cfg_precision_1_sva_st_100[1]) | (~ or_tmp_3017));
  assign mux_2191_nl = MUX_s_1_2_2((nor_1036_nl), or_tmp_3017, cfg_precision_1_sva_st_100[0]);
  assign and_3167_nl = main_stage_v_9 & (~((mux_2191_nl) | (~ (chn_inp_in_crt_sva_9_739_736_1[1]))));
  assign nor_1037_nl = ~((cfg_precision_1_sva_st_101[1]) | (~ or_tmp_3020));
  assign mux_2196_nl = MUX_s_1_2_2((nor_1037_nl), or_tmp_3020, cfg_precision_1_sva_st_101[0]);
  assign and_3168_nl = main_stage_v_10 & (~((mux_2196_nl) | (~ (chn_inp_in_crt_sva_10_739_736_1[1]))));
  assign mux_1293_nl = MUX_s_1_2_2((and_3168_nl), (and_3167_nl), or_11_cse);
  assign nor_1034_nl = ~((cfg_precision_1_sva_st_100[1]) | (~ or_tmp_3025));
  assign mux_1294_nl = MUX_s_1_2_2((nor_1034_nl), or_tmp_3025, cfg_precision_1_sva_st_100[0]);
  assign and_3165_nl = main_stage_v_9 & (~ (mux_1294_nl)) & (chn_inp_in_crt_sva_9_739_736_1[1]);
  assign nor_1035_nl = ~((cfg_precision_1_sva_st_101[1]) | (~ or_tmp_3029));
  assign mux_1296_nl = MUX_s_1_2_2((nor_1035_nl), or_tmp_3029, cfg_precision_1_sva_st_101[0]);
  assign and_3166_nl = main_stage_v_10 & (~ (mux_1296_nl)) & (chn_inp_in_crt_sva_10_739_736_1[1]);
  assign mux_1298_nl = MUX_s_1_2_2((and_3166_nl), (and_3165_nl), or_11_cse);
  assign mux_1300_nl = MUX_s_1_2_2(and_tmp_187, mux_tmp_1221, or_11_cse);
  assign nor_1032_nl = ~((cfg_precision_1_sva_st_112[1]) | (~ or_tmp_3035));
  assign mux_2190_nl = MUX_s_1_2_2((nor_1032_nl), or_tmp_3035, cfg_precision_1_sva_st_112[0]);
  assign and_3161_nl = main_stage_v_9 & (~((mux_2190_nl) | (~ (chn_inp_in_crt_sva_9_739_736_1[2]))));
  assign nor_1033_nl = ~((cfg_precision_1_sva_st_113[1]) | (~ or_tmp_3038));
  assign mux_2195_nl = MUX_s_1_2_2((nor_1033_nl), or_tmp_3038, cfg_precision_1_sva_st_113[0]);
  assign and_3162_nl = main_stage_v_10 & (~((mux_2195_nl) | (~ (chn_inp_in_crt_sva_10_739_736_1[2]))));
  assign mux_1305_nl = MUX_s_1_2_2((and_3162_nl), (and_3161_nl), or_11_cse);
  assign nor_1030_nl = ~((cfg_precision_1_sva_st_112[1]) | (~ or_tmp_3043));
  assign mux_1306_nl = MUX_s_1_2_2((nor_1030_nl), or_tmp_3043, cfg_precision_1_sva_st_112[0]);
  assign and_3159_nl = main_stage_v_9 & (~ (mux_1306_nl)) & (chn_inp_in_crt_sva_9_739_736_1[2]);
  assign nor_1031_nl = ~((cfg_precision_1_sva_st_113[1]) | (~ or_tmp_3047));
  assign mux_1308_nl = MUX_s_1_2_2((nor_1031_nl), or_tmp_3047, cfg_precision_1_sva_st_113[0]);
  assign and_3160_nl = main_stage_v_10 & (~ (mux_1308_nl)) & (chn_inp_in_crt_sva_10_739_736_1[2]);
  assign mux_1310_nl = MUX_s_1_2_2((and_3160_nl), (and_3159_nl), or_11_cse);
  assign mux_1312_nl = MUX_s_1_2_2(and_tmp_184, mux_tmp_1233, or_11_cse);
  assign nor_1028_nl = ~((cfg_precision_1_sva_st_124[1]) | (~ or_tmp_3053));
  assign mux_2189_nl = MUX_s_1_2_2((nor_1028_nl), or_tmp_3053, cfg_precision_1_sva_st_124[0]);
  assign and_3155_nl = main_stage_v_9 & (~((mux_2189_nl) | (~ (chn_inp_in_crt_sva_9_739_736_1[3]))));
  assign nor_1029_nl = ~((cfg_precision_1_sva_st_125[1]) | (~ or_tmp_3056));
  assign mux_2194_nl = MUX_s_1_2_2((nor_1029_nl), or_tmp_3056, cfg_precision_1_sva_st_125[0]);
  assign and_3156_nl = main_stage_v_10 & (~((mux_2194_nl) | (~ (chn_inp_in_crt_sva_10_739_736_1[3]))));
  assign mux_1317_nl = MUX_s_1_2_2((and_3156_nl), (and_3155_nl), or_11_cse);
  assign nor_1026_nl = ~((cfg_precision_1_sva_st_124[1]) | (~ or_tmp_3061));
  assign mux_1318_nl = MUX_s_1_2_2((nor_1026_nl), or_tmp_3061, cfg_precision_1_sva_st_124[0]);
  assign and_3153_nl = main_stage_v_9 & (~ (mux_1318_nl)) & (chn_inp_in_crt_sva_9_739_736_1[3]);
  assign nor_1027_nl = ~((cfg_precision_1_sva_st_125[1]) | (~ or_tmp_3065));
  assign mux_1320_nl = MUX_s_1_2_2((nor_1027_nl), or_tmp_3065, cfg_precision_1_sva_st_125[0]);
  assign and_3154_nl = main_stage_v_10 & (~ (mux_1320_nl)) & (chn_inp_in_crt_sva_10_739_736_1[3]);
  assign mux_1322_nl = MUX_s_1_2_2((and_3154_nl), (and_3153_nl), or_11_cse);
  assign mux_1324_nl = MUX_s_1_2_2(and_tmp_182, mux_tmp_1245, or_11_cse);
  assign nor_1362_nl = ~((~((~ (inp_lookup_2_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21]))
      | inp_lookup_2_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1)) | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_14);
  assign nor_1364_nl = ~((FpMul_6U_10U_2_p_mant_p1_2_sva[21]) | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_14);
  assign mux_872_nl = MUX_s_1_2_2((nor_1364_nl), (nor_1362_nl), nor_268_cse);
  assign nand_93_nl = ~(nor_267_cse & (mux_872_nl));
  assign mux_873_nl = MUX_s_1_2_2((nand_93_nl), IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_14,
      IsNaN_6U_10U_7_land_2_lpi_1_dfm_5);
  assign mux_875_nl = MUX_s_1_2_2(nand_tmp_94, (mux_873_nl), or_11_cse);
  assign mux_878_nl = MUX_s_1_2_2(not_tmp_793, (mux_875_nl), nor_266_cse);
  assign nor_1365_nl = ~((cfg_precision_1_sva_st_90!=2'b10) | (chn_inp_in_crt_sva_1_739_395_1[342]));
  assign nor_1366_nl = ~((~ chn_inp_in_rsci_bawt) | (cfg_precision_rsci_d!=2'b10)
      | (chn_inp_in_rsci_d_mxwt[737]));
  assign mux_879_nl = MUX_s_1_2_2((nor_1366_nl), (nor_1365_nl), main_stage_v_1);
  assign nor_1367_nl = ~((~ main_stage_v_1) | (cfg_precision_1_sva_st_90!=2'b10)
      | (chn_inp_in_crt_sva_1_739_395_1[342]));
  assign mux_880_nl = MUX_s_1_2_2(not_tmp_793, nand_tmp_94, nor_1367_nl);
  assign mux_881_nl = MUX_s_1_2_2((mux_880_nl), (mux_879_nl), or_11_cse);
  assign mux_882_nl = MUX_s_1_2_2((mux_881_nl), (mux_878_nl), main_stage_v_2);
  assign nand_378_nl = ~((FpFractionToFloat_35U_6U_10U_1_mux_tmp[4:3]==2'b11) & (IntLeadZero_35U_1_leading_sign_35_0_rtn_1_sva_2[5])
      & inp_lookup_1_FpMantRNE_36U_11U_1_else_and_svs_2 & (~ IsNaN_6U_10U_6_nor_tmp)
      & FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_st_2 & (FpFractionToFloat_35U_6U_10U_1_mux_tmp[2:0]==3'b111)
      & (~ (chn_inp_in_crt_sva_1_739_395_1[341])));
  assign mux_1326_nl = MUX_s_1_2_2((nand_378_nl), (chn_inp_in_crt_sva_1_739_395_1[341]),
      and_3149_cse);
  assign nor_1021_nl = ~((~ main_stage_v_1) | (cfg_precision_1_sva_st_90[0]) | (~((cfg_precision_1_sva_st_90[1])
      & (mux_1326_nl))));
  assign nor_1022_nl = ~((~((~(IsNaN_6U_10U_7_land_1_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_14))
      | (chn_inp_in_crt_sva_2_739_736_1[0]))) | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10));
  assign mux_1327_nl = MUX_s_1_2_2((nor_1022_nl), (nor_1021_nl), or_11_cse);
  assign nand_376_nl = ~((FpFractionToFloat_35U_6U_10U_1_mux_40_tmp==5'b11111) &
      (IntLeadZero_35U_1_leading_sign_35_0_rtn_2_sva_2[5]) & inp_lookup_2_FpMantRNE_36U_11U_1_else_and_svs_2
      & (~ IsNaN_6U_10U_6_nor_1_tmp) & FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_st_2
      & (~ (chn_inp_in_crt_sva_1_739_395_1[342])));
  assign mux_1328_nl = MUX_s_1_2_2((nand_376_nl), (chn_inp_in_crt_sva_1_739_395_1[342]),
      and_4145_cse);
  assign nor_1018_nl = ~((~ main_stage_v_1) | (cfg_precision_1_sva_st_90[0]) | (~((cfg_precision_1_sva_st_90[1])
      & (mux_1328_nl))));
  assign nor_1019_nl = ~((~((~ or_tmp_3087) | (chn_inp_in_crt_sva_2_739_736_1[1])))
      | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10));
  assign mux_1329_nl = MUX_s_1_2_2((nor_1019_nl), (nor_1018_nl), or_11_cse);
  assign nor_1014_nl = ~(((FpFractionToFloat_35U_6U_10U_1_mux_41_tmp==5'b11111) &
      (IntLeadZero_35U_1_leading_sign_35_0_rtn_3_sva_2[5]) & inp_lookup_3_FpMantRNE_36U_11U_1_else_and_svs_2
      & (~ IsNaN_6U_10U_6_nor_2_tmp) & FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_st_2
      & (~ (chn_inp_in_crt_sva_1_739_395_1[343]))) | (~ main_stage_v_1) | (cfg_precision_1_sva_st_90!=2'b10));
  assign mux_1330_nl = MUX_s_1_2_2((nor_1014_nl), and_3389_cse, and_3249_cse);
  assign nor_1015_nl = ~((~(nor_1017_cse | (chn_inp_in_crt_sva_2_739_736_1[2])))
      | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10));
  assign mux_1331_nl = MUX_s_1_2_2((nor_1015_nl), (mux_1330_nl), or_11_cse);
  assign and_3371_nl = (chn_inp_in_crt_sva_1_739_395_1[344]) & main_stage_v_1 & (cfg_precision_1_sva_st_90==2'b10);
  assign nor_1010_nl = ~(((FpFractionToFloat_35U_6U_10U_1_mux_42_tmp==5'b11111) &
      (IntLeadZero_35U_1_leading_sign_35_0_rtn_sva_2[5]) & inp_lookup_4_FpMantRNE_36U_11U_1_else_and_svs_2
      & (~ IsNaN_6U_10U_6_nor_3_tmp) & FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2
      & (~ (chn_inp_in_crt_sva_1_739_395_1[344]))) | (~ main_stage_v_1) | (cfg_precision_1_sva_st_90!=2'b10));
  assign mux_1332_nl = MUX_s_1_2_2((nor_1010_nl), (and_3371_nl), and_3361_cse_1);
  assign nor_1011_nl = ~((~((~(IsNaN_6U_10U_7_land_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_lpi_1_dfm_st_14))
      | (chn_inp_in_crt_sva_2_739_736_1[3]))) | (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10));
  assign mux_1333_nl = MUX_s_1_2_2((nor_1011_nl), (mux_1332_nl), or_11_cse);
  assign nor_1801_nl = ~((cfg_precision_1_sva_st_80!=2'b10) | (chn_inp_in_crt_sva_3_739_736_1[0])
      | (~ main_stage_v_3));
  assign or_5835_nl = IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_14 | IsNaN_6U_10U_7_land_1_lpi_1_dfm_5;
  assign mux_2001_nl = MUX_s_1_2_2((or_5835_nl), (nor_1801_nl), or_5800_cse);
  assign or_3116_nl = (~ (inp_lookup_2_FpMul_6U_10U_2_p_mant_p1_mul_tmp[21])) | inp_lookup_2_FpMul_6U_10U_2_else_2_else_if_if_acc_1_itm_5_1
      | (chn_inp_in_crt_sva_2_739_736_1[1]) | (cfg_precision_1_sva_st_91!=2'b10);
  assign or_3118_nl = (~ (FpMul_6U_10U_2_p_mant_p1_2_sva[21])) | (chn_inp_in_crt_sva_2_739_736_1[1])
      | (cfg_precision_1_sva_st_91!=2'b10);
  assign mux_1334_nl = MUX_s_1_2_2((or_3118_nl), (or_3116_nl), nor_268_cse);
  assign mux_1335_nl = MUX_s_1_2_2(or_tmp_736, (mux_1334_nl), nor_267_cse);
  assign or_3121_nl = or_tmp_3087 | (mux_1335_nl);
  assign mux_1336_nl = MUX_s_1_2_2(or_tmp_736, or_tmp_3123, main_stage_v_3);
  assign mux_1337_nl = MUX_s_1_2_2((mux_1336_nl), (or_3121_nl), or_11_cse);
  assign mux_1339_nl = MUX_s_1_2_2(or_740_cse, or_tmp_3123, main_stage_v_3);
  assign or_3130_nl = (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[1]) |
      (cfg_precision_1_sva_st_80!=2'b10) | IsNaN_6U_10U_6_land_2_lpi_1_dfm_5 | IsNaN_6U_10U_7_land_2_lpi_1_dfm_6
      | nor_1371_cse;
  assign mux_1340_nl = MUX_s_1_2_2((or_3130_nl), (mux_1339_nl), main_stage_v_1);
  assign mux_1341_nl = MUX_s_1_2_2((mux_1340_nl), mux_400_cse, or_11_cse);
  assign mux_1342_nl = MUX_s_1_2_2((mux_1341_nl), (mux_1337_nl), main_stage_v_2);
  assign and_994_nl = or_tmp_440 & or_tmp_439;
  assign nor_682_nl = ~((chn_inp_in_crt_sva_2_739_736_1[2]) | (~ main_stage_v_2));
  assign mux_1883_nl = MUX_s_1_2_2(or_tmp_440, (and_994_nl), nor_682_nl);
  assign or_4372_nl = (~ main_stage_v_3) | (chn_inp_in_crt_sva_3_739_736_1[2]);
  assign mux_1884_nl = MUX_s_1_2_2((mux_1883_nl), or_dcpl_167, or_4372_nl);
  assign or_5142_nl = main_stage_v_3 | (chn_inp_in_crt_sva_2_739_736_1[2]) | (~ main_stage_v_2)
      | (cfg_precision_1_sva_st_91!=2'b10);
  assign mux_1952_nl = MUX_s_1_2_2((or_5142_nl), (mux_1884_nl), or_11_cse);
  assign or_5834_nl = IsNaN_6U_10U_2_land_lpi_1_dfm_st_14 | IsNaN_6U_10U_7_land_lpi_1_dfm_5;
  assign mux_2002_nl = MUX_s_1_2_2((or_5834_nl), nor_1800_cse, or_5809_cse);
  assign or_nl = (fsm_output[1]) | IsNaN_6U_10U_2_land_lpi_1_dfm_st_14 | IsNaN_6U_10U_7_land_lpi_1_dfm_5;
  assign mux_2003_nl = MUX_s_1_2_2((or_nl), nor_1800_cse, or_5809_cse);
  assign nor_1005_nl = ~((~ inp_lookup_4_FpMantRNE_49U_24U_1_else_and_tmp) | (cfg_precision_1_sva_st_82[0])
      | not_tmp_374);
  assign nor_1006_nl = ~((~ or_tmp_3132) | (cfg_precision_1_sva_st_82[0]) | not_tmp_374);
  assign mux_1343_nl = MUX_s_1_2_2((nor_1006_nl), (nor_1005_nl), chn_inp_in_crt_sva_5_739_736_1[3]);
  assign mux_1344_nl = MUX_s_1_2_2(or_tmp_2695, inp_lookup_4_FpMantRNE_49U_24U_1_else_and_svs_2,
      chn_inp_in_crt_sva_6_739_736_1[3]);
  assign nor_1007_nl = ~((~ main_stage_v_6) | (cfg_precision_1_sva_st_83[0]) | (~((cfg_precision_1_sva_st_83[1])
      & (mux_1344_nl))));
  assign mux_1345_nl = MUX_s_1_2_2((nor_1007_nl), (mux_1343_nl), or_11_cse);
  assign nor_1003_nl = ~((chn_inp_in_crt_sva_5_739_736_1[3]) | (~ or_tmp_3132) |
      (cfg_precision_1_sva_st_82[0]) | not_tmp_374);
  assign nor_1004_nl = ~((chn_inp_in_crt_sva_6_739_736_1[3]) | (cfg_precision_1_sva_st_83!=2'b10)
      | not_tmp_1108);
  assign mux_1346_nl = MUX_s_1_2_2((nor_1004_nl), (nor_1003_nl), or_11_cse);
  assign mux_1348_nl = MUX_s_1_2_2(or_tmp_3156, or_tmp_3152, inp_lookup_3_FpMantRNE_49U_24U_1_else_and_tmp);
  assign mux_1349_nl = MUX_s_1_2_2(or_tmp_3160, or_tmp_2768, reg_inp_lookup_3_FpMantRNE_49U_24U_1_else_and_svs_1_cse);
  assign mux_1350_nl = MUX_s_1_2_2((mux_1349_nl), (mux_1348_nl), or_11_cse);
  assign mux_1351_nl = MUX_s_1_2_2(or_tmp_3160, or_tmp_3156, or_11_cse);
  assign mux_1352_nl = MUX_s_1_2_2(or_tmp_2768, or_tmp_3152, or_11_cse);
  assign FpMul_6U_10U_1_o_mant_or_nl = and_dcpl_1624 | (and_1185_tmp & mux_1958_m1c);
  assign FpMul_6U_10U_1_o_mant_and_8_nl = (~ and_1185_tmp) & mux_1958_m1c;
  assign nor_1864_nl = ~((chn_inp_in_crt_sva_5_739_736_1[2]) | (~ or_tmp_3153));
  assign nor_1865_nl = ~((FpAdd_8U_23U_1_int_mant_p1_3_sva_3[49]) | (~ or_2676_cse));
  assign mux_2127_nl = MUX_s_1_2_2((nor_1865_nl), or_2676_cse, inp_lookup_3_FpAdd_8U_23U_1_if_3_if_acc_1_itm_7);
  assign or_6120_nl = IsNaN_8U_23U_3_land_3_lpi_1_dfm_6 | (mux_2127_nl);
  assign mux_2128_nl = MUX_s_1_2_2(or_tmp_3153, (or_6120_nl), chn_inp_in_crt_sva_5_739_736_1[2]);
  assign mux_2129_nl = MUX_s_1_2_2((mux_2128_nl), (nor_1864_nl), IsNaN_8U_23U_2_land_3_lpi_1_dfm_9);
  assign and_3370_nl = inp_lookup_2_FpMantRNE_49U_24U_1_else_and_tmp & (cfg_precision_1_sva_st_82==2'b10)
      & main_stage_v_5;
  assign and_3140_nl = or_tmp_3180 & (cfg_precision_1_sva_st_82==2'b10) & main_stage_v_5;
  assign mux_1357_nl = MUX_s_1_2_2((and_3140_nl), (and_3370_nl), chn_inp_in_crt_sva_5_739_736_1[1]);
  assign mux_1358_nl = MUX_s_1_2_2(or_tmp_2738, inp_lookup_2_FpMantRNE_49U_24U_1_else_and_svs_2,
      chn_inp_in_crt_sva_6_739_736_1[1]);
  assign nor_996_nl = ~((~ main_stage_v_6) | (cfg_precision_1_sva_st_83[0]) | (~((cfg_precision_1_sva_st_83[1])
      & (mux_1358_nl))));
  assign mux_1359_nl = MUX_s_1_2_2((nor_996_nl), (mux_1357_nl), or_11_cse);
  assign nor_992_nl = ~((chn_inp_in_crt_sva_5_739_736_1[1]) | (~(or_tmp_3180 & (cfg_precision_1_sva_st_82==2'b10)
      & main_stage_v_5)));
  assign nor_993_nl = ~((chn_inp_in_crt_sva_6_739_736_1[1]) | (~ main_stage_v_6));
  assign nor_994_nl = ~((chn_inp_in_crt_sva_6_739_736_1[1]) | (~(IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_18
      & main_stage_v_6)));
  assign mux_1360_nl = MUX_s_1_2_2((nor_994_nl), (nor_993_nl), IsNaN_6U_10U_9_land_2_lpi_1_dfm_7);
  assign and_3139_nl = (~((cfg_precision_1_sva_st_83!=2'b10))) & (mux_1360_nl);
  assign mux_1361_nl = MUX_s_1_2_2((and_3139_nl), (nor_992_nl), or_11_cse);
  assign nor_988_nl = ~((~ inp_lookup_1_FpMantRNE_49U_24U_1_else_and_tmp) | (cfg_precision_1_sva_st_82[0])
      | not_tmp_374);
  assign nor_989_nl = ~((~ or_tmp_3200) | (cfg_precision_1_sva_st_82[0]) | not_tmp_374);
  assign mux_1363_nl = MUX_s_1_2_2((nor_989_nl), (nor_988_nl), chn_inp_in_crt_sva_5_739_736_1[0]);
  assign mux_1364_nl = MUX_s_1_2_2(or_tmp_2723, inp_lookup_1_FpMantRNE_49U_24U_1_else_and_svs_2,
      chn_inp_in_crt_sva_6_739_736_1[0]);
  assign nor_990_nl = ~((~ main_stage_v_6) | (cfg_precision_1_sva_st_83[0]) | (~((cfg_precision_1_sva_st_83[1])
      & (mux_1364_nl))));
  assign mux_1365_nl = MUX_s_1_2_2((nor_990_nl), (mux_1363_nl), or_11_cse);
  assign nor_986_nl = ~((chn_inp_in_crt_sva_5_739_736_1[0]) | (~ or_tmp_3200) | (cfg_precision_1_sva_st_82[0])
      | not_tmp_374);
  assign nor_987_nl = ~((cfg_precision_1_sva_st_83!=2'b10) | (chn_inp_in_crt_sva_6_739_736_1[0])
      | (~(or_tmp_2723 & main_stage_v_6)));
  assign mux_1366_nl = MUX_s_1_2_2((nor_987_nl), (nor_986_nl), or_11_cse);
  assign mux_1368_nl = MUX_s_1_2_2(nand_tmp_162, or_tmp_1255, or_11_cse);
  assign mux_1369_nl = MUX_s_1_2_2(nand_tmp_163, or_tmp_1302, or_11_cse);
  assign mux_1370_nl = MUX_s_1_2_2(nand_tmp_164, or_tmp_1312, or_11_cse);
  assign mux_1371_nl = MUX_s_1_2_2(nand_tmp_165, or_tmp_1340, or_11_cse);
  assign or_3241_nl = IsNaN_6U_10U_2_land_lpi_1_dfm_23 | (cfg_precision_1_sva_19!=2'b10)
      | (~((cfg_precision_1_sva_st_124!=2'b10) | (~ FpAdd_6U_10U_is_a_greater_acc_3_itm_6_1)
      | IsNaN_6U_10U_3_IsNaN_6U_10U_3_nor_3_tmp));
  assign mux_1379_nl = MUX_s_1_2_2(inp_lookup_else_unequal_tmp_35, (or_3241_nl),
      chn_inp_in_crt_sva_9_739_736_1[3]);
  assign and_3137_nl = main_stage_v_9 & (~ (mux_1379_nl));
  assign or_3246_nl = IsNaN_6U_10U_2_land_lpi_1_dfm_24 | (cfg_precision_1_sva_20!=2'b10)
      | (~(IsNaN_6U_10U_3_land_lpi_1_dfm_6 | (~ reg_inp_lookup_4_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse)));
  assign mux_1383_nl = MUX_s_1_2_2(inp_lookup_else_unequal_tmp_36, (or_3246_nl),
      chn_inp_in_crt_sva_10_739_736_1[3]);
  assign and_3138_nl = main_stage_v_10 & (~ (mux_1383_nl));
  assign mux_1384_nl = MUX_s_1_2_2((and_3138_nl), (and_3137_nl), or_11_cse);
  assign or_3252_nl = IsNaN_6U_10U_2_land_3_lpi_1_dfm_23 | (cfg_precision_1_sva_19!=2'b10)
      | (~((cfg_precision_1_sva_st_112!=2'b10) | (~ FpAdd_6U_10U_is_a_greater_acc_2_itm_6_1)
      | IsNaN_6U_10U_3_IsNaN_6U_10U_3_nor_2_tmp));
  assign mux_1388_nl = MUX_s_1_2_2(inp_lookup_else_unequal_tmp_35, (or_3252_nl),
      chn_inp_in_crt_sva_9_739_736_1[2]);
  assign and_3135_nl = main_stage_v_9 & (~ (mux_1388_nl));
  assign or_3257_nl = IsNaN_6U_10U_2_land_3_lpi_1_dfm_24 | (cfg_precision_1_sva_20!=2'b10)
      | (~(IsNaN_6U_10U_3_land_3_lpi_1_dfm_6 | (~ reg_inp_lookup_3_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse)));
  assign mux_1392_nl = MUX_s_1_2_2(inp_lookup_else_unequal_tmp_36, (or_3257_nl),
      chn_inp_in_crt_sva_10_739_736_1[2]);
  assign and_3136_nl = main_stage_v_10 & (~ (mux_1392_nl));
  assign mux_1393_nl = MUX_s_1_2_2((and_3136_nl), (and_3135_nl), or_11_cse);
  assign or_3263_nl = IsNaN_6U_10U_2_land_2_lpi_1_dfm_23 | (cfg_precision_1_sva_19!=2'b10)
      | (~((cfg_precision_1_sva_st_100!=2'b10) | (~ FpAdd_6U_10U_is_a_greater_acc_1_itm_6_1)
      | IsNaN_6U_10U_3_IsNaN_6U_10U_3_nor_1_tmp));
  assign mux_1397_nl = MUX_s_1_2_2(inp_lookup_else_unequal_tmp_35, (or_3263_nl),
      chn_inp_in_crt_sva_9_739_736_1[1]);
  assign and_3133_nl = main_stage_v_9 & (~ (mux_1397_nl));
  assign or_3268_nl = IsNaN_6U_10U_2_land_2_lpi_1_dfm_24 | (cfg_precision_1_sva_20!=2'b10)
      | (~(IsNaN_6U_10U_3_land_2_lpi_1_dfm_6 | (~ reg_inp_lookup_2_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse)));
  assign mux_1401_nl = MUX_s_1_2_2(inp_lookup_else_unequal_tmp_36, (or_3268_nl),
      chn_inp_in_crt_sva_10_739_736_1[1]);
  assign and_3134_nl = main_stage_v_10 & (~ (mux_1401_nl));
  assign mux_1402_nl = MUX_s_1_2_2((and_3134_nl), (and_3133_nl), or_11_cse);
  assign or_3274_nl = IsNaN_6U_10U_2_land_1_lpi_1_dfm_23 | (cfg_precision_1_sva_19!=2'b10)
      | (~((cfg_precision_1_sva_st_86!=2'b10) | (~ FpAdd_6U_10U_is_a_greater_acc_itm_6_1)
      | IsNaN_6U_10U_3_IsNaN_6U_10U_3_nor_tmp));
  assign mux_1406_nl = MUX_s_1_2_2(inp_lookup_else_unequal_tmp_35, (or_3274_nl),
      chn_inp_in_crt_sva_9_739_736_1[0]);
  assign and_3131_nl = main_stage_v_9 & (~ (mux_1406_nl));
  assign or_3279_nl = IsNaN_6U_10U_2_land_1_lpi_1_dfm_24 | (cfg_precision_1_sva_20!=2'b10)
      | (~(IsNaN_6U_10U_3_land_1_lpi_1_dfm_6 | (~ reg_inp_lookup_1_FpAdd_6U_10U_is_a_greater_slc_6_svs_1_cse)));
  assign mux_1410_nl = MUX_s_1_2_2(inp_lookup_else_unequal_tmp_36, (or_3279_nl),
      chn_inp_in_crt_sva_10_739_736_1[0]);
  assign and_3132_nl = main_stage_v_10 & (~ (mux_1410_nl));
  assign mux_1411_nl = MUX_s_1_2_2((and_3132_nl), (and_3131_nl), or_11_cse);
  assign or_3282_nl = (cfg_precision_1_sva_19!=2'b10) | not_tmp_1369;
  assign mux_1412_nl = MUX_s_1_2_2(not_tmp_1369, (or_3282_nl), chn_inp_in_crt_sva_9_739_736_1[0]);
  assign nor_975_nl = ~((cfg_precision_1_sva_19!=2'b10) | not_tmp_1369);
  assign nor_976_nl = ~(IsNaN_6U_10U_3_IsNaN_6U_10U_3_nor_tmp | (cfg_precision_1_sva_19!=2'b10)
      | not_tmp_1369);
  assign mux_1413_nl = MUX_s_1_2_2((nor_976_nl), (nor_975_nl), IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_21);
  assign nand_198_nl = ~((~((~ (chn_inp_in_crt_sva_9_739_736_1[0])) | (cfg_precision_1_sva_st_86!=2'b10)))
      & (mux_1413_nl));
  assign mux_1414_nl = MUX_s_1_2_2((nand_198_nl), (mux_1412_nl), IsNaN_6U_10U_2_land_1_lpi_1_dfm_23);
  assign or_3292_nl = IsNaN_6U_10U_3_land_1_lpi_1_dfm_6 | or_3291_cse;
  assign mux_1418_nl = MUX_s_1_2_2((or_3292_nl), or_3291_cse, IsNaN_6U_10U_2_land_1_lpi_1_dfm_24);
  assign nand_199_nl = ~(main_stage_v_10 & (chn_inp_in_crt_sva_10_739_736_1[0]) &
      (~ (mux_1418_nl)));
  assign mux_1419_nl = MUX_s_1_2_2((nand_199_nl), (mux_1414_nl), or_11_cse);
  assign and_3129_nl = ((chn_inp_in_crt_sva_10_739_736_1!=4'b0000)) & main_stage_v_10;
  assign mux_1420_nl = MUX_s_1_2_2((and_3129_nl), nor_tmp_464, or_11_cse);
  assign or_3298_nl = (cfg_precision_1_sva_19!=2'b10) | not_tmp_1373;
  assign mux_1421_nl = MUX_s_1_2_2(not_tmp_1373, (or_3298_nl), chn_inp_in_crt_sva_9_739_736_1[1]);
  assign nor_973_nl = ~((cfg_precision_1_sva_19!=2'b10) | not_tmp_1373);
  assign nor_974_nl = ~(IsNaN_6U_10U_3_IsNaN_6U_10U_3_nor_1_tmp | (cfg_precision_1_sva_19!=2'b10)
      | not_tmp_1373);
  assign mux_1422_nl = MUX_s_1_2_2((nor_974_nl), (nor_973_nl), IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_21);
  assign nand_200_nl = ~((~((~ (chn_inp_in_crt_sva_9_739_736_1[1])) | (cfg_precision_1_sva_st_100!=2'b10)))
      & (mux_1422_nl));
  assign mux_1423_nl = MUX_s_1_2_2((nand_200_nl), (mux_1421_nl), IsNaN_6U_10U_2_land_2_lpi_1_dfm_23);
  assign or_3308_nl = IsNaN_6U_10U_3_land_2_lpi_1_dfm_6 | or_3291_cse;
  assign mux_1427_nl = MUX_s_1_2_2((or_3308_nl), or_3291_cse, IsNaN_6U_10U_2_land_2_lpi_1_dfm_24);
  assign nand_201_nl = ~(main_stage_v_10 & (chn_inp_in_crt_sva_10_739_736_1[1]) &
      (~ (mux_1427_nl)));
  assign mux_1428_nl = MUX_s_1_2_2((nand_201_nl), (mux_1423_nl), or_11_cse);
  assign or_3311_nl = (cfg_precision_1_sva_19!=2'b10) | not_tmp_1377;
  assign mux_1429_nl = MUX_s_1_2_2(not_tmp_1377, (or_3311_nl), chn_inp_in_crt_sva_9_739_736_1[2]);
  assign nor_971_nl = ~((cfg_precision_1_sva_19!=2'b10) | not_tmp_1377);
  assign nor_972_nl = ~(IsNaN_6U_10U_3_IsNaN_6U_10U_3_nor_2_tmp | (cfg_precision_1_sva_19!=2'b10)
      | not_tmp_1377);
  assign mux_1430_nl = MUX_s_1_2_2((nor_972_nl), (nor_971_nl), IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_21);
  assign nand_202_nl = ~((~((~ (chn_inp_in_crt_sva_9_739_736_1[2])) | (cfg_precision_1_sva_st_112!=2'b10)))
      & (mux_1430_nl));
  assign mux_1431_nl = MUX_s_1_2_2((nand_202_nl), (mux_1429_nl), IsNaN_6U_10U_2_land_3_lpi_1_dfm_23);
  assign or_3321_nl = IsNaN_6U_10U_3_land_3_lpi_1_dfm_6 | or_3291_cse;
  assign mux_1435_nl = MUX_s_1_2_2((or_3321_nl), or_3291_cse, IsNaN_6U_10U_2_land_3_lpi_1_dfm_24);
  assign nand_203_nl = ~(main_stage_v_10 & (chn_inp_in_crt_sva_10_739_736_1[2]) &
      (~ (mux_1435_nl)));
  assign mux_1436_nl = MUX_s_1_2_2((nand_203_nl), (mux_1431_nl), or_11_cse);
  assign or_3324_nl = (cfg_precision_1_sva_19!=2'b10) | not_tmp_1381;
  assign mux_1437_nl = MUX_s_1_2_2(not_tmp_1381, (or_3324_nl), chn_inp_in_crt_sva_9_739_736_1[3]);
  assign nor_969_nl = ~((cfg_precision_1_sva_19!=2'b10) | not_tmp_1381);
  assign nor_970_nl = ~(IsNaN_6U_10U_3_IsNaN_6U_10U_3_nor_3_tmp | (cfg_precision_1_sva_19!=2'b10)
      | not_tmp_1381);
  assign mux_1438_nl = MUX_s_1_2_2((nor_970_nl), (nor_969_nl), IsNaN_6U_10U_2_land_lpi_1_dfm_st_20);
  assign nand_204_nl = ~((~((~ (chn_inp_in_crt_sva_9_739_736_1[3])) | (cfg_precision_1_sva_st_124!=2'b10)))
      & (mux_1438_nl));
  assign mux_1439_nl = MUX_s_1_2_2((nand_204_nl), (mux_1437_nl), IsNaN_6U_10U_2_land_lpi_1_dfm_23);
  assign or_3334_nl = IsNaN_6U_10U_3_land_lpi_1_dfm_6 | or_3291_cse;
  assign mux_1443_nl = MUX_s_1_2_2((or_3334_nl), or_3291_cse, IsNaN_6U_10U_2_land_lpi_1_dfm_24);
  assign nand_205_nl = ~(main_stage_v_10 & (chn_inp_in_crt_sva_10_739_736_1[3]) &
      (~ (mux_1443_nl)));
  assign mux_1444_nl = MUX_s_1_2_2((nand_205_nl), (mux_1439_nl), or_11_cse);
  assign nand_206_nl = ~(main_stage_v_2 & (chn_inp_in_crt_sva_2_739_736_1[0]) & (~
      mux_tmp_1367));
  assign mux_1446_nl = MUX_s_1_2_2((nand_206_nl), nand_694_cse, or_11_cse);
  assign or_3342_nl = nand_358_cse | not_tmp_1388;
  assign mux_1448_nl = MUX_s_1_2_2((or_3342_nl), or_tmp_213, or_11_cse);
  assign or_3345_nl = (~ (chn_inp_in_crt_sva_2_739_736_1[2])) | (~ main_stage_v_2)
      | (cfg_precision_1_sva_st_91[0]) | not_tmp_1391;
  assign mux_1450_nl = MUX_s_1_2_2((or_3345_nl), nand_693_cse, or_11_cse);
  assign mux_1451_nl = MUX_s_1_2_2((~ FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_7_0_1),
      FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_7_0_1, FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_7_1_1);
  assign or_3348_nl = (~ main_stage_v_2) | (~ (chn_inp_in_crt_sva_2_739_736_1[3]))
      | (cfg_precision_1_sva_st_91[0]) | (~((cfg_precision_1_sva_st_91[1]) & (mux_1451_nl)));
  assign mux_1452_nl = MUX_s_1_2_2((or_3348_nl), or_tmp_347, or_11_cse);
  assign mux_1453_nl = MUX_s_1_2_2(or_tmp_439, mux_tmp_1367, chn_inp_in_crt_sva_2_739_736_1[0]);
  assign and_3127_nl = main_stage_v_2 & (~ (mux_1453_nl));
  assign or_3350_nl = (cfg_precision_1_sva_st_80[0]) | not_tmp_940;
  assign mux_1454_nl = MUX_s_1_2_2(or_tmp_440, (or_3350_nl), chn_inp_in_crt_sva_3_739_736_1[0]);
  assign and_3128_nl = main_stage_v_3 & (~ (mux_1454_nl));
  assign mux_1455_nl = MUX_s_1_2_2((and_3128_nl), (and_3127_nl), or_11_cse);
  assign or_3353_nl = (cfg_precision_1_sva_st_91!=2'b10) | not_tmp_1388;
  assign mux_1456_nl = MUX_s_1_2_2(or_tmp_439, (or_3353_nl), chn_inp_in_crt_sva_2_739_736_1[1]);
  assign and_3125_nl = main_stage_v_2 & (~ (mux_1456_nl));
  assign mux_1457_nl = MUX_s_1_2_2(or_tmp_440, mux_tmp_950, chn_inp_in_crt_sva_3_739_736_1[1]);
  assign and_3126_nl = main_stage_v_3 & (~ (mux_1457_nl));
  assign mux_1458_nl = MUX_s_1_2_2((and_3126_nl), (and_3125_nl), or_11_cse);
  assign or_3356_nl = (~ main_stage_v_2) | (cfg_precision_1_sva_st_91[0]) | not_tmp_1391;
  assign mux_1459_nl = MUX_s_1_2_2(or_2176_cse, (or_3356_nl), chn_inp_in_crt_sva_2_739_736_1[2]);
  assign mux_1460_nl = MUX_s_1_2_2(or_tmp_440, mux_tmp_966, chn_inp_in_crt_sva_3_739_736_1[2]);
  assign nand_211_nl = ~(main_stage_v_3 & (~ (mux_1460_nl)));
  assign mux_1461_nl = MUX_s_1_2_2((nand_211_nl), (mux_1459_nl), or_11_cse);
  assign mux_1462_nl = MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_7_0_1,
      (~ FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_7_0_1), FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_lpi_1_dfm_7_1_1);
  assign nor_967_nl = ~((~ main_stage_v_2) | (cfg_precision_1_sva_st_91[0]) | (~((cfg_precision_1_sva_st_91[1])
      & (~((chn_inp_in_crt_sva_2_739_736_1[3]) & (mux_1462_nl))))));
  assign nor_968_nl = ~((~ main_stage_v_3) | (cfg_precision_1_sva_st_80[0]) | (~((cfg_precision_1_sva_st_80[1])
      & (~((chn_inp_in_crt_sva_3_739_736_1[3]) & mux_1061_cse)))));
  assign mux_1464_nl = MUX_s_1_2_2((nor_968_nl), (nor_967_nl), or_11_cse);
  assign inp_lookup_1_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_nl = (FpMul_6U_10U_2_o_mant_1_lpi_1_dfm_3_mx0w0!=10'b0000000000)
      | FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_3_5_mx1w1 | FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_3_4_mx0w0
      | (FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_3_3_0_mx0w0!=4'b0000);
  assign mux_1465_nl = MUX_s_1_2_2((~ inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4),
      inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4,
      inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4);
  assign or_3363_nl = (cfg_precision_1_sva_st_80[0]) | (~((cfg_precision_1_sva_st_80[1])
      & (mux_1465_nl)));
  assign mux_1466_nl = MUX_s_1_2_2((or_3363_nl), or_tmp_440, chn_inp_in_crt_sva_3_739_736_1[0]);
  assign nand_214_nl = ~(main_stage_v_3 & (~ (mux_1466_nl)));
  assign mux_1467_nl = MUX_s_1_2_2(nand_tmp_138, (nand_214_nl), or_11_cse);
  assign inp_lookup_2_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_nl = (FpMul_6U_10U_2_o_mant_2_lpi_1_dfm_3_mx0w0!=10'b0000000000)
      | FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_3_5_mx1w1 | FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_3_4_mx0w0
      | (FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_3_3_0_mx0w0!=4'b0000);
  assign mux_1468_nl = MUX_s_1_2_2(inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4,
      (~ inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4),
      inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4);
  assign or_3366_nl = (cfg_precision_1_sva_st_80!=2'b10) | (mux_1468_nl);
  assign mux_1469_nl = MUX_s_1_2_2((or_3366_nl), or_tmp_440, chn_inp_in_crt_sva_3_739_736_1[1]);
  assign nand_215_nl = ~(main_stage_v_3 & (~ (mux_1469_nl)));
  assign mux_1470_nl = MUX_s_1_2_2(nand_tmp_142, (nand_215_nl), or_11_cse);
  assign inp_lookup_3_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_nl = (FpMul_6U_10U_2_o_mant_3_lpi_1_dfm_3_mx1w1!=10'b0000000000)
      | FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_3_5_mx1w1 | FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_3_4_mx0w0
      | (FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_3_3_0_mx0w0!=4'b0000);
  assign mux_1471_nl = MUX_s_1_2_2(inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4,
      (~ inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4),
      inp_lookup_3_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4);
  assign or_3369_nl = (cfg_precision_1_sva_st_80!=2'b10) | (mux_1471_nl);
  assign mux_1472_nl = MUX_s_1_2_2((or_3369_nl), or_tmp_440, chn_inp_in_crt_sva_3_739_736_1[2]);
  assign nand_216_nl = ~(main_stage_v_3 & (~ (mux_1472_nl)));
  assign mux_1473_nl = MUX_s_1_2_2(nand_tmp_146, (nand_216_nl), or_11_cse);
  assign inp_lookup_4_FpAdd_6U_10U_1_IsZero_6U_10U_9_or_nl = (FpMul_6U_10U_2_o_mant_lpi_1_dfm_3_mx0w0!=10'b0000000000)
      | FpMul_6U_10U_2_o_expo_lpi_1_dfm_3_5_mx0w0 | FpMul_6U_10U_2_o_expo_lpi_1_dfm_3_4_mx0w0
      | (FpMul_6U_10U_2_o_expo_lpi_1_dfm_3_3_0_mx0w0!=4'b0000);
  assign nor_963_nl = ~((~(inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4
      | (chn_inp_in_crt_sva_3_739_736_1[3]))) | (cfg_precision_1_sva_st_80!=2'b10));
  assign nor_965_nl = ~((~((~ inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_4)
      | (chn_inp_in_crt_sva_3_739_736_1[3]))) | (cfg_precision_1_sva_st_80!=2'b10));
  assign mux_1474_nl = MUX_s_1_2_2((nor_965_nl), (nor_963_nl), inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_4);
  assign nand_217_nl = ~(main_stage_v_3 & (mux_1474_nl));
  assign mux_1475_nl = MUX_s_1_2_2(nand_tmp_148, (nand_217_nl), or_11_cse);
  assign mux_1478_nl = MUX_s_1_2_2(mux_1476_cse, nor_959_cse, chn_inp_in_crt_sva_4_739_736_1[3]);
  assign mux_1481_nl = MUX_s_1_2_2(mux_1480_cse, nor_1113_cse, chn_inp_in_crt_sva_5_739_736_1[3]);
  assign mux_1482_nl = MUX_s_1_2_2((mux_1481_nl), (mux_1478_nl), or_11_cse);
  assign mux_1484_nl = MUX_s_1_2_2(mux_1483_cse, nor_959_cse, chn_inp_in_crt_sva_4_739_736_1[3]);
  assign mux_1487_nl = MUX_s_1_2_2(mux_1480_cse, nor_1113_cse, or_5152_cse);
  assign mux_1488_nl = MUX_s_1_2_2((mux_1487_nl), (mux_1484_nl), or_11_cse);
  assign mux_1491_nl = MUX_s_1_2_2(mux_1476_cse, nor_950_cse, chn_inp_in_crt_sva_4_739_736_1[2]);
  assign mux_1494_nl = MUX_s_1_2_2(mux_1493_cse, nor_952_cse, chn_inp_in_crt_sva_5_739_736_1[2]);
  assign mux_1495_nl = MUX_s_1_2_2((mux_1494_nl), (mux_1491_nl), or_11_cse);
  assign mux_1497_nl = MUX_s_1_2_2(mux_1483_cse, nor_950_cse, chn_inp_in_crt_sva_4_739_736_1[2]);
  assign or_3417_nl = IsNaN_6U_10U_8_land_3_lpi_1_dfm_4 | (chn_inp_in_crt_sva_5_739_736_1[2]);
  assign mux_1500_nl = MUX_s_1_2_2(mux_1493_cse, nor_952_cse, or_3417_nl);
  assign mux_1501_nl = MUX_s_1_2_2((mux_1500_nl), (mux_1497_nl), or_11_cse);
  assign mux_1504_nl = MUX_s_1_2_2(mux_1476_cse, nor_941_cse, chn_inp_in_crt_sva_4_739_736_1[1]);
  assign mux_1507_nl = MUX_s_1_2_2(mux_1506_cse, nor_943_cse, chn_inp_in_crt_sva_5_739_736_1[1]);
  assign mux_1508_nl = MUX_s_1_2_2((mux_1507_nl), (mux_1504_nl), or_11_cse);
  assign mux_1510_nl = MUX_s_1_2_2(mux_1483_cse, nor_941_cse, chn_inp_in_crt_sva_4_739_736_1[1]);
  assign mux_1513_nl = MUX_s_1_2_2(mux_1506_cse, nor_943_cse, or_5154_cse);
  assign mux_1514_nl = MUX_s_1_2_2((mux_1513_nl), (mux_1510_nl), or_11_cse);
  assign mux_1517_nl = MUX_s_1_2_2(mux_1476_cse, nor_932_cse, chn_inp_in_crt_sva_4_739_736_1[0]);
  assign mux_1520_nl = MUX_s_1_2_2(mux_1519_cse, nor_1124_cse, chn_inp_in_crt_sva_5_739_736_1[0]);
  assign mux_1521_nl = MUX_s_1_2_2((mux_1520_nl), (mux_1517_nl), or_11_cse);
  assign mux_1523_nl = MUX_s_1_2_2(mux_1483_cse, nor_932_cse, chn_inp_in_crt_sva_4_739_736_1[0]);
  assign mux_1526_nl = MUX_s_1_2_2(mux_1519_cse, nor_1124_cse, or_5155_cse);
  assign mux_1527_nl = MUX_s_1_2_2((mux_1526_nl), (mux_1523_nl), or_11_cse);
  assign mux_1529_nl = MUX_s_1_2_2(and_3286_cse, mux_tmp_1450, or_11_cse);
  assign mux_1531_nl = MUX_s_1_2_2(and_3285_cse, mux_tmp_1452, or_11_cse);
  assign mux_1534_nl = MUX_s_1_2_2(and_3283_cse, main_stage_v_8, chn_inp_in_crt_sva_8_739_736_1[2]);
  assign mux_1535_nl = MUX_s_1_2_2((mux_1534_nl), mux_tmp_1454, or_11_cse);
  assign mux_1538_nl = MUX_s_1_2_2(and_3281_cse, main_stage_v_8, chn_inp_in_crt_sva_8_739_736_1[3]);
  assign mux_1539_nl = MUX_s_1_2_2((mux_1538_nl), mux_tmp_1458, or_11_cse);
  assign and_3550_nl = (~ IsInf_6U_23U_1_land_lpi_1_dfm_mx0w0) & or_11_cse;
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_mux_44_nl = MUX_v_4_2_2(FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_3_0_1,
      4'b1110, IsInf_6U_23U_1_land_lpi_1_dfm_mx0w0);
  assign nl_inp_lookup_4_FpExpoWidthInc_6U_8U_23U_0U_1U_1_else_acc_nl = conv_u2u_2_3({1'b1
      , FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_5_1}) + 3'b1;
  assign inp_lookup_4_FpExpoWidthInc_6U_8U_23U_0U_1U_1_else_acc_nl = nl_inp_lookup_4_FpExpoWidthInc_6U_8U_23U_0U_1U_1_else_acc_nl[2:0];
  assign IsZero_6U_23U_1_aelse_IsZero_6U_23U_1_or_3_nl = (FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_22_13_lpi_1_dfm_mx0w1!=10'b0000000000)
      | (FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_9_0_lpi_1_dfm!=10'b0000000000)
      | FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_5_1 | FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_4_1
      | (FpAdd_6U_10U_1_o_expo_lpi_1_dfm_10_3_0_1!=4'b0000);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_15_nl
      = MUX_v_3_2_2(3'b000, (inp_lookup_4_FpExpoWidthInc_6U_8U_23U_0U_1U_1_else_acc_nl),
      (IsZero_6U_23U_1_aelse_IsZero_6U_23U_1_or_3_nl));
  assign or_5264_nl = (cfg_precision_1_sva_st_85!=2'b10) | (chn_inp_in_crt_sva_8_739_736_1[3]);
  assign IsInf_6U_23U_1_aelse_mux_7_nl = MUX_s_1_2_2(IsInf_6U_23U_1_land_lpi_1_dfm_mx0w0,
      IsInf_6U_23U_1_land_lpi_1_dfm, or_5264_nl);
  assign and_4212_nl = mux_1541_cse & (chn_inp_in_crt_sva_8_739_736_1[3]);
  assign nor_1758_nl = ~((cfg_precision_1_sva_st_124[0]) | (~((cfg_precision_1_sva_st_124[1])
      & main_stage_v_9)));
  assign mux_2198_nl = MUX_s_1_2_2(main_stage_v_9, (nor_1758_nl), or_3489_cse);
  assign and_4214_nl = (mux_2198_nl) & (chn_inp_in_crt_sva_9_739_736_1[3]);
  assign mux_1547_nl = MUX_s_1_2_2((and_4214_nl), (and_4212_nl), or_11_cse);
  assign and_3552_nl = (~ IsInf_6U_23U_1_land_3_lpi_1_dfm_mx0w0) & or_11_cse;
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_mux_31_nl = MUX_v_4_2_2(FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_3_0_1,
      4'b1110, IsInf_6U_23U_1_land_3_lpi_1_dfm_mx0w0);
  assign nl_inp_lookup_3_FpExpoWidthInc_6U_8U_23U_0U_1U_1_else_acc_nl = conv_u2u_2_3({1'b1
      , FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_5_1}) + 3'b1;
  assign inp_lookup_3_FpExpoWidthInc_6U_8U_23U_0U_1U_1_else_acc_nl = nl_inp_lookup_3_FpExpoWidthInc_6U_8U_23U_0U_1U_1_else_acc_nl[2:0];
  assign IsZero_6U_23U_1_aelse_IsZero_6U_23U_1_or_2_nl = (FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_22_13_3_lpi_1_dfm_mx0w1!=10'b0000000000)
      | (FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_9_0_3_lpi_1_dfm!=10'b0000000000)
      | FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_5_1 | FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_4_1
      | (FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_10_3_0_1!=4'b0000);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_10_nl
      = MUX_v_3_2_2(3'b000, (inp_lookup_3_FpExpoWidthInc_6U_8U_23U_0U_1U_1_else_acc_nl),
      (IsZero_6U_23U_1_aelse_IsZero_6U_23U_1_or_2_nl));
  assign or_5260_nl = (cfg_precision_1_sva_st_85!=2'b10) | (chn_inp_in_crt_sva_8_739_736_1[2]);
  assign IsInf_6U_23U_1_aelse_mux_5_nl = MUX_s_1_2_2(IsInf_6U_23U_1_land_3_lpi_1_dfm_mx0w0,
      IsInf_6U_23U_1_land_3_lpi_1_dfm, or_5260_nl);
  assign and_4213_nl = mux_1541_cse & (chn_inp_in_crt_sva_8_739_736_1[2]);
  assign nor_1754_nl = ~((cfg_precision_1_sva_st_112[0]) | (~((cfg_precision_1_sva_st_112[1])
      & main_stage_v_9)));
  assign mux_2199_nl = MUX_s_1_2_2(main_stage_v_9, (nor_1754_nl), or_3489_cse);
  assign and_4215_nl = (mux_2199_nl) & (chn_inp_in_crt_sva_9_739_736_1[2]);
  assign mux_1555_nl = MUX_s_1_2_2((and_4215_nl), (and_4213_nl), or_11_cse);
  assign and_3554_nl = (~ IsInf_6U_23U_1_land_2_lpi_1_dfm_mx0w0) & or_11_cse;
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_mux_18_nl = MUX_v_4_2_2(FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_3_0_1,
      4'b1110, IsInf_6U_23U_1_land_2_lpi_1_dfm_mx0w0);
  assign nl_inp_lookup_2_FpExpoWidthInc_6U_8U_23U_0U_1U_1_else_acc_nl = conv_u2u_2_3({1'b1
      , FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_5_1}) + 3'b1;
  assign inp_lookup_2_FpExpoWidthInc_6U_8U_23U_0U_1U_1_else_acc_nl = nl_inp_lookup_2_FpExpoWidthInc_6U_8U_23U_0U_1U_1_else_acc_nl[2:0];
  assign IsZero_6U_23U_1_aelse_IsZero_6U_23U_1_or_1_nl = (FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_22_13_2_lpi_1_dfm_mx0w1!=10'b0000000000)
      | (FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_9_0_2_lpi_1_dfm!=10'b0000000000)
      | FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_5_1 | FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_4_1
      | (FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_10_3_0_1!=4'b0000);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_5_nl
      = MUX_v_3_2_2(3'b000, (inp_lookup_2_FpExpoWidthInc_6U_8U_23U_0U_1U_1_else_acc_nl),
      (IsZero_6U_23U_1_aelse_IsZero_6U_23U_1_or_1_nl));
  assign or_5256_nl = (~ (cfg_precision_1_sva_st_85[1])) | (chn_inp_in_crt_sva_8_739_736_1[1])
      | (cfg_precision_1_sva_st_85[0]);
  assign IsInf_6U_23U_1_aelse_mux_3_nl = MUX_s_1_2_2(IsInf_6U_23U_1_land_2_lpi_1_dfm_mx0w0,
      IsInf_6U_23U_1_land_2_lpi_1_dfm, or_5256_nl);
  assign and_3556_nl = (~ IsInf_6U_23U_1_land_1_lpi_1_dfm_mx0w0) & or_11_cse;
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_mux_48_nl = MUX_v_4_2_2(FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_3_0_1,
      4'b1110, IsInf_6U_23U_1_land_1_lpi_1_dfm_mx0w0);
  assign nl_inp_lookup_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_else_acc_nl = conv_u2u_2_3({1'b1
      , FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_5_1}) + 3'b1;
  assign inp_lookup_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_else_acc_nl = nl_inp_lookup_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_else_acc_nl[2:0];
  assign IsZero_6U_23U_1_aelse_IsZero_6U_23U_1_or_nl = (FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_22_13_1_lpi_1_dfm_mx0w1!=10'b0000000000)
      | (FpMantWidthInc_6U_10U_23U_0U_1U_1_o_mant_9_0_1_lpi_1_dfm!=10'b0000000000)
      | FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_5_1 | FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_4_1
      | (FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_10_3_0_1!=4'b0000);
  assign FpExpoWidthInc_6U_8U_23U_0U_1U_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_and_nl
      = MUX_v_3_2_2(3'b000, (inp_lookup_1_FpExpoWidthInc_6U_8U_23U_0U_1U_1_else_acc_nl),
      (IsZero_6U_23U_1_aelse_IsZero_6U_23U_1_or_nl));
  assign or_5251_nl = (cfg_precision_1_sva_st_85!=2'b10) | (chn_inp_in_crt_sva_8_739_736_1[0]);
  assign IsInf_6U_23U_1_aelse_mux_1_nl = MUX_s_1_2_2(IsInf_6U_23U_1_land_1_lpi_1_dfm_mx0w0,
      IsInf_6U_23U_1_land_1_lpi_1_dfm, or_5251_nl);
  assign mux_1564_nl = MUX_s_1_2_2(mux_tmp_1245, mux_tmp_1485, or_11_cse);
  assign mux_1567_nl = MUX_s_1_2_2(mux_tmp_1233, mux_tmp_1488, or_11_cse);
  assign mux_1570_nl = MUX_s_1_2_2(mux_tmp_1221, and_307_cse, or_11_cse);
  assign mux_1573_nl = MUX_s_1_2_2(mux_tmp_1209, mux_tmp_1494, or_11_cse);
  assign mux_1574_nl = MUX_s_1_2_2(nor_tmp_464, nor_tmp_522, or_11_cse);
  assign or_3533_nl = (chn_inp_in_crt_sva_8_739_736_1[0]) | nand_332_cse;
  assign mux_1579_nl = MUX_s_1_2_2((or_3533_nl), or_tmp_3530, or_11_cse);
  assign or_3537_nl = (chn_inp_in_crt_sva_8_739_736_1[1]) | nand_332_cse;
  assign mux_1580_nl = MUX_s_1_2_2((or_3537_nl), or_tmp_3534, or_11_cse);
  assign or_3541_nl = (chn_inp_in_crt_sva_8_739_736_1[2]) | nand_332_cse;
  assign mux_1581_nl = MUX_s_1_2_2((or_3541_nl), or_tmp_3538, or_11_cse);
  assign or_3545_nl = (chn_inp_in_crt_sva_8_739_736_1[3]) | nand_332_cse;
  assign mux_1582_nl = MUX_s_1_2_2((or_3545_nl), or_tmp_3542, or_11_cse);
  assign mux_1583_nl = MUX_s_1_2_2(mux_tmp_1450, nor_tmp_532, or_11_cse);
  assign mux_1584_nl = MUX_s_1_2_2(mux_tmp_1458, nor_tmp_533, or_11_cse);
  assign mux_1585_nl = MUX_s_1_2_2(mux_tmp_1452, nor_tmp_535, or_11_cse);
  assign mux_1588_nl = MUX_s_1_2_2(mux_tmp_1454, mux_tmp_1509, or_11_cse);
  assign mux_1590_nl = MUX_s_1_2_2(mux_tmp_1485, mux_tmp_1511, or_11_cse);
  assign mux_1592_nl = MUX_s_1_2_2(mux_tmp_1488, mux_tmp_1513, or_11_cse);
  assign mux_1595_nl = MUX_s_1_2_2(and_307_cse, and_312_cse, or_11_cse);
  assign mux_1597_nl = MUX_s_1_2_2(mux_tmp_1494, mux_tmp_1518, or_11_cse);
  assign mux_1598_nl = MUX_s_1_2_2(nor_tmp_522, nor_tmp_545, or_11_cse);
  assign mux_1599_nl = MUX_s_1_2_2(or_tmp_3510, or_tmp_3562, or_11_cse);
  assign mux_1600_nl = MUX_s_1_2_2(or_tmp_3512, or_tmp_3564, or_11_cse);
  assign mux_1601_nl = MUX_s_1_2_2(or_tmp_3514, or_tmp_3566, or_11_cse);
  assign mux_1602_nl = MUX_s_1_2_2(or_tmp_3516, or_tmp_3568, or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_46_nl = (~ FpMul_6U_10U_1_or_11_itm)
      & and_dcpl_655;
  assign nor_921_nl = ~((~ main_stage_v_4) | (cfg_precision_1_sva_st_81!=2'b10) |
      (~((~(FpAdd_6U_10U_1_is_a_greater_acc_itm_6 | (~ inp_lookup_1_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp)))
      | (chn_inp_in_crt_sva_4_739_736_1[0]) | IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_tmp
      | mux_476_cse)));
  assign mux_1604_nl = MUX_s_1_2_2((~ inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5),
      inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5,
      inp_lookup_1_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6);
  assign nor_923_nl = ~((cfg_precision_1_sva_st_82[0]) | (~((cfg_precision_1_sva_st_82[1])
      & main_stage_v_5 & (nor_1593_cse | (chn_inp_in_crt_sva_5_739_736_1[0]) | IsNaN_6U_10U_8_land_1_lpi_1_dfm_6
      | (mux_1604_nl)))));
  assign mux_1605_nl = MUX_s_1_2_2((nor_923_nl), (nor_921_nl), or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_45_nl = (~ FpMul_6U_10U_1_or_10_itm)
      & and_dcpl_663;
  assign nor_917_nl = ~((~ main_stage_v_4) | (cfg_precision_1_sva_st_81!=2'b10) |
      (~((~(FpAdd_6U_10U_1_is_a_greater_acc_1_itm_6 | (~ inp_lookup_2_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp)))
      | (chn_inp_in_crt_sva_4_739_736_1[1]) | IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_1_tmp
      | mux_485_cse)));
  assign mux_1607_nl = MUX_s_1_2_2((~ inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5),
      inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5,
      inp_lookup_2_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_6);
  assign nor_919_nl = ~((~ main_stage_v_5) | (cfg_precision_1_sva_st_82[0]) | (~((cfg_precision_1_sva_st_82[1])
      & (nor_1587_cse | (chn_inp_in_crt_sva_5_739_736_1[1]) | IsNaN_6U_10U_8_land_2_lpi_1_dfm_4
      | (mux_1607_nl)))));
  assign mux_1608_nl = MUX_s_1_2_2((nor_919_nl), (nor_917_nl), or_11_cse);
  assign FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_mant_and_44_nl = (~ FpMul_6U_10U_1_or_8_itm)
      & and_dcpl_679;
  assign nor_911_nl = ~((~ main_stage_v_4) | (cfg_precision_1_sva_st_81!=2'b10) |
      (~((~(FpAdd_6U_10U_1_is_a_greater_acc_3_itm_6_1 | (~ inp_lookup_4_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp)))
      | (chn_inp_in_crt_sva_4_739_736_1[3]) | IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_3_tmp
      | mux_1140_cse)));
  assign nor_913_nl = ~((~ main_stage_v_5) | (cfg_precision_1_sva_st_82!=2'b10));
  assign and_3394_nl = inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
      & main_stage_v_5 & (cfg_precision_1_sva_st_82==2'b10);
  assign nor_915_nl = ~(inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_5
      | (~ main_stage_v_5) | (cfg_precision_1_sva_st_82!=2'b10));
  assign mux_1610_nl = MUX_s_1_2_2((nor_915_nl), (and_3394_nl), inp_lookup_4_FpAdd_6U_10U_1_is_addition_FpAdd_6U_10U_1_is_addition_xnor_svs_st_5);
  assign or_3596_nl = nor_1130_cse | (chn_inp_in_crt_sva_5_739_736_1[3]) | IsNaN_6U_10U_8_land_lpi_1_dfm_4;
  assign mux_1611_nl = MUX_s_1_2_2((mux_1610_nl), (nor_913_nl), or_3596_nl);
  assign mux_1612_nl = MUX_s_1_2_2((mux_1611_nl), (nor_911_nl), or_11_cse);
  assign mux_1613_nl = MUX_s_1_2_2(nor_tmp_532, nor_tmp_551, or_11_cse);
  assign mux_1614_nl = MUX_s_1_2_2(nor_tmp_535, nor_tmp_552, or_11_cse);
  assign mux_1615_nl = MUX_s_1_2_2(mux_tmp_1509, nor_tmp_553, or_11_cse);
  assign mux_1616_nl = MUX_s_1_2_2(nor_tmp_533, nor_tmp_555, or_11_cse);
  assign mux_1617_nl = MUX_s_1_2_2(or_tmp_3542, or_tmp_3612, or_11_cse);
  assign mux_1618_nl = MUX_s_1_2_2(or_tmp_3538, or_tmp_3614, or_11_cse);
  assign mux_1619_nl = MUX_s_1_2_2(or_tmp_3534, or_tmp_3616, or_11_cse);
  assign mux_1620_nl = MUX_s_1_2_2(or_tmp_3530, or_tmp_3618, or_11_cse);
  assign mux_1622_nl = MUX_s_1_2_2(mux_tmp_1511, mux_tmp_1543, or_11_cse);
  assign mux_1624_nl = MUX_s_1_2_2(mux_tmp_1513, mux_tmp_1545, or_11_cse);
  assign mux_1629_nl = MUX_s_1_2_2(and_312_cse, mux_tmp_1548, or_11_cse);
  assign mux_1632_nl = MUX_s_1_2_2(mux_tmp_1518, mux_tmp_1553, or_11_cse);
  assign mux_1633_nl = MUX_s_1_2_2(nor_tmp_545, nor_tmp_569, or_11_cse);
  assign mux_1634_nl = MUX_s_1_2_2(or_tmp_3562, or_tmp_3627, or_11_cse);
  assign mux_1635_nl = MUX_s_1_2_2(or_tmp_3564, or_tmp_3629, or_11_cse);
  assign mux_1636_nl = MUX_s_1_2_2(or_tmp_3566, or_tmp_3631, or_11_cse);
  assign mux_1637_nl = MUX_s_1_2_2(or_tmp_3568, or_tmp_3633, or_11_cse);
  assign mux_1638_nl = MUX_s_1_2_2((FpMul_6U_10U_1_p_mant_p1_1_sva[21]), nor_905_cse,
      nor_1210_cse);
  assign nor_902_nl = ~((~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10) |
      (~((chn_inp_in_crt_sva_3_739_736_1[0]) | IsNaN_6U_10U_5_land_1_lpi_1_dfm_5
      | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_15 | (~((~ inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4)
      | FpMul_6U_10U_1_lor_6_lpi_1_dfm_5 | (mux_1638_nl))))));
  assign nor_907_nl = ~(nor_908_cse | (~ FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_1_st_2)
      | FpMul_6U_10U_1_lor_6_lpi_1_dfm_6 | (~ main_stage_v_4) | (cfg_precision_1_sva_st_81!=2'b10));
  assign or_3645_nl = (chn_inp_in_crt_sva_4_739_736_1[0]) | IsNaN_6U_10U_5_land_1_lpi_1_dfm_6
      | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_16;
  assign mux_1639_nl = MUX_s_1_2_2((nor_907_nl), nor_1221_cse, or_3645_nl);
  assign mux_1640_nl = MUX_s_1_2_2((mux_1639_nl), (nor_902_nl), or_11_cse);
  assign mux_1641_nl = MUX_s_1_2_2((FpMul_6U_10U_1_p_mant_p1_2_sva[21]), nor_898_cse,
      nor_1193_cse);
  assign nor_895_nl = ~((~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10) |
      (~((chn_inp_in_crt_sva_3_739_736_1[1]) | IsNaN_6U_10U_5_land_2_lpi_1_dfm_5
      | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_15 | (~((~ inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4)
      | FpMul_6U_10U_1_lor_7_lpi_1_dfm_5 | (mux_1641_nl))))));
  assign nor_900_nl = ~(nor_901_cse | (~ FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_1_st_2)
      | FpMul_6U_10U_1_lor_7_lpi_1_dfm_6 | (~ main_stage_v_4) | (cfg_precision_1_sva_st_81!=2'b10));
  assign or_3660_nl = (chn_inp_in_crt_sva_4_739_736_1[1]) | IsNaN_6U_10U_5_land_2_lpi_1_dfm_6
      | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_16;
  assign mux_1642_nl = MUX_s_1_2_2((nor_900_nl), nor_1221_cse, or_3660_nl);
  assign mux_1643_nl = MUX_s_1_2_2((mux_1642_nl), (nor_895_nl), or_11_cse);
  assign mux_1644_nl = MUX_s_1_2_2((~ (FpMul_6U_10U_1_p_mant_p1_sva[21])), or_5689_cse,
      nor_572_cse);
  assign nor_889_nl = ~((~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10) |
      (~((chn_inp_in_crt_sva_3_739_736_1[3]) | IsNaN_6U_10U_5_land_lpi_1_dfm_5 |
      IsNaN_6U_10U_2_land_lpi_1_dfm_st_15 | (~(FpMul_6U_10U_1_lor_1_lpi_1_dfm_5 |
      (~(inp_lookup_4_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs_2
      & (mux_1644_nl))))))));
  assign nor_893_nl = ~(nor_894_cse | (~ FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_1_st_2)
      | FpMul_6U_10U_1_lor_1_lpi_1_dfm_6 | (~ main_stage_v_4) | (cfg_precision_1_sva_st_81!=2'b10));
  assign or_3674_nl = (chn_inp_in_crt_sva_4_739_736_1[3]) | IsNaN_6U_10U_4_land_lpi_1_dfm_5
      | IsNaN_6U_10U_5_land_lpi_1_dfm_6;
  assign mux_1645_nl = MUX_s_1_2_2((nor_893_nl), nor_1221_cse, or_3674_nl);
  assign mux_1646_nl = MUX_s_1_2_2((mux_1645_nl), (nor_889_nl), or_11_cse);
  assign mux_1647_nl = MUX_s_1_2_2(nor_tmp_551, and_tmp_225, or_11_cse);
  assign mux_1648_nl = MUX_s_1_2_2(nor_tmp_555, and_tmp_226, or_11_cse);
  assign mux_1649_nl = MUX_s_1_2_2(nor_tmp_552, and_tmp_227, or_11_cse);
  assign mux_1650_nl = MUX_s_1_2_2(nor_tmp_553, and_tmp_228, or_11_cse);
  assign mux_1652_nl = MUX_s_1_2_2(or_tmp_3612, mux_tmp_1573, or_11_cse);
  assign mux_1654_nl = MUX_s_1_2_2(or_tmp_3614, mux_tmp_1575, or_11_cse);
  assign mux_1656_nl = MUX_s_1_2_2(or_tmp_3616, mux_tmp_1577, or_11_cse);
  assign mux_1658_nl = MUX_s_1_2_2(or_tmp_3618, mux_tmp_1579, or_11_cse);
  assign mux_1660_nl = MUX_s_1_2_2(mux_tmp_1543, mux_tmp_1581, or_11_cse);
  assign mux_1662_nl = MUX_s_1_2_2(mux_tmp_1545, mux_tmp_1583, or_11_cse);
  assign mux_1664_nl = MUX_s_1_2_2(mux_tmp_1548, mux_tmp_1585, or_11_cse);
  assign mux_1666_nl = MUX_s_1_2_2(mux_tmp_1553, mux_tmp_1587, or_11_cse);
  assign and_3089_nl = ((chn_inp_in_crt_sva_5_739_736_1!=4'b0000)) & main_stage_v_5;
  assign mux_1667_nl = MUX_s_1_2_2(nor_tmp_569, (and_3089_nl), or_11_cse);
  assign mux_1668_nl = MUX_s_1_2_2(or_tmp_3627, or_3716_cse, or_11_cse);
  assign mux_1669_nl = MUX_s_1_2_2(or_tmp_3629, or_3718_cse, or_11_cse);
  assign mux_1670_nl = MUX_s_1_2_2(or_tmp_3631, or_3720_cse, or_11_cse);
  assign mux_1671_nl = MUX_s_1_2_2(or_tmp_3633, or_3722_cse, or_11_cse);
  assign mux_1673_nl = MUX_s_1_2_2(mux_tmp_1579, nand_tmp_218, or_11_cse);
  assign mux_1675_nl = MUX_s_1_2_2(mux_tmp_1577, nand_tmp_219, or_11_cse);
  assign mux_1677_nl = MUX_s_1_2_2(mux_tmp_1575, nand_tmp_220, or_11_cse);
  assign mux_1679_nl = MUX_s_1_2_2(mux_tmp_1573, nand_tmp_221, or_11_cse);
  assign nand_320_nl = ~((~ IsNaN_6U_10U_4_nor_tmp) & inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_5_1
      & (inp_lookup_else_if_a0_15_10_1_lpi_1_dfm_6_4_0_1==5'b11111) & IsNaN_8U_23U_land_1_lpi_1_dfm_st_4
      & (~ (chn_inp_in_crt_sva_2_739_736_1[0])));
  assign mux_1680_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_2_739_736_1[0]), (nand_320_nl),
      and_3246_cse);
  assign nor_881_nl = ~((~ main_stage_v_2) | (cfg_precision_1_sva_st_91[0]) | (~((cfg_precision_1_sva_st_91[1])
      & (nor_35_cse | (mux_1680_nl)))));
  assign nor_883_nl = ~(FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_3 | (~ inp_lookup_1_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs)
      | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10));
  assign or_3742_nl = nor_884_cse | (chn_inp_in_crt_sva_3_739_736_1[0]);
  assign mux_1681_nl = MUX_s_1_2_2((nor_883_nl), nor_1217_cse, or_3742_nl);
  assign mux_1682_nl = MUX_s_1_2_2((mux_1681_nl), (nor_881_nl), or_11_cse);
  assign nand_318_nl = ~((~ IsNaN_6U_10U_4_nor_1_tmp) & inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_6_5_1
      & (inp_lookup_else_if_a0_15_10_2_lpi_1_dfm_6_4_0_1==5'b11111) & IsNaN_8U_23U_land_2_lpi_1_dfm_st_4
      & (~ (chn_inp_in_crt_sva_2_739_736_1[1])));
  assign mux_1683_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_2_739_736_1[1]), (nand_318_nl),
      and_3244_cse);
  assign nor_876_nl = ~((~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10) |
      (~(nor_584_cse | (mux_1683_nl))));
  assign nor_879_nl = ~(FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_3 | (~ inp_lookup_2_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs)
      | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10));
  assign or_3753_nl = nor_880_cse | (chn_inp_in_crt_sva_3_739_736_1[1]);
  assign mux_1684_nl = MUX_s_1_2_2((nor_879_nl), nor_1217_cse, or_3753_nl);
  assign mux_1685_nl = MUX_s_1_2_2((mux_1684_nl), (nor_876_nl), or_11_cse);
  assign nand_317_nl = ~((~ IsNaN_6U_10U_4_nor_3_tmp) & inp_lookup_else_if_a0_15_10_lpi_1_dfm_6_5_1
      & (inp_lookup_else_if_a0_15_10_lpi_1_dfm_6_4_0_1==5'b11111) & IsNaN_8U_23U_land_lpi_1_dfm_st_4
      & (~ (chn_inp_in_crt_sva_2_739_736_1[3])));
  assign mux_1686_nl = MUX_s_1_2_2((chn_inp_in_crt_sva_2_739_736_1[3]), (nand_317_nl),
      and_3240_cse);
  assign nor_871_nl = ~((~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10) |
      (~(nor_586_cse | (mux_1686_nl))));
  assign nor_874_nl = ~(FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_3 | (~ inp_lookup_4_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs)
      | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10));
  assign or_3764_nl = nor_875_cse | (chn_inp_in_crt_sva_3_739_736_1[3]);
  assign mux_1687_nl = MUX_s_1_2_2((nor_874_nl), nor_1217_cse, or_3764_nl);
  assign mux_1688_nl = MUX_s_1_2_2((mux_1687_nl), (nor_871_nl), or_11_cse);
  assign and_336_nl = main_stage_v_3 & (chn_inp_in_crt_sva_3_739_736_1[0]);
  assign mux_1689_nl = MUX_s_1_2_2(and_tmp_225, (and_336_nl), or_11_cse);
  assign and_337_nl = main_stage_v_3 & (chn_inp_in_crt_sva_3_739_736_1[3]);
  assign mux_1691_nl = MUX_s_1_2_2(and_tmp_226, (and_337_nl), or_11_cse);
  assign and_338_nl = main_stage_v_3 & (chn_inp_in_crt_sva_3_739_736_1[1]);
  assign mux_1692_nl = MUX_s_1_2_2(and_tmp_227, (and_338_nl), or_11_cse);
  assign and_339_nl = main_stage_v_3 & (chn_inp_in_crt_sva_3_739_736_1[2]);
  assign mux_1693_nl = MUX_s_1_2_2(and_tmp_228, (and_339_nl), or_11_cse);
  assign mux_1695_nl = MUX_s_1_2_2(nand_tmp_222, nand_661_cse, or_11_cse);
  assign mux_1696_nl = MUX_s_1_2_2(nand_tmp_222, or_2282_cse, or_11_cse);
  assign mux_1697_nl = MUX_s_1_2_2((mux_1696_nl), (mux_1695_nl), or_3779_cse);
  assign nor_860_nl = ~((chn_inp_in_crt_sva_3_739_736_1[0]) | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_15);
  assign or_5649_nl = (~((~((~ inp_lookup_1_FpAdd_8U_23U_1_is_a_greater_oif_equal_tmp)
      | FpAdd_8U_23U_1_is_a_greater_oif_aelse_acc_itm_23_1)) | FpAdd_8U_23U_1_is_a_greater_acc_itm_8_1))
      | IsNaN_8U_23U_3_IsNaN_8U_23U_3_nor_tmp;
  assign or_3788_nl = nor_905_cse | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_15;
  assign or_3789_nl = (FpMul_6U_10U_1_p_mant_p1_1_sva[21]) | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_15;
  assign mux_1699_nl = MUX_s_1_2_2((or_3789_nl), (or_3788_nl), nor_1210_cse);
  assign nor_862_nl = ~((~ inp_lookup_1_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4)
      | FpMul_6U_10U_1_lor_6_lpi_1_dfm_5 | (mux_1699_nl));
  assign mux_1700_nl = MUX_s_1_2_2((nor_862_nl), (or_5649_nl), chn_inp_in_crt_sva_3_739_736_1[0]);
  assign mux_1701_nl = MUX_s_1_2_2((mux_1700_nl), (nor_860_nl), IsNaN_6U_10U_5_land_1_lpi_1_dfm_5);
  assign and_3084_nl = nor_1217_cse & (mux_1701_nl);
  assign nor_864_nl = ~((~(FpMul_6U_10U_1_lor_6_lpi_1_dfm_st_4 | (~ FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_5)))
      | IsNaN_6U_10U_5_land_1_lpi_1_dfm_6);
  assign nor_865_nl = ~(IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_16 | (~((~(nor_908_cse
      | (~ FpAdd_8U_23U_1_is_a_greater_lor_1_lpi_1_dfm_1_st_2) | FpMul_6U_10U_1_lor_6_lpi_1_dfm_6))
      | IsNaN_6U_10U_5_land_1_lpi_1_dfm_6)));
  assign mux_1702_nl = MUX_s_1_2_2((nor_865_nl), (nor_864_nl), chn_inp_in_crt_sva_4_739_736_1[0]);
  assign and_3085_nl = nor_1221_cse & (mux_1702_nl);
  assign mux_1703_nl = MUX_s_1_2_2((and_3085_nl), (and_3084_nl), or_11_cse);
  assign mux_1705_nl = MUX_s_1_2_2(or_tmp_3802, or_tmp_3798, chn_inp_in_crt_sva_3_739_736_1[1]);
  assign or_3798_nl = IsNaN_6U_10U_5_land_2_lpi_1_dfm_5 | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_1706_nl = MUX_s_1_2_2(or_tmp_3798, (or_3798_nl), IsNaN_8U_23U_3_IsNaN_8U_23U_3_nor_1_tmp);
  assign or_3809_nl = (~((~(nor_898_cse | (~ inp_lookup_2_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4)
      | FpMul_6U_10U_1_lor_7_lpi_1_dfm_5)) | IsNaN_6U_10U_5_land_2_lpi_1_dfm_5))
      | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_15 | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_1707_nl = MUX_s_1_2_2(or_tmp_3802, (or_3809_nl), inp_lookup_2_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs);
  assign mux_1708_nl = MUX_s_1_2_2((mux_1707_nl), (mux_1706_nl), chn_inp_in_crt_sva_3_739_736_1[1]);
  assign mux_1709_nl = MUX_s_1_2_2((mux_1708_nl), (mux_1705_nl), FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_3);
  assign nor_853_nl = ~((~(FpMul_6U_10U_1_lor_7_lpi_1_dfm_st_4 | (~ FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_5)))
      | IsNaN_6U_10U_5_land_2_lpi_1_dfm_6);
  assign nor_854_nl = ~(IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_16 | (~((~(nor_901_cse
      | (~ FpAdd_8U_23U_1_is_a_greater_lor_2_lpi_1_dfm_1_st_2) | FpMul_6U_10U_1_lor_7_lpi_1_dfm_6))
      | IsNaN_6U_10U_5_land_2_lpi_1_dfm_6)));
  assign mux_1710_nl = MUX_s_1_2_2((nor_854_nl), (nor_853_nl), chn_inp_in_crt_sva_4_739_736_1[1]);
  assign nand_226_nl = ~(nor_1221_cse & (mux_1710_nl));
  assign mux_1711_nl = MUX_s_1_2_2((nand_226_nl), (mux_1709_nl), or_11_cse);
  assign or_3817_nl = (chn_inp_in_crt_sva_3_739_736_1[2]) | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_15
      | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10);
  assign mux_1713_nl = MUX_s_1_2_2(or_tmp_3819, or_2282_cse, IsNaN_8U_23U_3_IsNaN_8U_23U_3_nor_2_tmp);
  assign mux_1714_nl = MUX_s_1_2_2((mux_1713_nl), or_tmp_3819, FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_3);
  assign or_3825_nl = (~((~ (inp_lookup_3_FpMul_6U_10U_1_p_mant_p1_mul_tmp[21]))
      | inp_lookup_3_FpMul_6U_10U_1_else_2_else_if_if_acc_1_itm_5_1)) | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_15
      | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10);
  assign or_3827_nl = (FpMul_6U_10U_1_p_mant_p1_3_sva[21]) | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_15
      | (~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10);
  assign nor_600_nl = ~(FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_3 | (~ inp_lookup_3_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs));
  assign mux_1715_nl = MUX_s_1_2_2((or_3827_nl), (or_3825_nl), nor_600_nl);
  assign or_3828_nl = (~ inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_st_4)
      | FpMul_6U_10U_1_lor_8_lpi_1_dfm_5 | (mux_1715_nl);
  assign mux_1716_nl = MUX_s_1_2_2((or_3828_nl), (mux_1714_nl), chn_inp_in_crt_sva_3_739_736_1[2]);
  assign mux_1717_nl = MUX_s_1_2_2((mux_1716_nl), (or_3817_nl), IsNaN_6U_10U_5_land_3_lpi_1_dfm_5);
  assign nor_845_nl = ~((~(FpMul_6U_10U_1_lor_8_lpi_1_dfm_st_4 | (~ FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_5)))
      | IsNaN_6U_10U_5_land_3_lpi_1_dfm_6);
  assign nor_846_nl = ~(IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_16 | (~((~((~((~ FpExpoWidthInc_5U_6U_10U_1U_1U_2_o_expo_5_4_3_lpi_1_dfm_9_1)
      | inp_lookup_3_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_FpAdd_8U_23U_1_is_addition_xor_svs_5))
      | (~ FpAdd_8U_23U_1_is_a_greater_lor_3_lpi_1_dfm_1_st_2) | FpMul_6U_10U_1_lor_8_lpi_1_dfm_6))
      | IsNaN_6U_10U_5_land_3_lpi_1_dfm_6)));
  assign mux_1718_nl = MUX_s_1_2_2((nor_846_nl), (nor_845_nl), chn_inp_in_crt_sva_4_739_736_1[2]);
  assign nand_227_nl = ~(nor_1221_cse & (mux_1718_nl));
  assign mux_1719_nl = MUX_s_1_2_2((nand_227_nl), (mux_1717_nl), or_11_cse);
  assign or_3836_nl = FpAdd_8U_23U_1_is_a_greater_acc_3_itm_8_1 | IsNaN_6U_10U_5_land_lpi_1_dfm_5;
  assign mux_1720_nl = MUX_s_1_2_2((or_3836_nl), IsNaN_6U_10U_5_land_lpi_1_dfm_5,
      nor_605_cse);
  assign mux_1721_nl = MUX_s_1_2_2(or_tmp_3836, (mux_1720_nl), chn_inp_in_crt_sva_3_739_736_1[3]);
  assign or_3840_nl = nor_605_cse | FpAdd_8U_23U_1_is_a_greater_acc_3_itm_8_1 | IsNaN_6U_10U_5_land_lpi_1_dfm_5;
  assign or_3839_nl = IsNaN_8U_23U_3_IsNaN_8U_23U_3_nand_3_tmp | IsNaN_8U_23U_3_nor_3_tmp;
  assign mux_1722_nl = MUX_s_1_2_2(IsNaN_6U_10U_5_land_lpi_1_dfm_5, (or_3840_nl),
      or_3839_nl);
  assign or_3843_nl = (~((~((~((~ (inp_lookup_4_FpMul_6U_10U_1_p_mant_p1_mul_tmp[21]))
      | inp_lookup_4_FpMul_6U_10U_1_else_2_else_if_if_acc_1_itm_5_1)) | FpMul_6U_10U_1_lor_1_lpi_1_dfm_5
      | (~ inp_lookup_4_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs_2)))
      | IsNaN_6U_10U_5_land_lpi_1_dfm_5)) | IsNaN_6U_10U_2_land_lpi_1_dfm_st_15;
  assign mux_1723_nl = MUX_s_1_2_2(or_tmp_3836, (or_3843_nl), inp_lookup_4_FpMul_6U_10U_1_else_2_if_slc_FpMul_6U_10U_1_else_2_if_acc_6_svs);
  assign mux_1724_nl = MUX_s_1_2_2((mux_1723_nl), (mux_1722_nl), chn_inp_in_crt_sva_3_739_736_1[3]);
  assign mux_1725_nl = MUX_s_1_2_2((mux_1724_nl), (mux_1721_nl), FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_3);
  assign nor_836_nl = ~((~ main_stage_v_3) | (cfg_precision_1_sva_st_80!=2'b10) |
      (mux_1725_nl));
  assign nor_839_nl = ~(FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5 | FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_4
      | (~ main_stage_v_4) | (cfg_precision_1_sva_st_81!=2'b10));
  assign nor_840_nl = ~((or_tmp_2441 & FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_5)
      | FpMul_6U_10U_1_lor_1_lpi_1_dfm_st_4 | (~ main_stage_v_4) | (cfg_precision_1_sva_st_81!=2'b10));
  assign mux_1726_nl = MUX_s_1_2_2((nor_840_nl), (nor_839_nl), IsNaN_8U_23U_2_land_lpi_1_dfm_st_7);
  assign or_3853_nl = nor_894_cse | (~ FpAdd_8U_23U_1_is_a_greater_lor_lpi_1_dfm_1_st_2)
      | FpMul_6U_10U_1_lor_1_lpi_1_dfm_6 | (~ main_stage_v_4) | (cfg_precision_1_sva_st_81!=2'b10);
  assign mux_1727_nl = MUX_s_1_2_2((or_3853_nl), or_3850_cse, IsNaN_6U_10U_5_land_lpi_1_dfm_6);
  assign nor_841_nl = ~(IsNaN_6U_10U_4_land_lpi_1_dfm_5 | (mux_1727_nl));
  assign mux_1728_nl = MUX_s_1_2_2((nor_841_nl), (mux_1726_nl), chn_inp_in_crt_sva_4_739_736_1[3]);
  assign mux_1729_nl = MUX_s_1_2_2((mux_1728_nl), (nor_836_nl), or_11_cse);
  assign mux_1731_nl = MUX_s_1_2_2(mux_tmp_1581, and_tmp_240, or_11_cse);
  assign mux_1733_nl = MUX_s_1_2_2(mux_tmp_1583, and_tmp_242, or_11_cse);
  assign mux_1735_nl = MUX_s_1_2_2(mux_tmp_1585, and_tmp_244, or_11_cse);
  assign mux_1737_nl = MUX_s_1_2_2(mux_tmp_1587, and_tmp_246, or_11_cse);
  assign nor_833_nl = ~((~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[0])
      | (cfg_precision_1_sva_st_81!=2'b10) | ((~((~ IsNaN_6U_10U_9_nor_tmp) & FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_5_1
      & FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_4_1 & (FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_3_0_1==4'b1111)))
      & FpAdd_6U_10U_1_is_a_greater_acc_itm_6) | IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_tmp);
  assign or_3867_nl = (~ main_stage_v_5) | IsNaN_6U_10U_8_land_1_lpi_1_dfm_6;
  assign or_3870_nl = IsNaN_8U_23U_3_land_1_lpi_1_dfm_6 | (~ main_stage_v_5) | IsNaN_6U_10U_8_land_1_lpi_1_dfm_6;
  assign mux_1742_nl = MUX_s_1_2_2((or_3870_nl), (or_3867_nl), IsNaN_6U_10U_9_land_1_lpi_1_dfm_6);
  assign nor_1944_nl = ~((cfg_precision_1_sva_st_82!=2'b10) | (mux_1742_nl) | (chn_inp_in_crt_sva_5_739_736_1[0]));
  assign mux_1744_nl = MUX_s_1_2_2((nor_1944_nl), (nor_833_nl), or_11_cse);
  assign nor_825_nl = ~((~ IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_tmp) | (~ main_stage_v_4)
      | (chn_inp_in_crt_sva_4_739_736_1[0]) | (cfg_precision_1_sva_st_81!=2'b10));
  assign nor_826_nl = ~((~(FpAdd_6U_10U_1_is_a_greater_acc_itm_6 | inp_lookup_1_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp
      | IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_tmp)) | (~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[0])
      | (cfg_precision_1_sva_st_81!=2'b10));
  assign and_3081_nl = (~ IsNaN_6U_10U_9_nor_tmp) & FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_5_1
      & FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_4_1 & (FpMul_6U_10U_2_o_expo_1_lpi_1_dfm_6_3_0_1==4'b1111);
  assign mux_1745_nl = MUX_s_1_2_2((nor_826_nl), (nor_825_nl), and_3081_nl);
  assign nor_828_nl = ~((~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[0])
      | (cfg_precision_1_sva_st_81!=2'b10));
  assign mux_1746_nl = MUX_s_1_2_2((nor_828_nl), (mux_1745_nl), nor_956_cse);
  assign nand_779_nl = ~((nor_1593_cse | IsNaN_6U_10U_8_land_1_lpi_1_dfm_6) & main_stage_v_5);
  assign mux_1747_nl = MUX_s_1_2_2(or_3885_cse, (nand_779_nl), IsNaN_8U_23U_2_land_1_lpi_1_dfm_9);
  assign mux_1748_nl = MUX_s_1_2_2((mux_1747_nl), or_3722_cse, IsNaN_8U_23U_3_land_1_lpi_1_dfm_6);
  assign mux_1749_nl = MUX_s_1_2_2(or_3885_cse, (mux_1748_nl), nor_623_cse);
  assign mux_1750_nl = MUX_s_1_2_2((mux_1749_nl), or_3885_cse, IsNaN_6U_10U_9_land_1_lpi_1_dfm_6);
  assign nor_1953_nl = ~((cfg_precision_1_sva_st_82!=2'b10) | (mux_1750_nl) | (chn_inp_in_crt_sva_5_739_736_1[0]));
  assign mux_1752_nl = MUX_s_1_2_2((nor_1953_nl), (mux_1746_nl), or_11_cse);
  assign nor_822_nl = ~((~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[1])
      | (cfg_precision_1_sva_st_81!=2'b10) | ((~((~ IsNaN_6U_10U_9_nor_1_tmp) & FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_5_1
      & FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_4_1 & (FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_3_0_1==4'b1111)))
      & FpAdd_6U_10U_1_is_a_greater_acc_1_itm_6) | IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_1_tmp);
  assign or_3895_nl = (~ main_stage_v_5) | IsNaN_6U_10U_8_land_2_lpi_1_dfm_4;
  assign or_3898_nl = IsNaN_8U_23U_3_land_2_lpi_1_dfm_6 | (~ main_stage_v_5) | IsNaN_6U_10U_8_land_2_lpi_1_dfm_4;
  assign mux_1757_nl = MUX_s_1_2_2((or_3898_nl), (or_3895_nl), IsNaN_6U_10U_9_land_2_lpi_1_dfm_6);
  assign nor_1939_nl = ~((cfg_precision_1_sva_st_82!=2'b10) | (mux_1757_nl) | (chn_inp_in_crt_sva_5_739_736_1[1]));
  assign mux_1759_nl = MUX_s_1_2_2((nor_1939_nl), (nor_822_nl), or_11_cse);
  assign nor_814_nl = ~((~ IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_1_tmp) | (~ main_stage_v_4)
      | (chn_inp_in_crt_sva_4_739_736_1[1]) | (cfg_precision_1_sva_st_81!=2'b10));
  assign nor_815_nl = ~((~(FpAdd_6U_10U_1_is_a_greater_acc_1_itm_6 | inp_lookup_2_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp
      | IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_1_tmp)) | (~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[1])
      | (cfg_precision_1_sva_st_81!=2'b10));
  assign and_3079_nl = (~ IsNaN_6U_10U_9_nor_1_tmp) & FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_5_1
      & FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_4_1 & (FpMul_6U_10U_2_o_expo_2_lpi_1_dfm_6_3_0_1==4'b1111);
  assign mux_1760_nl = MUX_s_1_2_2((nor_815_nl), (nor_814_nl), and_3079_nl);
  assign nor_817_nl = ~((~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[1])
      | (cfg_precision_1_sva_st_81!=2'b10));
  assign mux_1761_nl = MUX_s_1_2_2((nor_817_nl), (mux_1760_nl), nor_956_cse);
  assign nand_778_nl = ~((nor_1587_cse | IsNaN_6U_10U_8_land_2_lpi_1_dfm_4) & main_stage_v_5);
  assign mux_1762_nl = MUX_s_1_2_2(or_3913_cse, (nand_778_nl), IsNaN_8U_23U_2_land_2_lpi_1_dfm_9);
  assign mux_1763_nl = MUX_s_1_2_2((mux_1762_nl), or_3720_cse, IsNaN_8U_23U_3_land_2_lpi_1_dfm_6);
  assign mux_1764_nl = MUX_s_1_2_2(or_3913_cse, (mux_1763_nl), nor_623_cse);
  assign mux_1765_nl = MUX_s_1_2_2((mux_1764_nl), or_3913_cse, IsNaN_6U_10U_9_land_2_lpi_1_dfm_6);
  assign nor_1952_nl = ~((cfg_precision_1_sva_st_82!=2'b10) | (mux_1765_nl) | (chn_inp_in_crt_sva_5_739_736_1[1]));
  assign mux_1767_nl = MUX_s_1_2_2((nor_1952_nl), (mux_1761_nl), or_11_cse);
  assign nor_811_nl = ~((~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[2])
      | (cfg_precision_1_sva_st_81!=2'b10) | ((~((~ IsNaN_6U_10U_9_nor_2_tmp) & FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_5_1
      & FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_4_1 & (FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_3_0_1==4'b1111)))
      & FpAdd_6U_10U_1_is_a_greater_acc_2_itm_6) | IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_2_tmp);
  assign or_3923_nl = (~ main_stage_v_5) | IsNaN_6U_10U_8_land_3_lpi_1_dfm_4;
  assign or_3926_nl = IsNaN_8U_23U_3_land_3_lpi_1_dfm_6 | (~ main_stage_v_5) | IsNaN_6U_10U_8_land_3_lpi_1_dfm_4;
  assign mux_1772_nl = MUX_s_1_2_2((or_3926_nl), (or_3923_nl), IsNaN_6U_10U_9_land_3_lpi_1_dfm_6);
  assign nor_1935_nl = ~((cfg_precision_1_sva_st_82!=2'b10) | (mux_1772_nl) | (chn_inp_in_crt_sva_5_739_736_1[2]));
  assign mux_1774_nl = MUX_s_1_2_2((nor_1935_nl), (nor_811_nl), or_11_cse);
  assign nor_803_nl = ~((~ IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_2_tmp) | (~ main_stage_v_4)
      | (chn_inp_in_crt_sva_4_739_736_1[2]) | (cfg_precision_1_sva_st_81!=2'b10));
  assign nor_804_nl = ~((~(FpAdd_6U_10U_1_is_a_greater_acc_2_itm_6 | inp_lookup_3_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp
      | IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_2_tmp)) | (~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[2])
      | (cfg_precision_1_sva_st_81!=2'b10));
  assign and_3077_nl = (~ IsNaN_6U_10U_9_nor_2_tmp) & FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_5_1
      & FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_4_1 & (FpMul_6U_10U_2_o_expo_3_lpi_1_dfm_6_3_0_1==4'b1111);
  assign mux_1775_nl = MUX_s_1_2_2((nor_804_nl), (nor_803_nl), and_3077_nl);
  assign nor_806_nl = ~((~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[2])
      | (cfg_precision_1_sva_st_81!=2'b10));
  assign mux_1776_nl = MUX_s_1_2_2((nor_806_nl), (mux_1775_nl), nor_956_cse);
  assign nand_777_nl = ~((nor_1584_cse | IsNaN_6U_10U_8_land_3_lpi_1_dfm_4) & main_stage_v_5);
  assign mux_1777_nl = MUX_s_1_2_2(or_3941_cse, (nand_777_nl), IsNaN_8U_23U_2_land_3_lpi_1_dfm_9);
  assign mux_1778_nl = MUX_s_1_2_2((mux_1777_nl), or_3718_cse, IsNaN_8U_23U_3_land_3_lpi_1_dfm_6);
  assign mux_1779_nl = MUX_s_1_2_2(or_3941_cse, (mux_1778_nl), nor_623_cse);
  assign mux_1780_nl = MUX_s_1_2_2((mux_1779_nl), or_3941_cse, IsNaN_6U_10U_9_land_3_lpi_1_dfm_6);
  assign nor_1951_nl = ~((cfg_precision_1_sva_st_82!=2'b10) | (mux_1780_nl) | (chn_inp_in_crt_sva_5_739_736_1[2]));
  assign mux_1782_nl = MUX_s_1_2_2((nor_1951_nl), (mux_1776_nl), or_11_cse);
  assign nor_800_nl = ~((~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[3])
      | (cfg_precision_1_sva_st_81!=2'b10) | ((~((~ IsNaN_6U_10U_9_nor_3_tmp) & FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_5_1
      & FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_4_1 & (FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_3_0_1==4'b1111)))
      & FpAdd_6U_10U_1_is_a_greater_acc_3_itm_6_1) | IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_3_tmp);
  assign or_3951_nl = (~ main_stage_v_5) | IsNaN_6U_10U_8_land_lpi_1_dfm_4;
  assign or_3954_nl = IsNaN_8U_23U_3_land_lpi_1_dfm_5 | (~ main_stage_v_5) | IsNaN_6U_10U_8_land_lpi_1_dfm_4;
  assign mux_1787_nl = MUX_s_1_2_2((or_3954_nl), (or_3951_nl), IsNaN_6U_10U_9_land_lpi_1_dfm_6);
  assign nor_1931_nl = ~((cfg_precision_1_sva_st_82!=2'b10) | (mux_1787_nl) | (chn_inp_in_crt_sva_5_739_736_1[3]));
  assign mux_1789_nl = MUX_s_1_2_2((nor_1931_nl), (nor_800_nl), or_11_cse);
  assign nor_792_nl = ~((~ IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_3_tmp) | (~ main_stage_v_4)
      | (chn_inp_in_crt_sva_4_739_736_1[3]) | (cfg_precision_1_sva_st_81!=2'b10));
  assign nor_793_nl = ~((~(FpAdd_6U_10U_1_is_a_greater_acc_3_itm_6_1 | inp_lookup_4_FpAdd_6U_10U_1_is_a_greater_oif_equal_tmp
      | IsNaN_6U_10U_8_IsNaN_6U_10U_8_nor_3_tmp)) | (~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[3])
      | (cfg_precision_1_sva_st_81!=2'b10));
  assign and_3075_nl = (~ IsNaN_6U_10U_9_nor_3_tmp) & FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_5_1
      & FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_4_1 & (FpMul_6U_10U_2_o_expo_lpi_1_dfm_6_3_0_1==4'b1111);
  assign mux_1790_nl = MUX_s_1_2_2((nor_793_nl), (nor_792_nl), and_3075_nl);
  assign nor_795_nl = ~((~ main_stage_v_4) | (chn_inp_in_crt_sva_4_739_736_1[3])
      | (cfg_precision_1_sva_st_81!=2'b10));
  assign mux_1791_nl = MUX_s_1_2_2((nor_795_nl), (mux_1790_nl), nor_956_cse);
  assign nand_780_nl = ~((nor_1130_cse | IsNaN_6U_10U_8_land_lpi_1_dfm_4) & main_stage_v_5);
  assign mux_1792_nl = MUX_s_1_2_2(or_3969_cse, (nand_780_nl), IsNaN_8U_23U_2_land_lpi_1_dfm_9);
  assign mux_1793_nl = MUX_s_1_2_2((mux_1792_nl), or_3716_cse, IsNaN_8U_23U_3_land_lpi_1_dfm_5);
  assign mux_1794_nl = MUX_s_1_2_2(or_3969_cse, (mux_1793_nl), nor_623_cse);
  assign mux_1795_nl = MUX_s_1_2_2((mux_1794_nl), or_3969_cse, IsNaN_6U_10U_9_land_lpi_1_dfm_6);
  assign nor_1954_nl = ~((cfg_precision_1_sva_st_82!=2'b10) | (mux_1795_nl) | (chn_inp_in_crt_sva_5_739_736_1[3]));
  assign mux_1797_nl = MUX_s_1_2_2((nor_1954_nl), (mux_1791_nl), or_11_cse);
  assign nor_791_nl = ~(nor_55_cse | and_348_cse);
  assign mux_1798_nl = MUX_s_1_2_2((nor_791_nl), FpFractionToFloat_35U_6U_10U_is_zero_3_lpi_1_dfm_5,
      chn_inp_in_crt_sva_2_739_736_1[2]);
  assign or_5648_nl = (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10) | (mux_1798_nl);
  assign mux_1799_nl = MUX_s_1_2_2(or_2282_cse, or_tmp_3973, IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_15);
  assign or_3978_nl = (chn_inp_in_crt_sva_3_739_736_1[2]) | (mux_1799_nl);
  assign mux_1800_nl = MUX_s_1_2_2(or_tmp_3973, or_2282_cse, chn_inp_in_crt_sva_3_739_736_1[2]);
  assign mux_1801_nl = MUX_s_1_2_2((mux_1800_nl), (or_3978_nl), IsNaN_6U_10U_5_land_3_lpi_1_dfm_5);
  assign mux_1802_nl = MUX_s_1_2_2((mux_1801_nl), (or_5648_nl), or_11_cse);
  assign mux_1805_nl = MUX_s_1_2_2(nand_tmp_221, nand_tmp_230, or_11_cse);
  assign mux_1808_nl = MUX_s_1_2_2(and_tmp_240, and_152_cse, or_11_cse);
  assign mux_1810_nl = MUX_s_1_2_2(nand_tmp_220, nand_tmp_231, or_11_cse);
  assign mux_1812_nl = MUX_s_1_2_2(and_tmp_242, and_144_cse, or_11_cse);
  assign mux_1814_nl = MUX_s_1_2_2(nand_tmp_219, nand_tmp_232, or_11_cse);
  assign mux_1816_nl = MUX_s_1_2_2(and_tmp_244, and_137_cse, or_11_cse);
  assign mux_1818_nl = MUX_s_1_2_2(nand_tmp_218, nand_tmp_233, or_11_cse);
  assign mux_1820_nl = MUX_s_1_2_2(and_tmp_246, and_131_cse, or_11_cse);
  assign mux_1822_nl = MUX_s_1_2_2(or_5800_cse, nand_tmp_234, or_11_cse);
  assign mux_1823_nl = MUX_s_1_2_2(or_2176_cse, nand_tmp_234, or_11_cse);
  assign mux_1824_nl = MUX_s_1_2_2((mux_1823_nl), (mux_1822_nl), FpFractionToFloat_35U_6U_10U_is_zero_1_lpi_1_dfm_5);
  assign mux_1826_nl = MUX_s_1_2_2(or_tmp_234, nand_tmp_235, or_11_cse);
  assign mux_1827_nl = MUX_s_1_2_2(or_2176_cse, nand_tmp_235, or_11_cse);
  assign mux_1828_nl = MUX_s_1_2_2((mux_1827_nl), (mux_1826_nl), FpFractionToFloat_35U_6U_10U_is_zero_2_lpi_1_dfm_5);
  assign or_4004_nl = (~ main_stage_v_1) | (cfg_precision_1_sva_st_90!=2'b10) | IsNaN_8U_23U_2_land_3_lpi_1_dfm_st_6;
  assign mux_1829_nl = MUX_s_1_2_2(or_tmp_8, (or_4004_nl), chn_inp_in_crt_sva_1_739_395_1[343]);
  assign or_4005_nl = (~ main_stage_v_2) | (cfg_precision_1_sva_st_91!=2'b10) | FpFractionToFloat_35U_6U_10U_is_zero_3_lpi_1_dfm_5;
  assign mux_1830_nl = MUX_s_1_2_2(or_2176_cse, (or_4005_nl), chn_inp_in_crt_sva_2_739_736_1[2]);
  assign mux_1831_nl = MUX_s_1_2_2((mux_1830_nl), (mux_1829_nl), or_11_cse);
  assign inp_lookup_4_IntShiftRight_69U_6U_32U_obits_fixed_and_nl = (reg_chn_inp_in_crt_sva_2_606_576_1_itm[0])
      & inp_lookup_4_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2;
  assign nl_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_1_sva_7 = (reg_chn_inp_in_crt_sva_2_606_576_1_itm[18:1])
      + conv_u2s_1_18(inp_lookup_4_IntShiftRight_69U_6U_32U_obits_fixed_and_nl);
  assign nand_236_nl = ~(main_stage_v_2 & (~(nor_1340_cse | (chn_inp_in_crt_sva_2_739_736_1[3]))));
  assign mux_1833_nl = MUX_s_1_2_2(nand_tmp_230, (nand_236_nl), or_11_cse);
  assign inp_lookup_3_IntShiftRight_69U_6U_32U_obits_fixed_and_nl = (reg_chn_inp_in_crt_sva_2_574_544_1_itm[0])
      & inp_lookup_3_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2;
  assign nl_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_4_sva_7 = (reg_chn_inp_in_crt_sva_2_574_544_1_itm[18:1])
      + conv_u2s_1_18(inp_lookup_3_IntShiftRight_69U_6U_32U_obits_fixed_and_nl);
  assign or_4013_nl = (~ main_stage_v_2) | nor_1340_cse | (chn_inp_in_crt_sva_2_739_736_1[2]);
  assign mux_1835_nl = MUX_s_1_2_2(nand_tmp_231, (or_4013_nl), or_11_cse);
  assign inp_lookup_2_IntShiftRight_69U_6U_32U_obits_fixed_and_nl = (reg_chn_inp_in_crt_sva_2_542_512_1_itm[0])
      & inp_lookup_2_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2;
  assign nl_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_3_sva_7 = (reg_chn_inp_in_crt_sva_2_542_512_1_itm[18:1])
      + conv_u2s_1_18(inp_lookup_2_IntShiftRight_69U_6U_32U_obits_fixed_and_nl);
  assign nand_237_nl = ~(main_stage_v_2 & (~(nor_1340_cse | (chn_inp_in_crt_sva_2_739_736_1[1]))));
  assign mux_1837_nl = MUX_s_1_2_2(nand_tmp_232, (nand_237_nl), or_11_cse);
  assign inp_lookup_1_IntShiftRight_69U_6U_32U_obits_fixed_and_nl = (reg_chn_inp_in_crt_sva_2_510_480_1_itm[0])
      & inp_lookup_1_IntShiftRight_69U_6U_32U_obits_fixed_or_itm_2;
  assign nl_IntShiftRight_69U_6U_32U_obits_fixed_acc_psp_2_sva_7 = (reg_chn_inp_in_crt_sva_2_510_480_1_itm[18:1])
      + conv_u2s_1_18(inp_lookup_1_IntShiftRight_69U_6U_32U_obits_fixed_and_nl);
  assign nand_238_nl = ~(main_stage_v_2 & (~((chn_inp_in_crt_sva_2_739_736_1[0])
      | nor_1340_cse)));
  assign mux_1840_nl = MUX_s_1_2_2(nand_tmp_233, (nand_238_nl), or_11_cse);
  assign inp_lookup_4_IsZero_6U_10U_1_IsZero_6U_10U_1_nor_nl = ~((chn_inp_in_rsci_d_mxwt[458])
      | FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_3_0_mx0w0 | (FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_3_mx0w0!=4'b0000));
  assign inp_lookup_1_IntShiftRight_69U_6U_32U_obits_fixed_or_nl = (inp_lookup_else_else_o_acc_psp_1_sva[0])
      | (inp_lookup_else_else_o_acc_psp_1_sva[1]) | (inp_lookup_else_else_o_acc_psp_1_sva[2])
      | (inp_lookup_else_else_o_acc_psp_1_sva[3]) | (inp_lookup_else_else_o_acc_psp_1_sva[4])
      | (inp_lookup_else_else_o_acc_psp_1_sva[5]) | (inp_lookup_else_else_o_acc_psp_1_sva[6])
      | (inp_lookup_else_else_o_acc_psp_1_sva[7]) | (inp_lookup_else_else_o_acc_psp_1_sva[8])
      | (inp_lookup_else_else_o_acc_psp_1_sva[9]) | (inp_lookup_else_else_o_acc_psp_1_sva[10])
      | (inp_lookup_else_else_o_acc_psp_1_sva[11]) | (inp_lookup_else_else_o_acc_psp_1_sva[12])
      | (inp_lookup_else_else_o_acc_psp_1_sva[13]) | (inp_lookup_else_else_o_acc_psp_1_sva[14])
      | (inp_lookup_else_else_o_acc_psp_1_sva[15]) | (inp_lookup_else_else_o_acc_psp_1_sva[16])
      | (inp_lookup_else_else_o_acc_psp_1_sva[17]) | (inp_lookup_else_else_o_acc_psp_1_sva[18])
      | (inp_lookup_else_else_o_acc_psp_1_sva[19]) | (inp_lookup_else_else_o_acc_psp_1_sva[20])
      | (inp_lookup_else_else_o_acc_psp_1_sva[21]) | (inp_lookup_else_else_o_acc_psp_1_sva[22])
      | (inp_lookup_else_else_o_acc_psp_1_sva[23]) | (inp_lookup_else_else_o_acc_psp_1_sva[24])
      | (inp_lookup_else_else_o_acc_psp_1_sva[25]) | (inp_lookup_else_else_o_acc_psp_1_sva[26])
      | (inp_lookup_else_else_o_acc_psp_1_sva[27]) | (inp_lookup_else_else_o_acc_psp_1_sva[28])
      | (inp_lookup_else_else_o_acc_psp_1_sva[29]) | (inp_lookup_else_else_o_acc_psp_1_sva[30])
      | (inp_lookup_else_else_o_acc_psp_1_sva[31]) | (inp_lookup_else_else_o_acc_psp_1_sva[32])
      | (inp_lookup_else_else_o_acc_psp_1_sva[33]) | (~ (inp_lookup_else_else_o_acc_psp_1_sva[52]));
  assign inp_lookup_1_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_nl = (IntSignedShiftRight_50U_5U_32U_mbits_fixed_1_sva[0])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_1_sva[1]) | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_1_sva[2])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_1_sva[3]) | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_1_sva[4])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_1_sva[5]) | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_1_sva[6])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_1_sva[7]) | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_1_sva[8])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_1_sva[9]) | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_1_sva[10])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_1_sva[11]) | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_1_sva[12])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_1_sva[13]) | (~ (IntSignedShiftRight_50U_5U_32U_mbits_fixed_1_sva[80]));
  assign nor_782_nl = ~(and_3149_cse | ((FpFractionToFloat_35U_6U_10U_1_mux_tmp[4:3]==2'b11)
      & (IntLeadZero_35U_1_leading_sign_35_0_rtn_1_sva_2[5]) & inp_lookup_1_FpMantRNE_36U_11U_1_else_and_svs_2
      & (~ IsNaN_6U_10U_6_nor_tmp) & FpAdd_8U_23U_is_a_greater_lor_1_lpi_1_dfm_1_st_2
      & (FpFractionToFloat_35U_6U_10U_1_mux_tmp[2:0]==3'b111)) | (chn_inp_in_crt_sva_1_739_395_1[341])
      | (~ main_stage_v_1));
  assign mux_1841_nl = MUX_s_1_2_2(nor_tmp_653, (nor_782_nl), cfg_precision_1_sva_st_90[1]);
  assign mux_1842_nl = MUX_s_1_2_2((mux_1841_nl), nor_tmp_653, cfg_precision_1_sva_st_90[0]);
  assign nor_783_nl = ~(IsNaN_6U_10U_7_land_1_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_1_lpi_1_dfm_st_14
      | (chn_inp_in_crt_sva_2_739_736_1[0]) | (~ main_stage_v_2));
  assign mux_1843_nl = MUX_s_1_2_2(nor_tmp_656, (nor_783_nl), cfg_precision_1_sva_st_91[1]);
  assign mux_1844_nl = MUX_s_1_2_2((mux_1843_nl), nor_tmp_656, cfg_precision_1_sva_st_91[0]);
  assign mux_1845_nl = MUX_s_1_2_2((mux_1844_nl), (mux_1842_nl), or_11_cse);
  assign inp_lookup_2_IntShiftRight_69U_6U_32U_obits_fixed_or_nl = (inp_lookup_else_else_o_acc_psp_2_sva[0])
      | (inp_lookup_else_else_o_acc_psp_2_sva[1]) | (inp_lookup_else_else_o_acc_psp_2_sva[2])
      | (inp_lookup_else_else_o_acc_psp_2_sva[3]) | (inp_lookup_else_else_o_acc_psp_2_sva[4])
      | (inp_lookup_else_else_o_acc_psp_2_sva[5]) | (inp_lookup_else_else_o_acc_psp_2_sva[6])
      | (inp_lookup_else_else_o_acc_psp_2_sva[7]) | (inp_lookup_else_else_o_acc_psp_2_sva[8])
      | (inp_lookup_else_else_o_acc_psp_2_sva[9]) | (inp_lookup_else_else_o_acc_psp_2_sva[10])
      | (inp_lookup_else_else_o_acc_psp_2_sva[11]) | (inp_lookup_else_else_o_acc_psp_2_sva[12])
      | (inp_lookup_else_else_o_acc_psp_2_sva[13]) | (inp_lookup_else_else_o_acc_psp_2_sva[14])
      | (inp_lookup_else_else_o_acc_psp_2_sva[15]) | (inp_lookup_else_else_o_acc_psp_2_sva[16])
      | (inp_lookup_else_else_o_acc_psp_2_sva[17]) | (inp_lookup_else_else_o_acc_psp_2_sva[18])
      | (inp_lookup_else_else_o_acc_psp_2_sva[19]) | (inp_lookup_else_else_o_acc_psp_2_sva[20])
      | (inp_lookup_else_else_o_acc_psp_2_sva[21]) | (inp_lookup_else_else_o_acc_psp_2_sva[22])
      | (inp_lookup_else_else_o_acc_psp_2_sva[23]) | (inp_lookup_else_else_o_acc_psp_2_sva[24])
      | (inp_lookup_else_else_o_acc_psp_2_sva[25]) | (inp_lookup_else_else_o_acc_psp_2_sva[26])
      | (inp_lookup_else_else_o_acc_psp_2_sva[27]) | (inp_lookup_else_else_o_acc_psp_2_sva[28])
      | (inp_lookup_else_else_o_acc_psp_2_sva[29]) | (inp_lookup_else_else_o_acc_psp_2_sva[30])
      | (inp_lookup_else_else_o_acc_psp_2_sva[31]) | (inp_lookup_else_else_o_acc_psp_2_sva[32])
      | (inp_lookup_else_else_o_acc_psp_2_sva[33]) | (~ (inp_lookup_else_else_o_acc_psp_2_sva[52]));
  assign inp_lookup_2_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_nl = (IntSignedShiftRight_50U_5U_32U_mbits_fixed_2_sva[0])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_2_sva[1]) | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_2_sva[2])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_2_sva[3]) | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_2_sva[4])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_2_sva[5]) | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_2_sva[6])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_2_sva[7]) | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_2_sva[8])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_2_sva[9]) | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_2_sva[10])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_2_sva[11]) | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_2_sva[12])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_2_sva[13]) | (~ (IntSignedShiftRight_50U_5U_32U_mbits_fixed_2_sva[80]));
  assign nor_776_nl = ~(and_4145_cse | ((FpFractionToFloat_35U_6U_10U_1_mux_40_tmp==5'b11111)
      & (IntLeadZero_35U_1_leading_sign_35_0_rtn_2_sva_2[5]) & inp_lookup_2_FpMantRNE_36U_11U_1_else_and_svs_2
      & (~ IsNaN_6U_10U_6_nor_1_tmp) & FpAdd_8U_23U_is_a_greater_lor_2_lpi_1_dfm_1_st_2)
      | (chn_inp_in_crt_sva_1_739_395_1[342]) | (~ main_stage_v_1));
  assign mux_1846_nl = MUX_s_1_2_2(nor_tmp_657, (nor_776_nl), cfg_precision_1_sva_st_90[1]);
  assign mux_1847_nl = MUX_s_1_2_2((mux_1846_nl), nor_tmp_657, cfg_precision_1_sva_st_90[0]);
  assign nor_777_nl = ~(IsNaN_6U_10U_7_land_2_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_2_lpi_1_dfm_st_14
      | (chn_inp_in_crt_sva_2_739_736_1[1]) | (~ main_stage_v_2));
  assign mux_1848_nl = MUX_s_1_2_2(nor_tmp_660, (nor_777_nl), cfg_precision_1_sva_st_91[1]);
  assign mux_1849_nl = MUX_s_1_2_2((mux_1848_nl), nor_tmp_660, cfg_precision_1_sva_st_91[0]);
  assign mux_1850_nl = MUX_s_1_2_2((mux_1849_nl), (mux_1847_nl), or_11_cse);
  assign inp_lookup_3_IntShiftRight_69U_6U_32U_obits_fixed_or_nl = (inp_lookup_else_else_o_acc_psp_3_sva[0])
      | (inp_lookup_else_else_o_acc_psp_3_sva[1]) | (inp_lookup_else_else_o_acc_psp_3_sva[2])
      | (inp_lookup_else_else_o_acc_psp_3_sva[3]) | (inp_lookup_else_else_o_acc_psp_3_sva[4])
      | (inp_lookup_else_else_o_acc_psp_3_sva[5]) | (inp_lookup_else_else_o_acc_psp_3_sva[6])
      | (inp_lookup_else_else_o_acc_psp_3_sva[7]) | (inp_lookup_else_else_o_acc_psp_3_sva[8])
      | (inp_lookup_else_else_o_acc_psp_3_sva[9]) | (inp_lookup_else_else_o_acc_psp_3_sva[10])
      | (inp_lookup_else_else_o_acc_psp_3_sva[11]) | (inp_lookup_else_else_o_acc_psp_3_sva[12])
      | (inp_lookup_else_else_o_acc_psp_3_sva[13]) | (inp_lookup_else_else_o_acc_psp_3_sva[14])
      | (inp_lookup_else_else_o_acc_psp_3_sva[15]) | (inp_lookup_else_else_o_acc_psp_3_sva[16])
      | (inp_lookup_else_else_o_acc_psp_3_sva[17]) | (inp_lookup_else_else_o_acc_psp_3_sva[18])
      | (inp_lookup_else_else_o_acc_psp_3_sva[19]) | (inp_lookup_else_else_o_acc_psp_3_sva[20])
      | (inp_lookup_else_else_o_acc_psp_3_sva[21]) | (inp_lookup_else_else_o_acc_psp_3_sva[22])
      | (inp_lookup_else_else_o_acc_psp_3_sva[23]) | (inp_lookup_else_else_o_acc_psp_3_sva[24])
      | (inp_lookup_else_else_o_acc_psp_3_sva[25]) | (inp_lookup_else_else_o_acc_psp_3_sva[26])
      | (inp_lookup_else_else_o_acc_psp_3_sva[27]) | (inp_lookup_else_else_o_acc_psp_3_sva[28])
      | (inp_lookup_else_else_o_acc_psp_3_sva[29]) | (inp_lookup_else_else_o_acc_psp_3_sva[30])
      | (inp_lookup_else_else_o_acc_psp_3_sva[31]) | (inp_lookup_else_else_o_acc_psp_3_sva[32])
      | (inp_lookup_else_else_o_acc_psp_3_sva[33]) | (~ (inp_lookup_else_else_o_acc_psp_3_sva[52]));
  assign inp_lookup_3_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_nl = (IntSignedShiftRight_50U_5U_32U_mbits_fixed_3_sva[0])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_3_sva[1]) | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_3_sva[2])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_3_sva[3]) | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_3_sva[4])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_3_sva[5]) | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_3_sva[6])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_3_sva[7]) | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_3_sva[8])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_3_sva[9]) | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_3_sva[10])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_3_sva[11]) | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_3_sva[12])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_3_sva[13]) | (~ (IntSignedShiftRight_50U_5U_32U_mbits_fixed_3_sva[80]));
  assign nor_770_nl = ~(and_3249_cse | ((FpFractionToFloat_35U_6U_10U_1_mux_41_tmp==5'b11111)
      & (IntLeadZero_35U_1_leading_sign_35_0_rtn_3_sva_2[5]) & inp_lookup_3_FpMantRNE_36U_11U_1_else_and_svs_2
      & (~ IsNaN_6U_10U_6_nor_2_tmp) & FpAdd_8U_23U_is_a_greater_lor_3_lpi_1_dfm_1_st_2)
      | (chn_inp_in_crt_sva_1_739_395_1[343]) | (~ main_stage_v_1));
  assign mux_1851_nl = MUX_s_1_2_2(nor_tmp_661, (nor_770_nl), cfg_precision_1_sva_st_90[1]);
  assign mux_1852_nl = MUX_s_1_2_2((mux_1851_nl), nor_tmp_661, cfg_precision_1_sva_st_90[0]);
  assign nor_771_nl = ~(IsNaN_6U_10U_7_land_3_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_3_lpi_1_dfm_st_14
      | (chn_inp_in_crt_sva_2_739_736_1[2]) | (~ main_stage_v_2));
  assign mux_1853_nl = MUX_s_1_2_2(nor_tmp_664, (nor_771_nl), cfg_precision_1_sva_st_91[1]);
  assign mux_1854_nl = MUX_s_1_2_2((mux_1853_nl), nor_tmp_664, cfg_precision_1_sva_st_91[0]);
  assign mux_1855_nl = MUX_s_1_2_2((mux_1854_nl), (mux_1852_nl), or_11_cse);
  assign inp_lookup_4_IntShiftRight_69U_6U_32U_obits_fixed_or_nl = (inp_lookup_else_else_o_acc_psp_sva[0])
      | (inp_lookup_else_else_o_acc_psp_sva[1]) | (inp_lookup_else_else_o_acc_psp_sva[2])
      | (inp_lookup_else_else_o_acc_psp_sva[3]) | (inp_lookup_else_else_o_acc_psp_sva[4])
      | (inp_lookup_else_else_o_acc_psp_sva[5]) | (inp_lookup_else_else_o_acc_psp_sva[6])
      | (inp_lookup_else_else_o_acc_psp_sva[7]) | (inp_lookup_else_else_o_acc_psp_sva[8])
      | (inp_lookup_else_else_o_acc_psp_sva[9]) | (inp_lookup_else_else_o_acc_psp_sva[10])
      | (inp_lookup_else_else_o_acc_psp_sva[11]) | (inp_lookup_else_else_o_acc_psp_sva[12])
      | (inp_lookup_else_else_o_acc_psp_sva[13]) | (inp_lookup_else_else_o_acc_psp_sva[14])
      | (inp_lookup_else_else_o_acc_psp_sva[15]) | (inp_lookup_else_else_o_acc_psp_sva[16])
      | (inp_lookup_else_else_o_acc_psp_sva[17]) | (inp_lookup_else_else_o_acc_psp_sva[18])
      | (inp_lookup_else_else_o_acc_psp_sva[19]) | (inp_lookup_else_else_o_acc_psp_sva[20])
      | (inp_lookup_else_else_o_acc_psp_sva[21]) | (inp_lookup_else_else_o_acc_psp_sva[22])
      | (inp_lookup_else_else_o_acc_psp_sva[23]) | (inp_lookup_else_else_o_acc_psp_sva[24])
      | (inp_lookup_else_else_o_acc_psp_sva[25]) | (inp_lookup_else_else_o_acc_psp_sva[26])
      | (inp_lookup_else_else_o_acc_psp_sva[27]) | (inp_lookup_else_else_o_acc_psp_sva[28])
      | (inp_lookup_else_else_o_acc_psp_sva[29]) | (inp_lookup_else_else_o_acc_psp_sva[30])
      | (inp_lookup_else_else_o_acc_psp_sva[31]) | (inp_lookup_else_else_o_acc_psp_sva[32])
      | (inp_lookup_else_else_o_acc_psp_sva[33]) | (~ (inp_lookup_else_else_o_acc_psp_sva[52]));
  assign inp_lookup_4_IntSignedShiftRight_50U_5U_32U_obits_fixed_or_nl = (IntSignedShiftRight_50U_5U_32U_mbits_fixed_sva[0])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_sva[1]) | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_sva[2])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_sva[3]) | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_sva[4])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_sva[5]) | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_sva[6])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_sva[7]) | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_sva[8])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_sva[9]) | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_sva[10])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_sva[11]) | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_sva[12])
      | (IntSignedShiftRight_50U_5U_32U_mbits_fixed_sva[13]) | (~ (IntSignedShiftRight_50U_5U_32U_mbits_fixed_sva[80]));
  assign nor_764_nl = ~(and_3361_cse_1 | ((FpFractionToFloat_35U_6U_10U_1_mux_42_tmp==5'b11111)
      & (IntLeadZero_35U_1_leading_sign_35_0_rtn_sva_2[5]) & inp_lookup_4_FpMantRNE_36U_11U_1_else_and_svs_2
      & (~ IsNaN_6U_10U_6_nor_3_tmp) & FpAdd_8U_23U_is_a_greater_lor_lpi_1_dfm_1_st_2)
      | (chn_inp_in_crt_sva_1_739_395_1[344]) | (~ main_stage_v_1));
  assign mux_1856_nl = MUX_s_1_2_2(nor_tmp_665, (nor_764_nl), cfg_precision_1_sva_st_90[1]);
  assign mux_1857_nl = MUX_s_1_2_2((mux_1856_nl), nor_tmp_665, cfg_precision_1_sva_st_90[0]);
  assign nor_765_nl = ~(IsNaN_6U_10U_7_land_lpi_1_dfm_5 | IsNaN_6U_10U_2_land_lpi_1_dfm_st_14
      | (chn_inp_in_crt_sva_2_739_736_1[3]) | (~ main_stage_v_2));
  assign mux_1858_nl = MUX_s_1_2_2(nor_tmp_668, (nor_765_nl), cfg_precision_1_sva_st_91[1]);
  assign mux_1859_nl = MUX_s_1_2_2((mux_1858_nl), nor_tmp_668, cfg_precision_1_sva_st_91[0]);
  assign mux_1860_nl = MUX_s_1_2_2((mux_1859_nl), (mux_1857_nl), or_11_cse);
  assign nl_inp_lookup_1_else_else_b1_mul_itm_2 = $signed((chn_inp_in_rsci_d_mxwt[347:332]))
      * $signed(conv_u2s_35_36(chn_inp_in_rsci_d_mxwt[162:128]));
  assign nor_761_nl = ~((chn_inp_in_rsci_d_mxwt[736]) | (~ and_dcpl_42));
  assign nor_762_nl = ~((~ main_stage_v_1) | (chn_inp_in_crt_sva_1_739_395_1[341])
      | nor_1336_cse_1);
  assign mux_1861_nl = MUX_s_1_2_2((nor_762_nl), (nor_761_nl), or_11_cse);
  assign nl_inp_lookup_2_else_else_b1_mul_itm_2 = $signed((chn_inp_in_rsci_d_mxwt[363:348]))
      * $signed(conv_u2s_35_36(chn_inp_in_rsci_d_mxwt[197:163]));
  assign nor_759_nl = ~((chn_inp_in_rsci_d_mxwt[737]) | (~ and_dcpl_42));
  assign nor_760_nl = ~((~ main_stage_v_1) | (chn_inp_in_crt_sva_1_739_395_1[342])
      | nor_1336_cse_1);
  assign mux_1862_nl = MUX_s_1_2_2((nor_760_nl), (nor_759_nl), or_11_cse);
  assign nl_inp_lookup_3_else_else_b1_mul_itm_2 = $signed((chn_inp_in_rsci_d_mxwt[379:364]))
      * $signed(conv_u2s_35_36(chn_inp_in_rsci_d_mxwt[232:198]));
  assign nor_757_nl = ~((chn_inp_in_rsci_d_mxwt[738]) | (~ and_dcpl_42));
  assign and_3058_nl = (~((chn_inp_in_crt_sva_1_739_395_1[343]) | (~ main_stage_v_1)))
      & nor_758_cse;
  assign mux_1863_nl = MUX_s_1_2_2((and_3058_nl), (nor_757_nl), or_11_cse);
  assign nl_inp_lookup_4_else_else_b1_mul_itm_2 = $signed((chn_inp_in_rsci_d_mxwt[395:380]))
      * $signed(conv_u2s_35_36(chn_inp_in_rsci_d_mxwt[267:233]));
  assign nor_755_nl = ~((chn_inp_in_rsci_d_mxwt[739]) | (~ and_dcpl_42));
  assign and_nl = (~((chn_inp_in_crt_sva_1_739_395_1[344]) | (~ main_stage_v_1)))
      & nor_756_cse;
  assign mux_1864_nl = MUX_s_1_2_2((and_nl), (nor_755_nl), or_11_cse);
  assign and_4121_nl = (inp_lookup_4_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[35:24]==12'b111111111111);
  assign mux_2130_nl = MUX_s_1_2_2((and_4121_nl), inp_lookup_4_FpMantRNE_36U_11U_1_else_and_svs,
      not_tmp_69);
  assign and_4120_nl = (inp_lookup_3_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[35:24]==12'b111111111111);
  assign mux_2131_nl = MUX_s_1_2_2(inp_lookup_3_FpMantRNE_36U_11U_1_else_and_svs,
      (and_4120_nl), or_79_cse);
  assign and_4119_nl = (inp_lookup_2_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[35:24]==12'b111111111111);
  assign mux_2132_nl = MUX_s_1_2_2((and_4119_nl), inp_lookup_2_FpMantRNE_36U_11U_1_else_and_svs,
      not_tmp_45);
  assign and_4118_nl = (inp_lookup_1_FpFractionToFloat_35U_6U_10U_1_if_shifted_frac_p1_lshift_tmp[35:24]==12'b111111111111);
  assign mux_2133_nl = MUX_s_1_2_2((and_4118_nl), inp_lookup_1_FpMantRNE_36U_11U_1_else_and_svs,
      not_tmp_34);
  assign FpAdd_8U_23U_if_2_mux_8_nl = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_qr_1_lpi_1_dfm_4,
      (~ FpAdd_8U_23U_addend_smaller_qr_1_lpi_1_dfm_4), FpAdd_8U_23U_else_2_and_tmp);
  assign FpAdd_8U_23U_if_2_FpAdd_8U_23U_if_2_nand_4_nl = ~((fsm_output[1]) & inp_lookup_1_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_4);
  assign FpAdd_8U_23U_if_2_mux_9_nl = MUX_v_49_2_2(FpAdd_8U_23U_addend_smaller_qr_1_lpi_1_dfm_4,
      FpAdd_8U_23U_addend_larger_qr_1_lpi_1_dfm_4, FpAdd_8U_23U_else_2_and_tmp);
  assign nl_acc_nl = ({FpAdd_8U_23U_else_2_and_tmp , (FpAdd_8U_23U_if_2_mux_8_nl)
      , (FpAdd_8U_23U_if_2_FpAdd_8U_23U_if_2_nand_4_nl)}) + conv_u2u_50_51({(FpAdd_8U_23U_if_2_mux_9_nl)
      , 1'b1});
  assign acc_nl = nl_acc_nl[50:0];
  assign z_out = readslicef_51_50_1((acc_nl));
  assign FpAdd_8U_23U_if_2_mux_10_nl = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_qr_2_lpi_1_dfm_4,
      (~ FpAdd_8U_23U_addend_smaller_qr_2_lpi_1_dfm_4), FpAdd_8U_23U_else_2_and_tmp_1);
  assign FpAdd_8U_23U_if_2_FpAdd_8U_23U_if_2_nand_5_nl = ~((fsm_output[1]) & inp_lookup_2_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_4);
  assign FpAdd_8U_23U_if_2_mux_11_nl = MUX_v_49_2_2(FpAdd_8U_23U_addend_smaller_qr_2_lpi_1_dfm_4,
      FpAdd_8U_23U_addend_larger_qr_2_lpi_1_dfm_4, FpAdd_8U_23U_else_2_and_tmp_1);
  assign nl_acc_1_nl = ({FpAdd_8U_23U_else_2_and_tmp_1 , (FpAdd_8U_23U_if_2_mux_10_nl)
      , (FpAdd_8U_23U_if_2_FpAdd_8U_23U_if_2_nand_5_nl)}) + conv_u2u_50_51({(FpAdd_8U_23U_if_2_mux_11_nl)
      , 1'b1});
  assign acc_1_nl = nl_acc_1_nl[50:0];
  assign z_out_1 = readslicef_51_50_1((acc_1_nl));
  assign FpAdd_8U_23U_if_2_mux_12_nl = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_qr_3_lpi_1_dfm_4,
      (~ FpAdd_8U_23U_addend_smaller_qr_3_lpi_1_dfm_4), FpAdd_8U_23U_else_2_and_tmp_2);
  assign FpAdd_8U_23U_if_2_FpAdd_8U_23U_if_2_nand_6_nl = ~((fsm_output[1]) & inp_lookup_3_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_4);
  assign FpAdd_8U_23U_if_2_mux_13_nl = MUX_v_49_2_2(FpAdd_8U_23U_addend_smaller_qr_3_lpi_1_dfm_4,
      FpAdd_8U_23U_addend_larger_qr_3_lpi_1_dfm_4, FpAdd_8U_23U_else_2_and_tmp_2);
  assign nl_acc_2_nl = ({FpAdd_8U_23U_else_2_and_tmp_2 , (FpAdd_8U_23U_if_2_mux_12_nl)
      , (FpAdd_8U_23U_if_2_FpAdd_8U_23U_if_2_nand_6_nl)}) + conv_u2u_50_51({(FpAdd_8U_23U_if_2_mux_13_nl)
      , 1'b1});
  assign acc_2_nl = nl_acc_2_nl[50:0];
  assign z_out_2 = readslicef_51_50_1((acc_2_nl));
  assign FpAdd_8U_23U_if_2_mux_14_nl = MUX_v_49_2_2(FpAdd_8U_23U_addend_larger_qr_lpi_1_dfm_4,
      (~ FpAdd_8U_23U_addend_smaller_qr_lpi_1_dfm_4), FpAdd_8U_23U_else_2_and_tmp_3);
  assign FpAdd_8U_23U_if_2_FpAdd_8U_23U_if_2_nand_7_nl = ~((fsm_output[1]) & inp_lookup_4_FpAdd_8U_23U_is_addition_FpAdd_8U_23U_is_addition_xnor_svs_4);
  assign FpAdd_8U_23U_if_2_mux_15_nl = MUX_v_49_2_2(FpAdd_8U_23U_addend_smaller_qr_lpi_1_dfm_4,
      FpAdd_8U_23U_addend_larger_qr_lpi_1_dfm_4, FpAdd_8U_23U_else_2_and_tmp_3);
  assign nl_acc_3_nl = ({FpAdd_8U_23U_else_2_and_tmp_3 , (FpAdd_8U_23U_if_2_mux_14_nl)
      , (FpAdd_8U_23U_if_2_FpAdd_8U_23U_if_2_nand_7_nl)}) + conv_u2u_50_51({(FpAdd_8U_23U_if_2_mux_15_nl)
      , 1'b1});
  assign acc_3_nl = nl_acc_3_nl[50:0];
  assign z_out_3 = readslicef_51_50_1((acc_3_nl));
  assign FpAdd_8U_23U_b_right_shift_qif_mux_8_nl = MUX_v_8_2_2((chn_inp_in_crt_sva_1_739_395_1[115:108]),
      (chn_inp_in_crt_sva_1_739_395_1[243:236]), FpAdd_8U_23U_a_right_shift_qelse_and_tmp);
  assign FpAdd_8U_23U_b_right_shift_qif_mux_9_nl = MUX_v_8_2_2((~ (chn_inp_in_crt_sva_1_739_395_1[243:236])),
      (~ (chn_inp_in_crt_sva_1_739_395_1[115:108])), FpAdd_8U_23U_a_right_shift_qelse_and_tmp);
  assign nl_acc_4_nl = ({(FpAdd_8U_23U_b_right_shift_qif_mux_8_nl) , 1'b1}) + ({(FpAdd_8U_23U_b_right_shift_qif_mux_9_nl)
      , 1'b1});
  assign acc_4_nl = nl_acc_4_nl[8:0];
  assign z_out_4 = readslicef_9_8_1((acc_4_nl));
  assign FpAdd_8U_23U_b_right_shift_qif_mux_10_nl = MUX_v_8_2_2((chn_inp_in_crt_sva_1_739_395_1[211:204]),
      (chn_inp_in_crt_sva_1_739_395_1[339:332]), FpAdd_8U_23U_a_right_shift_qelse_and_tmp_1);
  assign FpAdd_8U_23U_b_right_shift_qif_mux_11_nl = MUX_v_8_2_2((~ (chn_inp_in_crt_sva_1_739_395_1[339:332])),
      (~ (chn_inp_in_crt_sva_1_739_395_1[211:204])), FpAdd_8U_23U_a_right_shift_qelse_and_tmp_1);
  assign nl_acc_5_nl = ({(FpAdd_8U_23U_b_right_shift_qif_mux_10_nl) , 1'b1}) + ({(FpAdd_8U_23U_b_right_shift_qif_mux_11_nl)
      , 1'b1});
  assign acc_5_nl = nl_acc_5_nl[8:0];
  assign z_out_5 = readslicef_9_8_1((acc_5_nl));
  assign FpAdd_8U_23U_b_right_shift_qif_mux_12_nl = MUX_v_8_2_2((chn_inp_in_crt_sva_1_739_395_1[147:140]),
      (chn_inp_in_crt_sva_1_739_395_1[275:268]), FpAdd_8U_23U_a_right_shift_qelse_and_tmp_2);
  assign FpAdd_8U_23U_b_right_shift_qif_mux_13_nl = MUX_v_8_2_2((~ (chn_inp_in_crt_sva_1_739_395_1[275:268])),
      (~ (chn_inp_in_crt_sva_1_739_395_1[147:140])), FpAdd_8U_23U_a_right_shift_qelse_and_tmp_2);
  assign nl_acc_6_nl = ({(FpAdd_8U_23U_b_right_shift_qif_mux_12_nl) , 1'b1}) + ({(FpAdd_8U_23U_b_right_shift_qif_mux_13_nl)
      , 1'b1});
  assign acc_6_nl = nl_acc_6_nl[8:0];
  assign z_out_6 = readslicef_9_8_1((acc_6_nl));
  assign FpAdd_8U_23U_b_right_shift_qif_mux_14_nl = MUX_v_8_2_2((chn_inp_in_crt_sva_1_739_395_1[179:172]),
      (chn_inp_in_crt_sva_1_739_395_1[307:300]), FpAdd_8U_23U_a_right_shift_qelse_and_tmp_3);
  assign FpAdd_8U_23U_b_right_shift_qif_mux_15_nl = MUX_v_8_2_2((~ (chn_inp_in_crt_sva_1_739_395_1[307:300])),
      (~ (chn_inp_in_crt_sva_1_739_395_1[179:172])), FpAdd_8U_23U_a_right_shift_qelse_and_tmp_3);
  assign nl_acc_7_nl = ({(FpAdd_8U_23U_b_right_shift_qif_mux_14_nl) , 1'b1}) + ({(FpAdd_8U_23U_b_right_shift_qif_mux_15_nl)
      , 1'b1});
  assign acc_7_nl = nl_acc_7_nl[8:0];
  assign z_out_7 = readslicef_9_8_1((acc_7_nl));
  assign FpMul_6U_10U_oelse_1_FpMul_6U_10U_oelse_1_or_4_nl = FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_12_1_1
      | FpAdd_6U_10U_1_if_4_if_and_tmp;
  assign FpMul_6U_10U_oelse_1_mux_28_nl = MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_1_lpi_1_dfm_12_0_1,
      FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_5, FpAdd_6U_10U_1_if_4_if_and_tmp);
  assign FpMul_6U_10U_oelse_1_mux_29_nl = MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_1_lpi_1_dfm_21,
      ({FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_4 , (FpAdd_6U_10U_1_o_expo_1_lpi_1_dfm_2_3_0[3:1])}),
      FpAdd_6U_10U_1_if_4_if_and_tmp);
  assign nl_z_out_8 = conv_u2u_6_7({(FpMul_6U_10U_oelse_1_FpMul_6U_10U_oelse_1_or_4_nl)
      , (FpMul_6U_10U_oelse_1_mux_28_nl) , (FpMul_6U_10U_oelse_1_mux_29_nl)}) + conv_s2u_6_7({(~
      FpAdd_6U_10U_1_if_4_if_and_tmp) , 5'b1});
  assign z_out_8 = nl_z_out_8[6:0];
  assign FpMul_6U_10U_oelse_1_FpMul_6U_10U_oelse_1_or_5_nl = FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_12_1_1
      | FpAdd_6U_10U_1_if_4_if_and_tmp_1;
  assign FpMul_6U_10U_oelse_1_mux_30_nl = MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_2_lpi_1_dfm_12_0_1,
      FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_5, FpAdd_6U_10U_1_if_4_if_and_tmp_1);
  assign FpMul_6U_10U_oelse_1_mux_31_nl = MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_2_lpi_1_dfm_21,
      ({FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_4 , (FpAdd_6U_10U_1_o_expo_2_lpi_1_dfm_2_3_0[3:1])}),
      FpAdd_6U_10U_1_if_4_if_and_tmp_1);
  assign nl_z_out_9 = conv_u2u_6_7({(FpMul_6U_10U_oelse_1_FpMul_6U_10U_oelse_1_or_5_nl)
      , (FpMul_6U_10U_oelse_1_mux_30_nl) , (FpMul_6U_10U_oelse_1_mux_31_nl)}) + conv_s2u_6_7({(~
      FpAdd_6U_10U_1_if_4_if_and_tmp_1) , 5'b1});
  assign z_out_9 = nl_z_out_9[6:0];
  assign FpMul_6U_10U_oelse_1_FpMul_6U_10U_oelse_1_or_6_nl = FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_12_1_1
      | FpAdd_6U_10U_1_if_4_if_and_tmp_2;
  assign FpMul_6U_10U_oelse_1_mux_32_nl = MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_3_lpi_1_dfm_12_0_1,
      FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_5, FpAdd_6U_10U_1_if_4_if_and_tmp_2);
  assign FpMul_6U_10U_oelse_1_mux_33_nl = MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_3_lpi_1_dfm_21,
      ({FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_4 , (FpAdd_6U_10U_1_o_expo_3_lpi_1_dfm_2_3_0[3:1])}),
      FpAdd_6U_10U_1_if_4_if_and_tmp_2);
  assign nl_z_out_10 = conv_u2u_6_7({(FpMul_6U_10U_oelse_1_FpMul_6U_10U_oelse_1_or_6_nl)
      , (FpMul_6U_10U_oelse_1_mux_32_nl) , (FpMul_6U_10U_oelse_1_mux_33_nl)}) + conv_s2u_6_7({(~
      FpAdd_6U_10U_1_if_4_if_and_tmp_2) , 5'b1});
  assign z_out_10 = nl_z_out_10[6:0];
  assign FpMul_6U_10U_oelse_1_FpMul_6U_10U_oelse_1_or_7_nl = FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_12_1_1
      | FpAdd_6U_10U_1_if_4_if_and_tmp_3;
  assign FpMul_6U_10U_oelse_1_mux_34_nl = MUX_s_1_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_5_4_lpi_1_dfm_12_0_1,
      FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_5, FpAdd_6U_10U_1_if_4_if_and_tmp_3);
  assign FpMul_6U_10U_oelse_1_mux_35_nl = MUX_v_4_2_2(FpExpoWidthInc_5U_6U_10U_1U_1U_o_expo_3_0_lpi_1_dfm_21,
      ({FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_4 , (FpAdd_6U_10U_1_o_expo_lpi_1_dfm_2_3_0[3:1])}),
      FpAdd_6U_10U_1_if_4_if_and_tmp_3);
  assign nl_z_out_11 = conv_u2u_6_7({(FpMul_6U_10U_oelse_1_FpMul_6U_10U_oelse_1_or_7_nl)
      , (FpMul_6U_10U_oelse_1_mux_34_nl) , (FpMul_6U_10U_oelse_1_mux_35_nl)}) + conv_s2u_6_7({(~
      FpAdd_6U_10U_1_if_4_if_and_tmp_3) , 5'b1});
  assign z_out_11 = nl_z_out_11[6:0];
  assign FpAdd_6U_10U_a_right_shift_qelse_mux_24_nl = MUX_s_1_2_2(reg_FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_5_4_tmp,
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_15_tmp, FpAdd_6U_10U_b_right_shift_qif_and_tmp);
  assign FpAdd_6U_10U_a_right_shift_qelse_mux_25_nl = MUX_s_1_2_2(reg_FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_5_4_tmp_1,
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_15_tmp_1, FpAdd_6U_10U_b_right_shift_qif_and_tmp);
  assign FpAdd_6U_10U_a_right_shift_qelse_mux_26_nl = MUX_v_4_2_2(FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_3_0_1,
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_27, FpAdd_6U_10U_b_right_shift_qif_and_tmp);
  assign FpAdd_6U_10U_a_right_shift_qelse_mux_27_nl = MUX_s_1_2_2((~ reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_15_tmp),
      (~ reg_FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_5_4_tmp), FpAdd_6U_10U_b_right_shift_qif_and_tmp);
  assign FpAdd_6U_10U_a_right_shift_qelse_mux_28_nl = MUX_s_1_2_2((~ reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_1_lpi_1_dfm_15_tmp_1),
      (~ reg_FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_5_4_tmp_1), FpAdd_6U_10U_b_right_shift_qif_and_tmp);
  assign FpAdd_6U_10U_a_right_shift_qelse_mux_29_nl = MUX_v_4_2_2((~ FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_1_lpi_1_dfm_27),
      (~ FpMul_6U_10U_o_expo_1_lpi_1_dfm_6_3_0_1), FpAdd_6U_10U_b_right_shift_qif_and_tmp);
  assign nl_acc_12_nl = ({(FpAdd_6U_10U_a_right_shift_qelse_mux_24_nl) , (FpAdd_6U_10U_a_right_shift_qelse_mux_25_nl)
      , (FpAdd_6U_10U_a_right_shift_qelse_mux_26_nl) , 1'b1}) + ({(FpAdd_6U_10U_a_right_shift_qelse_mux_27_nl)
      , (FpAdd_6U_10U_a_right_shift_qelse_mux_28_nl) , (FpAdd_6U_10U_a_right_shift_qelse_mux_29_nl)
      , 1'b1});
  assign acc_12_nl = nl_acc_12_nl[6:0];
  assign z_out_12 = readslicef_7_6_1((acc_12_nl));
  assign FpAdd_6U_10U_a_right_shift_qelse_mux_30_nl = MUX_s_1_2_2(reg_FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_5_4_tmp,
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_15_tmp, FpAdd_6U_10U_b_right_shift_qif_and_tmp_1);
  assign FpAdd_6U_10U_a_right_shift_qelse_mux_31_nl = MUX_s_1_2_2(reg_FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_5_4_tmp_1,
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_15_tmp_1, FpAdd_6U_10U_b_right_shift_qif_and_tmp_1);
  assign FpAdd_6U_10U_a_right_shift_qelse_mux_32_nl = MUX_v_4_2_2(FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_3_0_1,
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_27, FpAdd_6U_10U_b_right_shift_qif_and_tmp_1);
  assign FpAdd_6U_10U_a_right_shift_qelse_mux_33_nl = MUX_s_1_2_2((~ reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_15_tmp),
      (~ reg_FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_5_4_tmp), FpAdd_6U_10U_b_right_shift_qif_and_tmp_1);
  assign FpAdd_6U_10U_a_right_shift_qelse_mux_34_nl = MUX_s_1_2_2((~ reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_2_lpi_1_dfm_15_tmp_1),
      (~ reg_FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_5_4_tmp_1), FpAdd_6U_10U_b_right_shift_qif_and_tmp_1);
  assign FpAdd_6U_10U_a_right_shift_qelse_mux_35_nl = MUX_v_4_2_2((~ FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_2_lpi_1_dfm_27),
      (~ FpMul_6U_10U_o_expo_2_lpi_1_dfm_6_3_0_1), FpAdd_6U_10U_b_right_shift_qif_and_tmp_1);
  assign nl_acc_13_nl = ({(FpAdd_6U_10U_a_right_shift_qelse_mux_30_nl) , (FpAdd_6U_10U_a_right_shift_qelse_mux_31_nl)
      , (FpAdd_6U_10U_a_right_shift_qelse_mux_32_nl) , 1'b1}) + ({(FpAdd_6U_10U_a_right_shift_qelse_mux_33_nl)
      , (FpAdd_6U_10U_a_right_shift_qelse_mux_34_nl) , (FpAdd_6U_10U_a_right_shift_qelse_mux_35_nl)
      , 1'b1});
  assign acc_13_nl = nl_acc_13_nl[6:0];
  assign z_out_13 = readslicef_7_6_1((acc_13_nl));
  assign FpAdd_6U_10U_a_right_shift_qelse_mux_36_nl = MUX_s_1_2_2(reg_FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_5_4_tmp,
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_15_tmp, FpAdd_6U_10U_b_right_shift_qif_and_tmp_2);
  assign FpAdd_6U_10U_a_right_shift_qelse_mux_37_nl = MUX_s_1_2_2(reg_FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_5_4_tmp_1,
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_15_tmp_1, FpAdd_6U_10U_b_right_shift_qif_and_tmp_2);
  assign FpAdd_6U_10U_a_right_shift_qelse_mux_38_nl = MUX_v_4_2_2(FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_3_0_1,
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_27, FpAdd_6U_10U_b_right_shift_qif_and_tmp_2);
  assign FpAdd_6U_10U_a_right_shift_qelse_mux_39_nl = MUX_s_1_2_2((~ reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_15_tmp),
      (~ reg_FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_5_4_tmp), FpAdd_6U_10U_b_right_shift_qif_and_tmp_2);
  assign FpAdd_6U_10U_a_right_shift_qelse_mux_40_nl = MUX_s_1_2_2((~ reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_3_lpi_1_dfm_15_tmp_1),
      (~ reg_FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_5_4_tmp_1), FpAdd_6U_10U_b_right_shift_qif_and_tmp_2);
  assign FpAdd_6U_10U_a_right_shift_qelse_mux_41_nl = MUX_v_4_2_2((~ FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_3_lpi_1_dfm_27),
      (~ FpMul_6U_10U_o_expo_3_lpi_1_dfm_6_3_0_1), FpAdd_6U_10U_b_right_shift_qif_and_tmp_2);
  assign nl_acc_14_nl = ({(FpAdd_6U_10U_a_right_shift_qelse_mux_36_nl) , (FpAdd_6U_10U_a_right_shift_qelse_mux_37_nl)
      , (FpAdd_6U_10U_a_right_shift_qelse_mux_38_nl) , 1'b1}) + ({(FpAdd_6U_10U_a_right_shift_qelse_mux_39_nl)
      , (FpAdd_6U_10U_a_right_shift_qelse_mux_40_nl) , (FpAdd_6U_10U_a_right_shift_qelse_mux_41_nl)
      , 1'b1});
  assign acc_14_nl = nl_acc_14_nl[6:0];
  assign z_out_14 = readslicef_7_6_1((acc_14_nl));
  assign FpAdd_6U_10U_a_right_shift_qelse_mux_42_nl = MUX_s_1_2_2(reg_FpMul_6U_10U_o_expo_lpi_1_dfm_6_5_4_tmp,
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_15_tmp, FpAdd_6U_10U_b_right_shift_qif_and_tmp_3);
  assign FpAdd_6U_10U_a_right_shift_qelse_mux_43_nl = MUX_s_1_2_2(reg_FpMul_6U_10U_o_expo_lpi_1_dfm_6_5_4_tmp_1,
      reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_15_tmp_1, FpAdd_6U_10U_b_right_shift_qif_and_tmp_3);
  assign FpAdd_6U_10U_a_right_shift_qelse_mux_44_nl = MUX_v_4_2_2(FpMul_6U_10U_o_expo_lpi_1_dfm_6_3_0_1,
      FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_27, FpAdd_6U_10U_b_right_shift_qif_and_tmp_3);
  assign FpAdd_6U_10U_a_right_shift_qelse_mux_45_nl = MUX_s_1_2_2((~ reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_15_tmp),
      (~ reg_FpMul_6U_10U_o_expo_lpi_1_dfm_6_5_4_tmp), FpAdd_6U_10U_b_right_shift_qif_and_tmp_3);
  assign FpAdd_6U_10U_a_right_shift_qelse_mux_46_nl = MUX_s_1_2_2((~ reg_FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_5_4_lpi_1_dfm_15_tmp_1),
      (~ reg_FpMul_6U_10U_o_expo_lpi_1_dfm_6_5_4_tmp_1), FpAdd_6U_10U_b_right_shift_qif_and_tmp_3);
  assign FpAdd_6U_10U_a_right_shift_qelse_mux_47_nl = MUX_v_4_2_2((~ FpExpoWidthInc_5U_6U_10U_1U_1U_1_o_expo_3_0_lpi_1_dfm_27),
      (~ FpMul_6U_10U_o_expo_lpi_1_dfm_6_3_0_1), FpAdd_6U_10U_b_right_shift_qif_and_tmp_3);
  assign nl_acc_15_nl = ({(FpAdd_6U_10U_a_right_shift_qelse_mux_42_nl) , (FpAdd_6U_10U_a_right_shift_qelse_mux_43_nl)
      , (FpAdd_6U_10U_a_right_shift_qelse_mux_44_nl) , 1'b1}) + ({(FpAdd_6U_10U_a_right_shift_qelse_mux_45_nl)
      , (FpAdd_6U_10U_a_right_shift_qelse_mux_46_nl) , (FpAdd_6U_10U_a_right_shift_qelse_mux_47_nl)
      , 1'b1});
  assign acc_15_nl = nl_acc_15_nl[6:0];
  assign z_out_15 = readslicef_7_6_1((acc_15_nl));
  function [0:0] MUX1HOT_s_1_1_2;
    input [0:0] input_0;
    input [0:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    MUX1HOT_s_1_1_2 = result;
  end
  endfunction
  function [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction
  function [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction
  function [9:0] MUX1HOT_v_10_3_2;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [2:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | ( input_1 & {10{sel[1]}});
    result = result | ( input_2 & {10{sel[2]}});
    MUX1HOT_v_10_3_2 = result;
  end
  endfunction
  function [9:0] MUX1HOT_v_10_4_2;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [3:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | ( input_1 & {10{sel[1]}});
    result = result | ( input_2 & {10{sel[2]}});
    result = result | ( input_3 & {10{sel[3]}});
    MUX1HOT_v_10_4_2 = result;
  end
  endfunction
  function [9:0] MUX1HOT_v_10_5_2;
    input [9:0] input_4;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [4:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | ( input_1 & {10{sel[1]}});
    result = result | ( input_2 & {10{sel[2]}});
    result = result | ( input_3 & {10{sel[3]}});
    result = result | ( input_4 & {10{sel[4]}});
    MUX1HOT_v_10_5_2 = result;
  end
  endfunction
  function [22:0] MUX1HOT_v_23_3_2;
    input [22:0] input_2;
    input [22:0] input_1;
    input [22:0] input_0;
    input [2:0] sel;
    reg [22:0] result;
  begin
    result = input_0 & {23{sel[0]}};
    result = result | ( input_1 & {23{sel[1]}});
    result = result | ( input_2 & {23{sel[2]}});
    MUX1HOT_v_23_3_2 = result;
  end
  endfunction
  function [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction
  function [30:0] MUX1HOT_v_31_3_2;
    input [30:0] input_2;
    input [30:0] input_1;
    input [30:0] input_0;
    input [2:0] sel;
    reg [30:0] result;
  begin
    result = input_0 & {31{sel[0]}};
    result = result | ( input_1 & {31{sel[1]}});
    result = result | ( input_2 & {31{sel[2]}});
    MUX1HOT_v_31_3_2 = result;
  end
  endfunction
  function [31:0] MUX1HOT_v_32_3_2;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [2:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    MUX1HOT_v_32_3_2 = result;
  end
  endfunction
  function [35:0] MUX1HOT_v_36_3_2;
    input [35:0] input_2;
    input [35:0] input_1;
    input [35:0] input_0;
    input [2:0] sel;
    reg [35:0] result;
  begin
    result = input_0 & {36{sel[0]}};
    result = result | ( input_1 & {36{sel[1]}});
    result = result | ( input_2 & {36{sel[2]}});
    MUX1HOT_v_36_3_2 = result;
  end
  endfunction
  function [2:0] MUX1HOT_v_3_4_2;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [3:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    result = result | ( input_3 & {3{sel[3]}});
    MUX1HOT_v_3_4_2 = result;
  end
  endfunction
  function [3:0] MUX1HOT_v_4_3_2;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [2:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    MUX1HOT_v_4_3_2 = result;
  end
  endfunction
  function [3:0] MUX1HOT_v_4_4_2;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [3:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    result = result | ( input_3 & {4{sel[3]}});
    MUX1HOT_v_4_4_2 = result;
  end
  endfunction
  function [4:0] MUX1HOT_v_5_4_2;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [3:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | ( input_1 & {5{sel[1]}});
    result = result | ( input_2 & {5{sel[2]}});
    result = result | ( input_3 & {5{sel[3]}});
    MUX1HOT_v_5_4_2 = result;
  end
  endfunction
  function [5:0] MUX1HOT_v_6_3_2;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [2:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | ( input_1 & {6{sel[1]}});
    result = result | ( input_2 & {6{sel[2]}});
    MUX1HOT_v_6_3_2 = result;
  end
  endfunction
  function [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction
  function [7:0] MUX1HOT_v_8_4_2;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [3:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    result = result | ( input_3 & {8{sel[3]}});
    MUX1HOT_v_8_4_2 = result;
  end
  endfunction
  function [8:0] MUX1HOT_v_9_3_2;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [2:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | ( input_1 & {9{sel[1]}});
    result = result | ( input_2 & {9{sel[2]}});
    MUX1HOT_v_9_3_2 = result;
  end
  endfunction
  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction
  function [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction
  function [16:0] MUX_v_17_2_2;
    input [16:0] input_0;
    input [16:0] input_1;
    input [0:0] sel;
    reg [16:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_17_2_2 = result;
  end
  endfunction
  function [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input [0:0] sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction
  function [20:0] MUX_v_21_2_2;
    input [20:0] input_0;
    input [20:0] input_1;
    input [0:0] sel;
    reg [20:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_21_2_2 = result;
  end
  endfunction
  function [21:0] MUX_v_22_2_2;
    input [21:0] input_0;
    input [21:0] input_1;
    input [0:0] sel;
    reg [21:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_22_2_2 = result;
  end
  endfunction
  function [22:0] MUX_v_23_2_2;
    input [22:0] input_0;
    input [22:0] input_1;
    input [0:0] sel;
    reg [22:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_23_2_2 = result;
  end
  endfunction
  function [23:0] MUX_v_24_2_2;
    input [23:0] input_0;
    input [23:0] input_1;
    input [0:0] sel;
    reg [23:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_24_2_2 = result;
  end
  endfunction
  function [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction
  function [29:0] MUX_v_30_2_2;
    input [29:0] input_0;
    input [29:0] input_1;
    input [0:0] sel;
    reg [29:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_30_2_2 = result;
  end
  endfunction
  function [30:0] MUX_v_31_2_2;
    input [30:0] input_0;
    input [30:0] input_1;
    input [0:0] sel;
    reg [30:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_31_2_2 = result;
  end
  endfunction
  function [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction
  function [48:0] MUX_v_49_2_2;
    input [48:0] input_0;
    input [48:0] input_1;
    input [0:0] sel;
    reg [48:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_49_2_2 = result;
  end
  endfunction
  function [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction
  function [49:0] MUX_v_50_2_2;
    input [49:0] input_0;
    input [49:0] input_1;
    input [0:0] sel;
    reg [49:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_50_2_2 = result;
  end
  endfunction
  function [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction
  function [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction
  function [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction
  function [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [0:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction
  function [0:0] readslicef_11_1_10;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_11_1_10 = tmp[0:0];
  end
  endfunction
  function [0:0] readslicef_24_1_23;
    input [23:0] vector;
    reg [23:0] tmp;
  begin
    tmp = vector >> 23;
    readslicef_24_1_23 = tmp[0:0];
  end
  endfunction
  function [0:0] readslicef_3_1_2;
    input [2:0] vector;
    reg [2:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_3_1_2 = tmp[0:0];
  end
  endfunction
  function [49:0] readslicef_51_50_1;
    input [50:0] vector;
    reg [50:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_51_50_1 = tmp[49:0];
  end
  endfunction
  function [0:0] readslicef_5_1_4;
    input [4:0] vector;
    reg [4:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_5_1_4 = tmp[0:0];
  end
  endfunction
  function [0:0] readslicef_6_1_5;
    input [5:0] vector;
    reg [5:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_6_1_5 = tmp[0:0];
  end
  endfunction
  function [0:0] readslicef_7_1_6;
    input [6:0] vector;
    reg [6:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_7_1_6 = tmp[0:0];
  end
  endfunction
  function [5:0] readslicef_7_6_1;
    input [6:0] vector;
    reg [6:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_7_6_1 = tmp[5:0];
  end
  endfunction
  function [0:0] readslicef_8_1_7;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_8_1_7 = tmp[0:0];
  end
  endfunction
  function [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction
  function [7:0] readslicef_9_8_1;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_9_8_1 = tmp[7:0];
  end
  endfunction
  function [9:0] signext_10_1;
    input [0:0] vector;
  begin
    signext_10_1= {{9{vector[0]}}, vector};
  end
  endfunction
  function [9:0] signext_10_5;
    input [4:0] vector;
  begin
    signext_10_5= {{5{vector[4]}}, vector};
  end
  endfunction
  function [2:0] signext_3_1;
    input [0:0] vector;
  begin
    signext_3_1= {{2{vector[0]}}, vector};
  end
  endfunction
  function [3:0] signext_4_1;
    input [0:0] vector;
  begin
    signext_4_1= {{3{vector[0]}}, vector};
  end
  endfunction
  function [7:0] conv_s2s_7_8 ;
    input [6:0] vector ;
  begin
    conv_s2s_7_8 = {vector[6], vector};
  end
  endfunction
  function [32:0] conv_s2s_16_33 ;
    input [15:0] vector ;
  begin
    conv_s2s_16_33 = {{17{vector[15]}}, vector};
  end
  endfunction
  function [32:0] conv_s2s_32_33 ;
    input [31:0] vector ;
  begin
    conv_s2s_32_33 = {vector[31], vector};
  end
  endfunction
  function [52:0] conv_s2s_51_53 ;
    input [50:0] vector ;
  begin
    conv_s2s_51_53 = {{2{vector[50]}}, vector};
  end
  endfunction
  function [52:0] conv_s2s_52_53 ;
    input [51:0] vector ;
  begin
    conv_s2s_52_53 = {vector[51], vector};
  end
  endfunction
  function [66:0] conv_s2s_66_67 ;
    input [65:0] vector ;
  begin
    conv_s2s_66_67 = {vector[65], vector};
  end
  endfunction
  function [2:0] conv_s2u_2_3 ;
    input [1:0] vector ;
  begin
    conv_s2u_2_3 = {vector[1], vector};
  end
  endfunction
  function [6:0] conv_s2u_6_7 ;
    input [5:0] vector ;
  begin
    conv_s2u_6_7 = {vector[5], vector};
  end
  endfunction
  function [33:0] conv_s2u_33_34 ;
    input [32:0] vector ;
  begin
    conv_s2u_33_34 = {vector[32], vector};
  end
  endfunction
  function [49:0] conv_s2u_50_50 ;
    input [49:0] vector ;
  begin
    conv_s2u_50_50 = vector;
  end
  endfunction
  function [17:0] conv_u2s_1_18 ;
    input [0:0] vector ;
  begin
    conv_u2s_1_18 = {{17{1'b0}}, vector};
  end
  endfunction
  function [66:0] conv_u2s_1_67 ;
    input [0:0] vector ;
  begin
    conv_u2s_1_67 = {{66{1'b0}}, vector};
  end
  endfunction
  function [6:0] conv_u2s_5_7 ;
    input [4:0] vector ;
  begin
    conv_u2s_5_7 = {{2{1'b0}}, vector};
  end
  endfunction
  function [6:0] conv_u2s_6_7 ;
    input [5:0] vector ;
  begin
    conv_u2s_6_7 = {1'b0, vector};
  end
  endfunction
  function [7:0] conv_u2s_6_8 ;
    input [5:0] vector ;
  begin
    conv_u2s_6_8 = {{2{1'b0}}, vector};
  end
  endfunction
  function [8:0] conv_u2s_6_9 ;
    input [5:0] vector ;
  begin
    conv_u2s_6_9 = {{3{1'b0}}, vector};
  end
  endfunction
  function [8:0] conv_u2s_8_9 ;
    input [7:0] vector ;
  begin
    conv_u2s_8_9 = {1'b0, vector};
  end
  endfunction
  function [35:0] conv_u2s_35_36 ;
    input [34:0] vector ;
  begin
    conv_u2s_35_36 = {1'b0, vector};
  end
  endfunction
  function [36:0] conv_u2s_36_37 ;
    input [35:0] vector ;
  begin
    conv_u2s_36_37 = {1'b0, vector};
  end
  endfunction
  function [9:0] conv_u2u_1_10 ;
    input [0:0] vector ;
  begin
    conv_u2u_1_10 = {{9{1'b0}}, vector};
  end
  endfunction
  function [10:0] conv_u2u_1_11 ;
    input [0:0] vector ;
  begin
    conv_u2u_1_11 = {{10{1'b0}}, vector};
  end
  endfunction
  function [22:0] conv_u2u_1_23 ;
    input [0:0] vector ;
  begin
    conv_u2u_1_23 = {{22{1'b0}}, vector};
  end
  endfunction
  function [2:0] conv_u2u_2_3 ;
    input [1:0] vector ;
  begin
    conv_u2u_2_3 = {1'b0, vector};
  end
  endfunction
  function [4:0] conv_u2u_4_5 ;
    input [3:0] vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction
  function [5:0] conv_u2u_5_6 ;
    input [4:0] vector ;
  begin
    conv_u2u_5_6 = {1'b0, vector};
  end
  endfunction
  function [6:0] conv_u2u_6_7 ;
    input [5:0] vector ;
  begin
    conv_u2u_6_7 = {1'b0, vector};
  end
  endfunction
  function [7:0] conv_u2u_7_8 ;
    input [6:0] vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction
  function [8:0] conv_u2u_8_9 ;
    input [7:0] vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction
  function [10:0] conv_u2u_10_11 ;
    input [9:0] vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction
  function [21:0] conv_u2u_22_22 ;
    input [21:0] vector ;
  begin
    conv_u2u_22_22 = vector;
  end
  endfunction
  function [23:0] conv_u2u_23_24 ;
    input [22:0] vector ;
  begin
    conv_u2u_23_24 = {1'b0, vector};
  end
  endfunction
  function [49:0] conv_u2u_49_50 ;
    input [48:0] vector ;
  begin
    conv_u2u_49_50 = {1'b0, vector};
  end
  endfunction
  function [50:0] conv_u2u_50_51 ;
    input [49:0] vector ;
  begin
    conv_u2u_50_51 = {1'b0, vector};
  end
  endfunction
endmodule
// ------------------------------------------------------------------
// Design Unit: NV_NVDLA_SDP_CORE_Y_inp
// ------------------------------------------------------------------
module NV_NVDLA_SDP_CORE_Y_inp (
  nvdla_core_clk, nvdla_core_rstn, chn_inp_in_rsc_z, chn_inp_in_rsc_vz, chn_inp_in_rsc_lz,
      cfg_precision_rsc_z, chn_inp_out_rsc_z, chn_inp_out_rsc_vz, chn_inp_out_rsc_lz
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [739:0] chn_inp_in_rsc_z;
  input chn_inp_in_rsc_vz;
  output chn_inp_in_rsc_lz;
  input [1:0] cfg_precision_rsc_z;
  output [127:0] chn_inp_out_rsc_z;
  input chn_inp_out_rsc_vz;
  output chn_inp_out_rsc_lz;
// Interconnect Declarations
  wire chn_inp_in_rsci_oswt;
  wire chn_inp_in_rsci_oswt_unreg;
  wire chn_inp_out_rsci_oswt;
  wire chn_inp_out_rsci_oswt_unreg;
// Interconnect Declarations for Component Instantiations
  SDP_Y_INP_chn_inp_in_rsci_unreg chn_inp_in_rsci_unreg_inst (
      .in_0(chn_inp_in_rsci_oswt_unreg),
      .outsig(chn_inp_in_rsci_oswt)
    );
  SDP_Y_INP_chn_inp_out_rsci_unreg chn_inp_out_rsci_unreg_inst (
      .in_0(chn_inp_out_rsci_oswt_unreg),
      .outsig(chn_inp_out_rsci_oswt)
    );
  NV_NVDLA_SDP_CORE_Y_inp_core NV_NVDLA_SDP_CORE_Y_inp_core_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_inp_in_rsc_z(chn_inp_in_rsc_z),
      .chn_inp_in_rsc_vz(chn_inp_in_rsc_vz),
      .chn_inp_in_rsc_lz(chn_inp_in_rsc_lz),
      .cfg_precision_rsc_z(cfg_precision_rsc_z),
      .chn_inp_out_rsc_z(chn_inp_out_rsc_z),
      .chn_inp_out_rsc_vz(chn_inp_out_rsc_vz),
      .chn_inp_out_rsc_lz(chn_inp_out_rsc_lz),
      .chn_inp_in_rsci_oswt(chn_inp_in_rsci_oswt),
      .chn_inp_in_rsci_oswt_unreg(chn_inp_in_rsci_oswt_unreg),
      .chn_inp_out_rsci_oswt(chn_inp_out_rsci_oswt),
      .chn_inp_out_rsci_oswt_unreg(chn_inp_out_rsci_oswt_unreg)
    );
endmodule
