`timescale 10ps/1ps
module NV_NVDLA_PDP_CORE_med2d_lut(
    input  [7 : 0] encoding,
    input  [7 : 0] decoding,
    input  [7 : 0][3 : 0][3 : 0] msbs_i,
    input  [7 : 0][3 : 0][3 : 0] msbs_j,
    input  [7 : 0][3 : 0][3 : 0] msbs_k,
    input  [7 : 0][3 : 0][3 : 0] msbs_w,
    output [7 : 0][3 : 0][11 : 0] code_o,
    input  [7 : 0][3 : 0][11 : 0] to_decode,
    output  [7 : 0][3 : 0][3 : 0] decoded_msbs_i,
    output  [7 : 0][3 : 0][3 : 0] decoded_msbs_j,
    output  [7 : 0][3 : 0][3 : 0] decoded_msbs_k,
    output  [7 : 0][3 : 0][3 : 0] decoded_msbs_w
);

wire [3876 : 1][15 : 0] lut_table; 
reg  [7 : 0][3 : 0][11 : 0] code;
reg  [7 : 0][3 : 0][3 : 0] decoded_msbs_i_reg;
reg  [7 : 0][3 : 0][3 : 0] decoded_msbs_j_reg;
reg  [7 : 0][3 : 0][3 : 0] decoded_msbs_k_reg;
reg  [7 : 0][3 : 0][3 : 0] decoded_msbs_w_reg;


assign lut_table[1] = 16'b0000000000000000; 
assign lut_table[2] = 16'b0000000000000001; 
assign lut_table[3] = 16'b0000000000000010; 
assign lut_table[4] = 16'b0000000000000011; 
assign lut_table[5] = 16'b0000000000000100; 
assign lut_table[6] = 16'b0000000000000101; 
assign lut_table[7] = 16'b0000000000000110; 
assign lut_table[8] = 16'b0000000000000111; 
assign lut_table[9] = 16'b0000000000001000; 
assign lut_table[10] = 16'b0000000000001001; 
assign lut_table[11] = 16'b0000000000001010; 
assign lut_table[12] = 16'b0000000000001011; 
assign lut_table[13] = 16'b0000000000001100; 
assign lut_table[14] = 16'b0000000000001101; 
assign lut_table[15] = 16'b0000000000001110; 
assign lut_table[16] = 16'b0000000000001111; 
assign lut_table[17] = 16'b0000000000010001; 
assign lut_table[18] = 16'b0000000000010010; 
assign lut_table[19] = 16'b0000000000010011; 
assign lut_table[20] = 16'b0000000000010100; 
assign lut_table[21] = 16'b0000000000010101; 
assign lut_table[22] = 16'b0000000000010110; 
assign lut_table[23] = 16'b0000000000010111; 
assign lut_table[24] = 16'b0000000000011000; 
assign lut_table[25] = 16'b0000000000011001; 
assign lut_table[26] = 16'b0000000000011010; 
assign lut_table[27] = 16'b0000000000011011; 
assign lut_table[28] = 16'b0000000000011100; 
assign lut_table[29] = 16'b0000000000011101; 
assign lut_table[30] = 16'b0000000000011110; 
assign lut_table[31] = 16'b0000000000011111; 
assign lut_table[32] = 16'b0000000000100010; 
assign lut_table[33] = 16'b0000000000100011; 
assign lut_table[34] = 16'b0000000000100100; 
assign lut_table[35] = 16'b0000000000100101; 
assign lut_table[36] = 16'b0000000000100110; 
assign lut_table[37] = 16'b0000000000100111; 
assign lut_table[38] = 16'b0000000000101000; 
assign lut_table[39] = 16'b0000000000101001; 
assign lut_table[40] = 16'b0000000000101010; 
assign lut_table[41] = 16'b0000000000101011; 
assign lut_table[42] = 16'b0000000000101100; 
assign lut_table[43] = 16'b0000000000101101; 
assign lut_table[44] = 16'b0000000000101110; 
assign lut_table[45] = 16'b0000000000101111; 
assign lut_table[46] = 16'b0000000000110011; 
assign lut_table[47] = 16'b0000000000110100; 
assign lut_table[48] = 16'b0000000000110101; 
assign lut_table[49] = 16'b0000000000110110; 
assign lut_table[50] = 16'b0000000000110111; 
assign lut_table[51] = 16'b0000000000111000; 
assign lut_table[52] = 16'b0000000000111001; 
assign lut_table[53] = 16'b0000000000111010; 
assign lut_table[54] = 16'b0000000000111011; 
assign lut_table[55] = 16'b0000000000111100; 
assign lut_table[56] = 16'b0000000000111101; 
assign lut_table[57] = 16'b0000000000111110; 
assign lut_table[58] = 16'b0000000000111111; 
assign lut_table[59] = 16'b0000000001000100; 
assign lut_table[60] = 16'b0000000001000101; 
assign lut_table[61] = 16'b0000000001000110; 
assign lut_table[62] = 16'b0000000001000111; 
assign lut_table[63] = 16'b0000000001001000; 
assign lut_table[64] = 16'b0000000001001001; 
assign lut_table[65] = 16'b0000000001001010; 
assign lut_table[66] = 16'b0000000001001011; 
assign lut_table[67] = 16'b0000000001001100; 
assign lut_table[68] = 16'b0000000001001101; 
assign lut_table[69] = 16'b0000000001001110; 
assign lut_table[70] = 16'b0000000001001111; 
assign lut_table[71] = 16'b0000000001010101; 
assign lut_table[72] = 16'b0000000001010110; 
assign lut_table[73] = 16'b0000000001010111; 
assign lut_table[74] = 16'b0000000001011000; 
assign lut_table[75] = 16'b0000000001011001; 
assign lut_table[76] = 16'b0000000001011010; 
assign lut_table[77] = 16'b0000000001011011; 
assign lut_table[78] = 16'b0000000001011100; 
assign lut_table[79] = 16'b0000000001011101; 
assign lut_table[80] = 16'b0000000001011110; 
assign lut_table[81] = 16'b0000000001011111; 
assign lut_table[82] = 16'b0000000001100110; 
assign lut_table[83] = 16'b0000000001100111; 
assign lut_table[84] = 16'b0000000001101000; 
assign lut_table[85] = 16'b0000000001101001; 
assign lut_table[86] = 16'b0000000001101010; 
assign lut_table[87] = 16'b0000000001101011; 
assign lut_table[88] = 16'b0000000001101100; 
assign lut_table[89] = 16'b0000000001101101; 
assign lut_table[90] = 16'b0000000001101110; 
assign lut_table[91] = 16'b0000000001101111; 
assign lut_table[92] = 16'b0000000001110111; 
assign lut_table[93] = 16'b0000000001111000; 
assign lut_table[94] = 16'b0000000001111001; 
assign lut_table[95] = 16'b0000000001111010; 
assign lut_table[96] = 16'b0000000001111011; 
assign lut_table[97] = 16'b0000000001111100; 
assign lut_table[98] = 16'b0000000001111101; 
assign lut_table[99] = 16'b0000000001111110; 
assign lut_table[100] = 16'b0000000001111111; 
assign lut_table[101] = 16'b0000000010001000; 
assign lut_table[102] = 16'b0000000010001001; 
assign lut_table[103] = 16'b0000000010001010; 
assign lut_table[104] = 16'b0000000010001011; 
assign lut_table[105] = 16'b0000000010001100; 
assign lut_table[106] = 16'b0000000010001101; 
assign lut_table[107] = 16'b0000000010001110; 
assign lut_table[108] = 16'b0000000010001111; 
assign lut_table[109] = 16'b0000000010011001; 
assign lut_table[110] = 16'b0000000010011010; 
assign lut_table[111] = 16'b0000000010011011; 
assign lut_table[112] = 16'b0000000010011100; 
assign lut_table[113] = 16'b0000000010011101; 
assign lut_table[114] = 16'b0000000010011110; 
assign lut_table[115] = 16'b0000000010011111; 
assign lut_table[116] = 16'b0000000010101010; 
assign lut_table[117] = 16'b0000000010101011; 
assign lut_table[118] = 16'b0000000010101100; 
assign lut_table[119] = 16'b0000000010101101; 
assign lut_table[120] = 16'b0000000010101110; 
assign lut_table[121] = 16'b0000000010101111; 
assign lut_table[122] = 16'b0000000010111011; 
assign lut_table[123] = 16'b0000000010111100; 
assign lut_table[124] = 16'b0000000010111101; 
assign lut_table[125] = 16'b0000000010111110; 
assign lut_table[126] = 16'b0000000010111111; 
assign lut_table[127] = 16'b0000000011001100; 
assign lut_table[128] = 16'b0000000011001101; 
assign lut_table[129] = 16'b0000000011001110; 
assign lut_table[130] = 16'b0000000011001111; 
assign lut_table[131] = 16'b0000000011011101; 
assign lut_table[132] = 16'b0000000011011110; 
assign lut_table[133] = 16'b0000000011011111; 
assign lut_table[134] = 16'b0000000011101110; 
assign lut_table[135] = 16'b0000000011101111; 
assign lut_table[136] = 16'b0000000011111111; 
assign lut_table[137] = 16'b0000000100010001; 
assign lut_table[138] = 16'b0000000100010010; 
assign lut_table[139] = 16'b0000000100010011; 
assign lut_table[140] = 16'b0000000100010100; 
assign lut_table[141] = 16'b0000000100010101; 
assign lut_table[142] = 16'b0000000100010110; 
assign lut_table[143] = 16'b0000000100010111; 
assign lut_table[144] = 16'b0000000100011000; 
assign lut_table[145] = 16'b0000000100011001; 
assign lut_table[146] = 16'b0000000100011010; 
assign lut_table[147] = 16'b0000000100011011; 
assign lut_table[148] = 16'b0000000100011100; 
assign lut_table[149] = 16'b0000000100011101; 
assign lut_table[150] = 16'b0000000100011110; 
assign lut_table[151] = 16'b0000000100011111; 
assign lut_table[152] = 16'b0000000100100010; 
assign lut_table[153] = 16'b0000000100100011; 
assign lut_table[154] = 16'b0000000100100100; 
assign lut_table[155] = 16'b0000000100100101; 
assign lut_table[156] = 16'b0000000100100110; 
assign lut_table[157] = 16'b0000000100100111; 
assign lut_table[158] = 16'b0000000100101000; 
assign lut_table[159] = 16'b0000000100101001; 
assign lut_table[160] = 16'b0000000100101010; 
assign lut_table[161] = 16'b0000000100101011; 
assign lut_table[162] = 16'b0000000100101100; 
assign lut_table[163] = 16'b0000000100101101; 
assign lut_table[164] = 16'b0000000100101110; 
assign lut_table[165] = 16'b0000000100101111; 
assign lut_table[166] = 16'b0000000100110011; 
assign lut_table[167] = 16'b0000000100110100; 
assign lut_table[168] = 16'b0000000100110101; 
assign lut_table[169] = 16'b0000000100110110; 
assign lut_table[170] = 16'b0000000100110111; 
assign lut_table[171] = 16'b0000000100111000; 
assign lut_table[172] = 16'b0000000100111001; 
assign lut_table[173] = 16'b0000000100111010; 
assign lut_table[174] = 16'b0000000100111011; 
assign lut_table[175] = 16'b0000000100111100; 
assign lut_table[176] = 16'b0000000100111101; 
assign lut_table[177] = 16'b0000000100111110; 
assign lut_table[178] = 16'b0000000100111111; 
assign lut_table[179] = 16'b0000000101000100; 
assign lut_table[180] = 16'b0000000101000101; 
assign lut_table[181] = 16'b0000000101000110; 
assign lut_table[182] = 16'b0000000101000111; 
assign lut_table[183] = 16'b0000000101001000; 
assign lut_table[184] = 16'b0000000101001001; 
assign lut_table[185] = 16'b0000000101001010; 
assign lut_table[186] = 16'b0000000101001011; 
assign lut_table[187] = 16'b0000000101001100; 
assign lut_table[188] = 16'b0000000101001101; 
assign lut_table[189] = 16'b0000000101001110; 
assign lut_table[190] = 16'b0000000101001111; 
assign lut_table[191] = 16'b0000000101010101; 
assign lut_table[192] = 16'b0000000101010110; 
assign lut_table[193] = 16'b0000000101010111; 
assign lut_table[194] = 16'b0000000101011000; 
assign lut_table[195] = 16'b0000000101011001; 
assign lut_table[196] = 16'b0000000101011010; 
assign lut_table[197] = 16'b0000000101011011; 
assign lut_table[198] = 16'b0000000101011100; 
assign lut_table[199] = 16'b0000000101011101; 
assign lut_table[200] = 16'b0000000101011110; 
assign lut_table[201] = 16'b0000000101011111; 
assign lut_table[202] = 16'b0000000101100110; 
assign lut_table[203] = 16'b0000000101100111; 
assign lut_table[204] = 16'b0000000101101000; 
assign lut_table[205] = 16'b0000000101101001; 
assign lut_table[206] = 16'b0000000101101010; 
assign lut_table[207] = 16'b0000000101101011; 
assign lut_table[208] = 16'b0000000101101100; 
assign lut_table[209] = 16'b0000000101101101; 
assign lut_table[210] = 16'b0000000101101110; 
assign lut_table[211] = 16'b0000000101101111; 
assign lut_table[212] = 16'b0000000101110111; 
assign lut_table[213] = 16'b0000000101111000; 
assign lut_table[214] = 16'b0000000101111001; 
assign lut_table[215] = 16'b0000000101111010; 
assign lut_table[216] = 16'b0000000101111011; 
assign lut_table[217] = 16'b0000000101111100; 
assign lut_table[218] = 16'b0000000101111101; 
assign lut_table[219] = 16'b0000000101111110; 
assign lut_table[220] = 16'b0000000101111111; 
assign lut_table[221] = 16'b0000000110001000; 
assign lut_table[222] = 16'b0000000110001001; 
assign lut_table[223] = 16'b0000000110001010; 
assign lut_table[224] = 16'b0000000110001011; 
assign lut_table[225] = 16'b0000000110001100; 
assign lut_table[226] = 16'b0000000110001101; 
assign lut_table[227] = 16'b0000000110001110; 
assign lut_table[228] = 16'b0000000110001111; 
assign lut_table[229] = 16'b0000000110011001; 
assign lut_table[230] = 16'b0000000110011010; 
assign lut_table[231] = 16'b0000000110011011; 
assign lut_table[232] = 16'b0000000110011100; 
assign lut_table[233] = 16'b0000000110011101; 
assign lut_table[234] = 16'b0000000110011110; 
assign lut_table[235] = 16'b0000000110011111; 
assign lut_table[236] = 16'b0000000110101010; 
assign lut_table[237] = 16'b0000000110101011; 
assign lut_table[238] = 16'b0000000110101100; 
assign lut_table[239] = 16'b0000000110101101; 
assign lut_table[240] = 16'b0000000110101110; 
assign lut_table[241] = 16'b0000000110101111; 
assign lut_table[242] = 16'b0000000110111011; 
assign lut_table[243] = 16'b0000000110111100; 
assign lut_table[244] = 16'b0000000110111101; 
assign lut_table[245] = 16'b0000000110111110; 
assign lut_table[246] = 16'b0000000110111111; 
assign lut_table[247] = 16'b0000000111001100; 
assign lut_table[248] = 16'b0000000111001101; 
assign lut_table[249] = 16'b0000000111001110; 
assign lut_table[250] = 16'b0000000111001111; 
assign lut_table[251] = 16'b0000000111011101; 
assign lut_table[252] = 16'b0000000111011110; 
assign lut_table[253] = 16'b0000000111011111; 
assign lut_table[254] = 16'b0000000111101110; 
assign lut_table[255] = 16'b0000000111101111; 
assign lut_table[256] = 16'b0000000111111111; 
assign lut_table[257] = 16'b0000001000100010; 
assign lut_table[258] = 16'b0000001000100011; 
assign lut_table[259] = 16'b0000001000100100; 
assign lut_table[260] = 16'b0000001000100101; 
assign lut_table[261] = 16'b0000001000100110; 
assign lut_table[262] = 16'b0000001000100111; 
assign lut_table[263] = 16'b0000001000101000; 
assign lut_table[264] = 16'b0000001000101001; 
assign lut_table[265] = 16'b0000001000101010; 
assign lut_table[266] = 16'b0000001000101011; 
assign lut_table[267] = 16'b0000001000101100; 
assign lut_table[268] = 16'b0000001000101101; 
assign lut_table[269] = 16'b0000001000101110; 
assign lut_table[270] = 16'b0000001000101111; 
assign lut_table[271] = 16'b0000001000110011; 
assign lut_table[272] = 16'b0000001000110100; 
assign lut_table[273] = 16'b0000001000110101; 
assign lut_table[274] = 16'b0000001000110110; 
assign lut_table[275] = 16'b0000001000110111; 
assign lut_table[276] = 16'b0000001000111000; 
assign lut_table[277] = 16'b0000001000111001; 
assign lut_table[278] = 16'b0000001000111010; 
assign lut_table[279] = 16'b0000001000111011; 
assign lut_table[280] = 16'b0000001000111100; 
assign lut_table[281] = 16'b0000001000111101; 
assign lut_table[282] = 16'b0000001000111110; 
assign lut_table[283] = 16'b0000001000111111; 
assign lut_table[284] = 16'b0000001001000100; 
assign lut_table[285] = 16'b0000001001000101; 
assign lut_table[286] = 16'b0000001001000110; 
assign lut_table[287] = 16'b0000001001000111; 
assign lut_table[288] = 16'b0000001001001000; 
assign lut_table[289] = 16'b0000001001001001; 
assign lut_table[290] = 16'b0000001001001010; 
assign lut_table[291] = 16'b0000001001001011; 
assign lut_table[292] = 16'b0000001001001100; 
assign lut_table[293] = 16'b0000001001001101; 
assign lut_table[294] = 16'b0000001001001110; 
assign lut_table[295] = 16'b0000001001001111; 
assign lut_table[296] = 16'b0000001001010101; 
assign lut_table[297] = 16'b0000001001010110; 
assign lut_table[298] = 16'b0000001001010111; 
assign lut_table[299] = 16'b0000001001011000; 
assign lut_table[300] = 16'b0000001001011001; 
assign lut_table[301] = 16'b0000001001011010; 
assign lut_table[302] = 16'b0000001001011011; 
assign lut_table[303] = 16'b0000001001011100; 
assign lut_table[304] = 16'b0000001001011101; 
assign lut_table[305] = 16'b0000001001011110; 
assign lut_table[306] = 16'b0000001001011111; 
assign lut_table[307] = 16'b0000001001100110; 
assign lut_table[308] = 16'b0000001001100111; 
assign lut_table[309] = 16'b0000001001101000; 
assign lut_table[310] = 16'b0000001001101001; 
assign lut_table[311] = 16'b0000001001101010; 
assign lut_table[312] = 16'b0000001001101011; 
assign lut_table[313] = 16'b0000001001101100; 
assign lut_table[314] = 16'b0000001001101101; 
assign lut_table[315] = 16'b0000001001101110; 
assign lut_table[316] = 16'b0000001001101111; 
assign lut_table[317] = 16'b0000001001110111; 
assign lut_table[318] = 16'b0000001001111000; 
assign lut_table[319] = 16'b0000001001111001; 
assign lut_table[320] = 16'b0000001001111010; 
assign lut_table[321] = 16'b0000001001111011; 
assign lut_table[322] = 16'b0000001001111100; 
assign lut_table[323] = 16'b0000001001111101; 
assign lut_table[324] = 16'b0000001001111110; 
assign lut_table[325] = 16'b0000001001111111; 
assign lut_table[326] = 16'b0000001010001000; 
assign lut_table[327] = 16'b0000001010001001; 
assign lut_table[328] = 16'b0000001010001010; 
assign lut_table[329] = 16'b0000001010001011; 
assign lut_table[330] = 16'b0000001010001100; 
assign lut_table[331] = 16'b0000001010001101; 
assign lut_table[332] = 16'b0000001010001110; 
assign lut_table[333] = 16'b0000001010001111; 
assign lut_table[334] = 16'b0000001010011001; 
assign lut_table[335] = 16'b0000001010011010; 
assign lut_table[336] = 16'b0000001010011011; 
assign lut_table[337] = 16'b0000001010011100; 
assign lut_table[338] = 16'b0000001010011101; 
assign lut_table[339] = 16'b0000001010011110; 
assign lut_table[340] = 16'b0000001010011111; 
assign lut_table[341] = 16'b0000001010101010; 
assign lut_table[342] = 16'b0000001010101011; 
assign lut_table[343] = 16'b0000001010101100; 
assign lut_table[344] = 16'b0000001010101101; 
assign lut_table[345] = 16'b0000001010101110; 
assign lut_table[346] = 16'b0000001010101111; 
assign lut_table[347] = 16'b0000001010111011; 
assign lut_table[348] = 16'b0000001010111100; 
assign lut_table[349] = 16'b0000001010111101; 
assign lut_table[350] = 16'b0000001010111110; 
assign lut_table[351] = 16'b0000001010111111; 
assign lut_table[352] = 16'b0000001011001100; 
assign lut_table[353] = 16'b0000001011001101; 
assign lut_table[354] = 16'b0000001011001110; 
assign lut_table[355] = 16'b0000001011001111; 
assign lut_table[356] = 16'b0000001011011101; 
assign lut_table[357] = 16'b0000001011011110; 
assign lut_table[358] = 16'b0000001011011111; 
assign lut_table[359] = 16'b0000001011101110; 
assign lut_table[360] = 16'b0000001011101111; 
assign lut_table[361] = 16'b0000001011111111; 
assign lut_table[362] = 16'b0000001100110011; 
assign lut_table[363] = 16'b0000001100110100; 
assign lut_table[364] = 16'b0000001100110101; 
assign lut_table[365] = 16'b0000001100110110; 
assign lut_table[366] = 16'b0000001100110111; 
assign lut_table[367] = 16'b0000001100111000; 
assign lut_table[368] = 16'b0000001100111001; 
assign lut_table[369] = 16'b0000001100111010; 
assign lut_table[370] = 16'b0000001100111011; 
assign lut_table[371] = 16'b0000001100111100; 
assign lut_table[372] = 16'b0000001100111101; 
assign lut_table[373] = 16'b0000001100111110; 
assign lut_table[374] = 16'b0000001100111111; 
assign lut_table[375] = 16'b0000001101000100; 
assign lut_table[376] = 16'b0000001101000101; 
assign lut_table[377] = 16'b0000001101000110; 
assign lut_table[378] = 16'b0000001101000111; 
assign lut_table[379] = 16'b0000001101001000; 
assign lut_table[380] = 16'b0000001101001001; 
assign lut_table[381] = 16'b0000001101001010; 
assign lut_table[382] = 16'b0000001101001011; 
assign lut_table[383] = 16'b0000001101001100; 
assign lut_table[384] = 16'b0000001101001101; 
assign lut_table[385] = 16'b0000001101001110; 
assign lut_table[386] = 16'b0000001101001111; 
assign lut_table[387] = 16'b0000001101010101; 
assign lut_table[388] = 16'b0000001101010110; 
assign lut_table[389] = 16'b0000001101010111; 
assign lut_table[390] = 16'b0000001101011000; 
assign lut_table[391] = 16'b0000001101011001; 
assign lut_table[392] = 16'b0000001101011010; 
assign lut_table[393] = 16'b0000001101011011; 
assign lut_table[394] = 16'b0000001101011100; 
assign lut_table[395] = 16'b0000001101011101; 
assign lut_table[396] = 16'b0000001101011110; 
assign lut_table[397] = 16'b0000001101011111; 
assign lut_table[398] = 16'b0000001101100110; 
assign lut_table[399] = 16'b0000001101100111; 
assign lut_table[400] = 16'b0000001101101000; 
assign lut_table[401] = 16'b0000001101101001; 
assign lut_table[402] = 16'b0000001101101010; 
assign lut_table[403] = 16'b0000001101101011; 
assign lut_table[404] = 16'b0000001101101100; 
assign lut_table[405] = 16'b0000001101101101; 
assign lut_table[406] = 16'b0000001101101110; 
assign lut_table[407] = 16'b0000001101101111; 
assign lut_table[408] = 16'b0000001101110111; 
assign lut_table[409] = 16'b0000001101111000; 
assign lut_table[410] = 16'b0000001101111001; 
assign lut_table[411] = 16'b0000001101111010; 
assign lut_table[412] = 16'b0000001101111011; 
assign lut_table[413] = 16'b0000001101111100; 
assign lut_table[414] = 16'b0000001101111101; 
assign lut_table[415] = 16'b0000001101111110; 
assign lut_table[416] = 16'b0000001101111111; 
assign lut_table[417] = 16'b0000001110001000; 
assign lut_table[418] = 16'b0000001110001001; 
assign lut_table[419] = 16'b0000001110001010; 
assign lut_table[420] = 16'b0000001110001011; 
assign lut_table[421] = 16'b0000001110001100; 
assign lut_table[422] = 16'b0000001110001101; 
assign lut_table[423] = 16'b0000001110001110; 
assign lut_table[424] = 16'b0000001110001111; 
assign lut_table[425] = 16'b0000001110011001; 
assign lut_table[426] = 16'b0000001110011010; 
assign lut_table[427] = 16'b0000001110011011; 
assign lut_table[428] = 16'b0000001110011100; 
assign lut_table[429] = 16'b0000001110011101; 
assign lut_table[430] = 16'b0000001110011110; 
assign lut_table[431] = 16'b0000001110011111; 
assign lut_table[432] = 16'b0000001110101010; 
assign lut_table[433] = 16'b0000001110101011; 
assign lut_table[434] = 16'b0000001110101100; 
assign lut_table[435] = 16'b0000001110101101; 
assign lut_table[436] = 16'b0000001110101110; 
assign lut_table[437] = 16'b0000001110101111; 
assign lut_table[438] = 16'b0000001110111011; 
assign lut_table[439] = 16'b0000001110111100; 
assign lut_table[440] = 16'b0000001110111101; 
assign lut_table[441] = 16'b0000001110111110; 
assign lut_table[442] = 16'b0000001110111111; 
assign lut_table[443] = 16'b0000001111001100; 
assign lut_table[444] = 16'b0000001111001101; 
assign lut_table[445] = 16'b0000001111001110; 
assign lut_table[446] = 16'b0000001111001111; 
assign lut_table[447] = 16'b0000001111011101; 
assign lut_table[448] = 16'b0000001111011110; 
assign lut_table[449] = 16'b0000001111011111; 
assign lut_table[450] = 16'b0000001111101110; 
assign lut_table[451] = 16'b0000001111101111; 
assign lut_table[452] = 16'b0000001111111111; 
assign lut_table[453] = 16'b0000010001000100; 
assign lut_table[454] = 16'b0000010001000101; 
assign lut_table[455] = 16'b0000010001000110; 
assign lut_table[456] = 16'b0000010001000111; 
assign lut_table[457] = 16'b0000010001001000; 
assign lut_table[458] = 16'b0000010001001001; 
assign lut_table[459] = 16'b0000010001001010; 
assign lut_table[460] = 16'b0000010001001011; 
assign lut_table[461] = 16'b0000010001001100; 
assign lut_table[462] = 16'b0000010001001101; 
assign lut_table[463] = 16'b0000010001001110; 
assign lut_table[464] = 16'b0000010001001111; 
assign lut_table[465] = 16'b0000010001010101; 
assign lut_table[466] = 16'b0000010001010110; 
assign lut_table[467] = 16'b0000010001010111; 
assign lut_table[468] = 16'b0000010001011000; 
assign lut_table[469] = 16'b0000010001011001; 
assign lut_table[470] = 16'b0000010001011010; 
assign lut_table[471] = 16'b0000010001011011; 
assign lut_table[472] = 16'b0000010001011100; 
assign lut_table[473] = 16'b0000010001011101; 
assign lut_table[474] = 16'b0000010001011110; 
assign lut_table[475] = 16'b0000010001011111; 
assign lut_table[476] = 16'b0000010001100110; 
assign lut_table[477] = 16'b0000010001100111; 
assign lut_table[478] = 16'b0000010001101000; 
assign lut_table[479] = 16'b0000010001101001; 
assign lut_table[480] = 16'b0000010001101010; 
assign lut_table[481] = 16'b0000010001101011; 
assign lut_table[482] = 16'b0000010001101100; 
assign lut_table[483] = 16'b0000010001101101; 
assign lut_table[484] = 16'b0000010001101110; 
assign lut_table[485] = 16'b0000010001101111; 
assign lut_table[486] = 16'b0000010001110111; 
assign lut_table[487] = 16'b0000010001111000; 
assign lut_table[488] = 16'b0000010001111001; 
assign lut_table[489] = 16'b0000010001111010; 
assign lut_table[490] = 16'b0000010001111011; 
assign lut_table[491] = 16'b0000010001111100; 
assign lut_table[492] = 16'b0000010001111101; 
assign lut_table[493] = 16'b0000010001111110; 
assign lut_table[494] = 16'b0000010001111111; 
assign lut_table[495] = 16'b0000010010001000; 
assign lut_table[496] = 16'b0000010010001001; 
assign lut_table[497] = 16'b0000010010001010; 
assign lut_table[498] = 16'b0000010010001011; 
assign lut_table[499] = 16'b0000010010001100; 
assign lut_table[500] = 16'b0000010010001101; 
assign lut_table[501] = 16'b0000010010001110; 
assign lut_table[502] = 16'b0000010010001111; 
assign lut_table[503] = 16'b0000010010011001; 
assign lut_table[504] = 16'b0000010010011010; 
assign lut_table[505] = 16'b0000010010011011; 
assign lut_table[506] = 16'b0000010010011100; 
assign lut_table[507] = 16'b0000010010011101; 
assign lut_table[508] = 16'b0000010010011110; 
assign lut_table[509] = 16'b0000010010011111; 
assign lut_table[510] = 16'b0000010010101010; 
assign lut_table[511] = 16'b0000010010101011; 
assign lut_table[512] = 16'b0000010010101100; 
assign lut_table[513] = 16'b0000010010101101; 
assign lut_table[514] = 16'b0000010010101110; 
assign lut_table[515] = 16'b0000010010101111; 
assign lut_table[516] = 16'b0000010010111011; 
assign lut_table[517] = 16'b0000010010111100; 
assign lut_table[518] = 16'b0000010010111101; 
assign lut_table[519] = 16'b0000010010111110; 
assign lut_table[520] = 16'b0000010010111111; 
assign lut_table[521] = 16'b0000010011001100; 
assign lut_table[522] = 16'b0000010011001101; 
assign lut_table[523] = 16'b0000010011001110; 
assign lut_table[524] = 16'b0000010011001111; 
assign lut_table[525] = 16'b0000010011011101; 
assign lut_table[526] = 16'b0000010011011110; 
assign lut_table[527] = 16'b0000010011011111; 
assign lut_table[528] = 16'b0000010011101110; 
assign lut_table[529] = 16'b0000010011101111; 
assign lut_table[530] = 16'b0000010011111111; 
assign lut_table[531] = 16'b0000010101010101; 
assign lut_table[532] = 16'b0000010101010110; 
assign lut_table[533] = 16'b0000010101010111; 
assign lut_table[534] = 16'b0000010101011000; 
assign lut_table[535] = 16'b0000010101011001; 
assign lut_table[536] = 16'b0000010101011010; 
assign lut_table[537] = 16'b0000010101011011; 
assign lut_table[538] = 16'b0000010101011100; 
assign lut_table[539] = 16'b0000010101011101; 
assign lut_table[540] = 16'b0000010101011110; 
assign lut_table[541] = 16'b0000010101011111; 
assign lut_table[542] = 16'b0000010101100110; 
assign lut_table[543] = 16'b0000010101100111; 
assign lut_table[544] = 16'b0000010101101000; 
assign lut_table[545] = 16'b0000010101101001; 
assign lut_table[546] = 16'b0000010101101010; 
assign lut_table[547] = 16'b0000010101101011; 
assign lut_table[548] = 16'b0000010101101100; 
assign lut_table[549] = 16'b0000010101101101; 
assign lut_table[550] = 16'b0000010101101110; 
assign lut_table[551] = 16'b0000010101101111; 
assign lut_table[552] = 16'b0000010101110111; 
assign lut_table[553] = 16'b0000010101111000; 
assign lut_table[554] = 16'b0000010101111001; 
assign lut_table[555] = 16'b0000010101111010; 
assign lut_table[556] = 16'b0000010101111011; 
assign lut_table[557] = 16'b0000010101111100; 
assign lut_table[558] = 16'b0000010101111101; 
assign lut_table[559] = 16'b0000010101111110; 
assign lut_table[560] = 16'b0000010101111111; 
assign lut_table[561] = 16'b0000010110001000; 
assign lut_table[562] = 16'b0000010110001001; 
assign lut_table[563] = 16'b0000010110001010; 
assign lut_table[564] = 16'b0000010110001011; 
assign lut_table[565] = 16'b0000010110001100; 
assign lut_table[566] = 16'b0000010110001101; 
assign lut_table[567] = 16'b0000010110001110; 
assign lut_table[568] = 16'b0000010110001111; 
assign lut_table[569] = 16'b0000010110011001; 
assign lut_table[570] = 16'b0000010110011010; 
assign lut_table[571] = 16'b0000010110011011; 
assign lut_table[572] = 16'b0000010110011100; 
assign lut_table[573] = 16'b0000010110011101; 
assign lut_table[574] = 16'b0000010110011110; 
assign lut_table[575] = 16'b0000010110011111; 
assign lut_table[576] = 16'b0000010110101010; 
assign lut_table[577] = 16'b0000010110101011; 
assign lut_table[578] = 16'b0000010110101100; 
assign lut_table[579] = 16'b0000010110101101; 
assign lut_table[580] = 16'b0000010110101110; 
assign lut_table[581] = 16'b0000010110101111; 
assign lut_table[582] = 16'b0000010110111011; 
assign lut_table[583] = 16'b0000010110111100; 
assign lut_table[584] = 16'b0000010110111101; 
assign lut_table[585] = 16'b0000010110111110; 
assign lut_table[586] = 16'b0000010110111111; 
assign lut_table[587] = 16'b0000010111001100; 
assign lut_table[588] = 16'b0000010111001101; 
assign lut_table[589] = 16'b0000010111001110; 
assign lut_table[590] = 16'b0000010111001111; 
assign lut_table[591] = 16'b0000010111011101; 
assign lut_table[592] = 16'b0000010111011110; 
assign lut_table[593] = 16'b0000010111011111; 
assign lut_table[594] = 16'b0000010111101110; 
assign lut_table[595] = 16'b0000010111101111; 
assign lut_table[596] = 16'b0000010111111111; 
assign lut_table[597] = 16'b0000011001100110; 
assign lut_table[598] = 16'b0000011001100111; 
assign lut_table[599] = 16'b0000011001101000; 
assign lut_table[600] = 16'b0000011001101001; 
assign lut_table[601] = 16'b0000011001101010; 
assign lut_table[602] = 16'b0000011001101011; 
assign lut_table[603] = 16'b0000011001101100; 
assign lut_table[604] = 16'b0000011001101101; 
assign lut_table[605] = 16'b0000011001101110; 
assign lut_table[606] = 16'b0000011001101111; 
assign lut_table[607] = 16'b0000011001110111; 
assign lut_table[608] = 16'b0000011001111000; 
assign lut_table[609] = 16'b0000011001111001; 
assign lut_table[610] = 16'b0000011001111010; 
assign lut_table[611] = 16'b0000011001111011; 
assign lut_table[612] = 16'b0000011001111100; 
assign lut_table[613] = 16'b0000011001111101; 
assign lut_table[614] = 16'b0000011001111110; 
assign lut_table[615] = 16'b0000011001111111; 
assign lut_table[616] = 16'b0000011010001000; 
assign lut_table[617] = 16'b0000011010001001; 
assign lut_table[618] = 16'b0000011010001010; 
assign lut_table[619] = 16'b0000011010001011; 
assign lut_table[620] = 16'b0000011010001100; 
assign lut_table[621] = 16'b0000011010001101; 
assign lut_table[622] = 16'b0000011010001110; 
assign lut_table[623] = 16'b0000011010001111; 
assign lut_table[624] = 16'b0000011010011001; 
assign lut_table[625] = 16'b0000011010011010; 
assign lut_table[626] = 16'b0000011010011011; 
assign lut_table[627] = 16'b0000011010011100; 
assign lut_table[628] = 16'b0000011010011101; 
assign lut_table[629] = 16'b0000011010011110; 
assign lut_table[630] = 16'b0000011010011111; 
assign lut_table[631] = 16'b0000011010101010; 
assign lut_table[632] = 16'b0000011010101011; 
assign lut_table[633] = 16'b0000011010101100; 
assign lut_table[634] = 16'b0000011010101101; 
assign lut_table[635] = 16'b0000011010101110; 
assign lut_table[636] = 16'b0000011010101111; 
assign lut_table[637] = 16'b0000011010111011; 
assign lut_table[638] = 16'b0000011010111100; 
assign lut_table[639] = 16'b0000011010111101; 
assign lut_table[640] = 16'b0000011010111110; 
assign lut_table[641] = 16'b0000011010111111; 
assign lut_table[642] = 16'b0000011011001100; 
assign lut_table[643] = 16'b0000011011001101; 
assign lut_table[644] = 16'b0000011011001110; 
assign lut_table[645] = 16'b0000011011001111; 
assign lut_table[646] = 16'b0000011011011101; 
assign lut_table[647] = 16'b0000011011011110; 
assign lut_table[648] = 16'b0000011011011111; 
assign lut_table[649] = 16'b0000011011101110; 
assign lut_table[650] = 16'b0000011011101111; 
assign lut_table[651] = 16'b0000011011111111; 
assign lut_table[652] = 16'b0000011101110111; 
assign lut_table[653] = 16'b0000011101111000; 
assign lut_table[654] = 16'b0000011101111001; 
assign lut_table[655] = 16'b0000011101111010; 
assign lut_table[656] = 16'b0000011101111011; 
assign lut_table[657] = 16'b0000011101111100; 
assign lut_table[658] = 16'b0000011101111101; 
assign lut_table[659] = 16'b0000011101111110; 
assign lut_table[660] = 16'b0000011101111111; 
assign lut_table[661] = 16'b0000011110001000; 
assign lut_table[662] = 16'b0000011110001001; 
assign lut_table[663] = 16'b0000011110001010; 
assign lut_table[664] = 16'b0000011110001011; 
assign lut_table[665] = 16'b0000011110001100; 
assign lut_table[666] = 16'b0000011110001101; 
assign lut_table[667] = 16'b0000011110001110; 
assign lut_table[668] = 16'b0000011110001111; 
assign lut_table[669] = 16'b0000011110011001; 
assign lut_table[670] = 16'b0000011110011010; 
assign lut_table[671] = 16'b0000011110011011; 
assign lut_table[672] = 16'b0000011110011100; 
assign lut_table[673] = 16'b0000011110011101; 
assign lut_table[674] = 16'b0000011110011110; 
assign lut_table[675] = 16'b0000011110011111; 
assign lut_table[676] = 16'b0000011110101010; 
assign lut_table[677] = 16'b0000011110101011; 
assign lut_table[678] = 16'b0000011110101100; 
assign lut_table[679] = 16'b0000011110101101; 
assign lut_table[680] = 16'b0000011110101110; 
assign lut_table[681] = 16'b0000011110101111; 
assign lut_table[682] = 16'b0000011110111011; 
assign lut_table[683] = 16'b0000011110111100; 
assign lut_table[684] = 16'b0000011110111101; 
assign lut_table[685] = 16'b0000011110111110; 
assign lut_table[686] = 16'b0000011110111111; 
assign lut_table[687] = 16'b0000011111001100; 
assign lut_table[688] = 16'b0000011111001101; 
assign lut_table[689] = 16'b0000011111001110; 
assign lut_table[690] = 16'b0000011111001111; 
assign lut_table[691] = 16'b0000011111011101; 
assign lut_table[692] = 16'b0000011111011110; 
assign lut_table[693] = 16'b0000011111011111; 
assign lut_table[694] = 16'b0000011111101110; 
assign lut_table[695] = 16'b0000011111101111; 
assign lut_table[696] = 16'b0000011111111111; 
assign lut_table[697] = 16'b0000100010001000; 
assign lut_table[698] = 16'b0000100010001001; 
assign lut_table[699] = 16'b0000100010001010; 
assign lut_table[700] = 16'b0000100010001011; 
assign lut_table[701] = 16'b0000100010001100; 
assign lut_table[702] = 16'b0000100010001101; 
assign lut_table[703] = 16'b0000100010001110; 
assign lut_table[704] = 16'b0000100010001111; 
assign lut_table[705] = 16'b0000100010011001; 
assign lut_table[706] = 16'b0000100010011010; 
assign lut_table[707] = 16'b0000100010011011; 
assign lut_table[708] = 16'b0000100010011100; 
assign lut_table[709] = 16'b0000100010011101; 
assign lut_table[710] = 16'b0000100010011110; 
assign lut_table[711] = 16'b0000100010011111; 
assign lut_table[712] = 16'b0000100010101010; 
assign lut_table[713] = 16'b0000100010101011; 
assign lut_table[714] = 16'b0000100010101100; 
assign lut_table[715] = 16'b0000100010101101; 
assign lut_table[716] = 16'b0000100010101110; 
assign lut_table[717] = 16'b0000100010101111; 
assign lut_table[718] = 16'b0000100010111011; 
assign lut_table[719] = 16'b0000100010111100; 
assign lut_table[720] = 16'b0000100010111101; 
assign lut_table[721] = 16'b0000100010111110; 
assign lut_table[722] = 16'b0000100010111111; 
assign lut_table[723] = 16'b0000100011001100; 
assign lut_table[724] = 16'b0000100011001101; 
assign lut_table[725] = 16'b0000100011001110; 
assign lut_table[726] = 16'b0000100011001111; 
assign lut_table[727] = 16'b0000100011011101; 
assign lut_table[728] = 16'b0000100011011110; 
assign lut_table[729] = 16'b0000100011011111; 
assign lut_table[730] = 16'b0000100011101110; 
assign lut_table[731] = 16'b0000100011101111; 
assign lut_table[732] = 16'b0000100011111111; 
assign lut_table[733] = 16'b0000100110011001; 
assign lut_table[734] = 16'b0000100110011010; 
assign lut_table[735] = 16'b0000100110011011; 
assign lut_table[736] = 16'b0000100110011100; 
assign lut_table[737] = 16'b0000100110011101; 
assign lut_table[738] = 16'b0000100110011110; 
assign lut_table[739] = 16'b0000100110011111; 
assign lut_table[740] = 16'b0000100110101010; 
assign lut_table[741] = 16'b0000100110101011; 
assign lut_table[742] = 16'b0000100110101100; 
assign lut_table[743] = 16'b0000100110101101; 
assign lut_table[744] = 16'b0000100110101110; 
assign lut_table[745] = 16'b0000100110101111; 
assign lut_table[746] = 16'b0000100110111011; 
assign lut_table[747] = 16'b0000100110111100; 
assign lut_table[748] = 16'b0000100110111101; 
assign lut_table[749] = 16'b0000100110111110; 
assign lut_table[750] = 16'b0000100110111111; 
assign lut_table[751] = 16'b0000100111001100; 
assign lut_table[752] = 16'b0000100111001101; 
assign lut_table[753] = 16'b0000100111001110; 
assign lut_table[754] = 16'b0000100111001111; 
assign lut_table[755] = 16'b0000100111011101; 
assign lut_table[756] = 16'b0000100111011110; 
assign lut_table[757] = 16'b0000100111011111; 
assign lut_table[758] = 16'b0000100111101110; 
assign lut_table[759] = 16'b0000100111101111; 
assign lut_table[760] = 16'b0000100111111111; 
assign lut_table[761] = 16'b0000101010101010; 
assign lut_table[762] = 16'b0000101010101011; 
assign lut_table[763] = 16'b0000101010101100; 
assign lut_table[764] = 16'b0000101010101101; 
assign lut_table[765] = 16'b0000101010101110; 
assign lut_table[766] = 16'b0000101010101111; 
assign lut_table[767] = 16'b0000101010111011; 
assign lut_table[768] = 16'b0000101010111100; 
assign lut_table[769] = 16'b0000101010111101; 
assign lut_table[770] = 16'b0000101010111110; 
assign lut_table[771] = 16'b0000101010111111; 
assign lut_table[772] = 16'b0000101011001100; 
assign lut_table[773] = 16'b0000101011001101; 
assign lut_table[774] = 16'b0000101011001110; 
assign lut_table[775] = 16'b0000101011001111; 
assign lut_table[776] = 16'b0000101011011101; 
assign lut_table[777] = 16'b0000101011011110; 
assign lut_table[778] = 16'b0000101011011111; 
assign lut_table[779] = 16'b0000101011101110; 
assign lut_table[780] = 16'b0000101011101111; 
assign lut_table[781] = 16'b0000101011111111; 
assign lut_table[782] = 16'b0000101110111011; 
assign lut_table[783] = 16'b0000101110111100; 
assign lut_table[784] = 16'b0000101110111101; 
assign lut_table[785] = 16'b0000101110111110; 
assign lut_table[786] = 16'b0000101110111111; 
assign lut_table[787] = 16'b0000101111001100; 
assign lut_table[788] = 16'b0000101111001101; 
assign lut_table[789] = 16'b0000101111001110; 
assign lut_table[790] = 16'b0000101111001111; 
assign lut_table[791] = 16'b0000101111011101; 
assign lut_table[792] = 16'b0000101111011110; 
assign lut_table[793] = 16'b0000101111011111; 
assign lut_table[794] = 16'b0000101111101110; 
assign lut_table[795] = 16'b0000101111101111; 
assign lut_table[796] = 16'b0000101111111111; 
assign lut_table[797] = 16'b0000110011001100; 
assign lut_table[798] = 16'b0000110011001101; 
assign lut_table[799] = 16'b0000110011001110; 
assign lut_table[800] = 16'b0000110011001111; 
assign lut_table[801] = 16'b0000110011011101; 
assign lut_table[802] = 16'b0000110011011110; 
assign lut_table[803] = 16'b0000110011011111; 
assign lut_table[804] = 16'b0000110011101110; 
assign lut_table[805] = 16'b0000110011101111; 
assign lut_table[806] = 16'b0000110011111111; 
assign lut_table[807] = 16'b0000110111011101; 
assign lut_table[808] = 16'b0000110111011110; 
assign lut_table[809] = 16'b0000110111011111; 
assign lut_table[810] = 16'b0000110111101110; 
assign lut_table[811] = 16'b0000110111101111; 
assign lut_table[812] = 16'b0000110111111111; 
assign lut_table[813] = 16'b0000111011101110; 
assign lut_table[814] = 16'b0000111011101111; 
assign lut_table[815] = 16'b0000111011111111; 
assign lut_table[816] = 16'b0000111111111111; 
assign lut_table[817] = 16'b0001000100010001; 
assign lut_table[818] = 16'b0001000100010010; 
assign lut_table[819] = 16'b0001000100010011; 
assign lut_table[820] = 16'b0001000100010100; 
assign lut_table[821] = 16'b0001000100010101; 
assign lut_table[822] = 16'b0001000100010110; 
assign lut_table[823] = 16'b0001000100010111; 
assign lut_table[824] = 16'b0001000100011000; 
assign lut_table[825] = 16'b0001000100011001; 
assign lut_table[826] = 16'b0001000100011010; 
assign lut_table[827] = 16'b0001000100011011; 
assign lut_table[828] = 16'b0001000100011100; 
assign lut_table[829] = 16'b0001000100011101; 
assign lut_table[830] = 16'b0001000100011110; 
assign lut_table[831] = 16'b0001000100011111; 
assign lut_table[832] = 16'b0001000100100010; 
assign lut_table[833] = 16'b0001000100100011; 
assign lut_table[834] = 16'b0001000100100100; 
assign lut_table[835] = 16'b0001000100100101; 
assign lut_table[836] = 16'b0001000100100110; 
assign lut_table[837] = 16'b0001000100100111; 
assign lut_table[838] = 16'b0001000100101000; 
assign lut_table[839] = 16'b0001000100101001; 
assign lut_table[840] = 16'b0001000100101010; 
assign lut_table[841] = 16'b0001000100101011; 
assign lut_table[842] = 16'b0001000100101100; 
assign lut_table[843] = 16'b0001000100101101; 
assign lut_table[844] = 16'b0001000100101110; 
assign lut_table[845] = 16'b0001000100101111; 
assign lut_table[846] = 16'b0001000100110011; 
assign lut_table[847] = 16'b0001000100110100; 
assign lut_table[848] = 16'b0001000100110101; 
assign lut_table[849] = 16'b0001000100110110; 
assign lut_table[850] = 16'b0001000100110111; 
assign lut_table[851] = 16'b0001000100111000; 
assign lut_table[852] = 16'b0001000100111001; 
assign lut_table[853] = 16'b0001000100111010; 
assign lut_table[854] = 16'b0001000100111011; 
assign lut_table[855] = 16'b0001000100111100; 
assign lut_table[856] = 16'b0001000100111101; 
assign lut_table[857] = 16'b0001000100111110; 
assign lut_table[858] = 16'b0001000100111111; 
assign lut_table[859] = 16'b0001000101000100; 
assign lut_table[860] = 16'b0001000101000101; 
assign lut_table[861] = 16'b0001000101000110; 
assign lut_table[862] = 16'b0001000101000111; 
assign lut_table[863] = 16'b0001000101001000; 
assign lut_table[864] = 16'b0001000101001001; 
assign lut_table[865] = 16'b0001000101001010; 
assign lut_table[866] = 16'b0001000101001011; 
assign lut_table[867] = 16'b0001000101001100; 
assign lut_table[868] = 16'b0001000101001101; 
assign lut_table[869] = 16'b0001000101001110; 
assign lut_table[870] = 16'b0001000101001111; 
assign lut_table[871] = 16'b0001000101010101; 
assign lut_table[872] = 16'b0001000101010110; 
assign lut_table[873] = 16'b0001000101010111; 
assign lut_table[874] = 16'b0001000101011000; 
assign lut_table[875] = 16'b0001000101011001; 
assign lut_table[876] = 16'b0001000101011010; 
assign lut_table[877] = 16'b0001000101011011; 
assign lut_table[878] = 16'b0001000101011100; 
assign lut_table[879] = 16'b0001000101011101; 
assign lut_table[880] = 16'b0001000101011110; 
assign lut_table[881] = 16'b0001000101011111; 
assign lut_table[882] = 16'b0001000101100110; 
assign lut_table[883] = 16'b0001000101100111; 
assign lut_table[884] = 16'b0001000101101000; 
assign lut_table[885] = 16'b0001000101101001; 
assign lut_table[886] = 16'b0001000101101010; 
assign lut_table[887] = 16'b0001000101101011; 
assign lut_table[888] = 16'b0001000101101100; 
assign lut_table[889] = 16'b0001000101101101; 
assign lut_table[890] = 16'b0001000101101110; 
assign lut_table[891] = 16'b0001000101101111; 
assign lut_table[892] = 16'b0001000101110111; 
assign lut_table[893] = 16'b0001000101111000; 
assign lut_table[894] = 16'b0001000101111001; 
assign lut_table[895] = 16'b0001000101111010; 
assign lut_table[896] = 16'b0001000101111011; 
assign lut_table[897] = 16'b0001000101111100; 
assign lut_table[898] = 16'b0001000101111101; 
assign lut_table[899] = 16'b0001000101111110; 
assign lut_table[900] = 16'b0001000101111111; 
assign lut_table[901] = 16'b0001000110001000; 
assign lut_table[902] = 16'b0001000110001001; 
assign lut_table[903] = 16'b0001000110001010; 
assign lut_table[904] = 16'b0001000110001011; 
assign lut_table[905] = 16'b0001000110001100; 
assign lut_table[906] = 16'b0001000110001101; 
assign lut_table[907] = 16'b0001000110001110; 
assign lut_table[908] = 16'b0001000110001111; 
assign lut_table[909] = 16'b0001000110011001; 
assign lut_table[910] = 16'b0001000110011010; 
assign lut_table[911] = 16'b0001000110011011; 
assign lut_table[912] = 16'b0001000110011100; 
assign lut_table[913] = 16'b0001000110011101; 
assign lut_table[914] = 16'b0001000110011110; 
assign lut_table[915] = 16'b0001000110011111; 
assign lut_table[916] = 16'b0001000110101010; 
assign lut_table[917] = 16'b0001000110101011; 
assign lut_table[918] = 16'b0001000110101100; 
assign lut_table[919] = 16'b0001000110101101; 
assign lut_table[920] = 16'b0001000110101110; 
assign lut_table[921] = 16'b0001000110101111; 
assign lut_table[922] = 16'b0001000110111011; 
assign lut_table[923] = 16'b0001000110111100; 
assign lut_table[924] = 16'b0001000110111101; 
assign lut_table[925] = 16'b0001000110111110; 
assign lut_table[926] = 16'b0001000110111111; 
assign lut_table[927] = 16'b0001000111001100; 
assign lut_table[928] = 16'b0001000111001101; 
assign lut_table[929] = 16'b0001000111001110; 
assign lut_table[930] = 16'b0001000111001111; 
assign lut_table[931] = 16'b0001000111011101; 
assign lut_table[932] = 16'b0001000111011110; 
assign lut_table[933] = 16'b0001000111011111; 
assign lut_table[934] = 16'b0001000111101110; 
assign lut_table[935] = 16'b0001000111101111; 
assign lut_table[936] = 16'b0001000111111111; 
assign lut_table[937] = 16'b0001001000100010; 
assign lut_table[938] = 16'b0001001000100011; 
assign lut_table[939] = 16'b0001001000100100; 
assign lut_table[940] = 16'b0001001000100101; 
assign lut_table[941] = 16'b0001001000100110; 
assign lut_table[942] = 16'b0001001000100111; 
assign lut_table[943] = 16'b0001001000101000; 
assign lut_table[944] = 16'b0001001000101001; 
assign lut_table[945] = 16'b0001001000101010; 
assign lut_table[946] = 16'b0001001000101011; 
assign lut_table[947] = 16'b0001001000101100; 
assign lut_table[948] = 16'b0001001000101101; 
assign lut_table[949] = 16'b0001001000101110; 
assign lut_table[950] = 16'b0001001000101111; 
assign lut_table[951] = 16'b0001001000110011; 
assign lut_table[952] = 16'b0001001000110100; 
assign lut_table[953] = 16'b0001001000110101; 
assign lut_table[954] = 16'b0001001000110110; 
assign lut_table[955] = 16'b0001001000110111; 
assign lut_table[956] = 16'b0001001000111000; 
assign lut_table[957] = 16'b0001001000111001; 
assign lut_table[958] = 16'b0001001000111010; 
assign lut_table[959] = 16'b0001001000111011; 
assign lut_table[960] = 16'b0001001000111100; 
assign lut_table[961] = 16'b0001001000111101; 
assign lut_table[962] = 16'b0001001000111110; 
assign lut_table[963] = 16'b0001001000111111; 
assign lut_table[964] = 16'b0001001001000100; 
assign lut_table[965] = 16'b0001001001000101; 
assign lut_table[966] = 16'b0001001001000110; 
assign lut_table[967] = 16'b0001001001000111; 
assign lut_table[968] = 16'b0001001001001000; 
assign lut_table[969] = 16'b0001001001001001; 
assign lut_table[970] = 16'b0001001001001010; 
assign lut_table[971] = 16'b0001001001001011; 
assign lut_table[972] = 16'b0001001001001100; 
assign lut_table[973] = 16'b0001001001001101; 
assign lut_table[974] = 16'b0001001001001110; 
assign lut_table[975] = 16'b0001001001001111; 
assign lut_table[976] = 16'b0001001001010101; 
assign lut_table[977] = 16'b0001001001010110; 
assign lut_table[978] = 16'b0001001001010111; 
assign lut_table[979] = 16'b0001001001011000; 
assign lut_table[980] = 16'b0001001001011001; 
assign lut_table[981] = 16'b0001001001011010; 
assign lut_table[982] = 16'b0001001001011011; 
assign lut_table[983] = 16'b0001001001011100; 
assign lut_table[984] = 16'b0001001001011101; 
assign lut_table[985] = 16'b0001001001011110; 
assign lut_table[986] = 16'b0001001001011111; 
assign lut_table[987] = 16'b0001001001100110; 
assign lut_table[988] = 16'b0001001001100111; 
assign lut_table[989] = 16'b0001001001101000; 
assign lut_table[990] = 16'b0001001001101001; 
assign lut_table[991] = 16'b0001001001101010; 
assign lut_table[992] = 16'b0001001001101011; 
assign lut_table[993] = 16'b0001001001101100; 
assign lut_table[994] = 16'b0001001001101101; 
assign lut_table[995] = 16'b0001001001101110; 
assign lut_table[996] = 16'b0001001001101111; 
assign lut_table[997] = 16'b0001001001110111; 
assign lut_table[998] = 16'b0001001001111000; 
assign lut_table[999] = 16'b0001001001111001; 
assign lut_table[1000] = 16'b0001001001111010; 
assign lut_table[1001] = 16'b0001001001111011; 
assign lut_table[1002] = 16'b0001001001111100; 
assign lut_table[1003] = 16'b0001001001111101; 
assign lut_table[1004] = 16'b0001001001111110; 
assign lut_table[1005] = 16'b0001001001111111; 
assign lut_table[1006] = 16'b0001001010001000; 
assign lut_table[1007] = 16'b0001001010001001; 
assign lut_table[1008] = 16'b0001001010001010; 
assign lut_table[1009] = 16'b0001001010001011; 
assign lut_table[1010] = 16'b0001001010001100; 
assign lut_table[1011] = 16'b0001001010001101; 
assign lut_table[1012] = 16'b0001001010001110; 
assign lut_table[1013] = 16'b0001001010001111; 
assign lut_table[1014] = 16'b0001001010011001; 
assign lut_table[1015] = 16'b0001001010011010; 
assign lut_table[1016] = 16'b0001001010011011; 
assign lut_table[1017] = 16'b0001001010011100; 
assign lut_table[1018] = 16'b0001001010011101; 
assign lut_table[1019] = 16'b0001001010011110; 
assign lut_table[1020] = 16'b0001001010011111; 
assign lut_table[1021] = 16'b0001001010101010; 
assign lut_table[1022] = 16'b0001001010101011; 
assign lut_table[1023] = 16'b0001001010101100; 
assign lut_table[1024] = 16'b0001001010101101; 
assign lut_table[1025] = 16'b0001001010101110; 
assign lut_table[1026] = 16'b0001001010101111; 
assign lut_table[1027] = 16'b0001001010111011; 
assign lut_table[1028] = 16'b0001001010111100; 
assign lut_table[1029] = 16'b0001001010111101; 
assign lut_table[1030] = 16'b0001001010111110; 
assign lut_table[1031] = 16'b0001001010111111; 
assign lut_table[1032] = 16'b0001001011001100; 
assign lut_table[1033] = 16'b0001001011001101; 
assign lut_table[1034] = 16'b0001001011001110; 
assign lut_table[1035] = 16'b0001001011001111; 
assign lut_table[1036] = 16'b0001001011011101; 
assign lut_table[1037] = 16'b0001001011011110; 
assign lut_table[1038] = 16'b0001001011011111; 
assign lut_table[1039] = 16'b0001001011101110; 
assign lut_table[1040] = 16'b0001001011101111; 
assign lut_table[1041] = 16'b0001001011111111; 
assign lut_table[1042] = 16'b0001001100110011; 
assign lut_table[1043] = 16'b0001001100110100; 
assign lut_table[1044] = 16'b0001001100110101; 
assign lut_table[1045] = 16'b0001001100110110; 
assign lut_table[1046] = 16'b0001001100110111; 
assign lut_table[1047] = 16'b0001001100111000; 
assign lut_table[1048] = 16'b0001001100111001; 
assign lut_table[1049] = 16'b0001001100111010; 
assign lut_table[1050] = 16'b0001001100111011; 
assign lut_table[1051] = 16'b0001001100111100; 
assign lut_table[1052] = 16'b0001001100111101; 
assign lut_table[1053] = 16'b0001001100111110; 
assign lut_table[1054] = 16'b0001001100111111; 
assign lut_table[1055] = 16'b0001001101000100; 
assign lut_table[1056] = 16'b0001001101000101; 
assign lut_table[1057] = 16'b0001001101000110; 
assign lut_table[1058] = 16'b0001001101000111; 
assign lut_table[1059] = 16'b0001001101001000; 
assign lut_table[1060] = 16'b0001001101001001; 
assign lut_table[1061] = 16'b0001001101001010; 
assign lut_table[1062] = 16'b0001001101001011; 
assign lut_table[1063] = 16'b0001001101001100; 
assign lut_table[1064] = 16'b0001001101001101; 
assign lut_table[1065] = 16'b0001001101001110; 
assign lut_table[1066] = 16'b0001001101001111; 
assign lut_table[1067] = 16'b0001001101010101; 
assign lut_table[1068] = 16'b0001001101010110; 
assign lut_table[1069] = 16'b0001001101010111; 
assign lut_table[1070] = 16'b0001001101011000; 
assign lut_table[1071] = 16'b0001001101011001; 
assign lut_table[1072] = 16'b0001001101011010; 
assign lut_table[1073] = 16'b0001001101011011; 
assign lut_table[1074] = 16'b0001001101011100; 
assign lut_table[1075] = 16'b0001001101011101; 
assign lut_table[1076] = 16'b0001001101011110; 
assign lut_table[1077] = 16'b0001001101011111; 
assign lut_table[1078] = 16'b0001001101100110; 
assign lut_table[1079] = 16'b0001001101100111; 
assign lut_table[1080] = 16'b0001001101101000; 
assign lut_table[1081] = 16'b0001001101101001; 
assign lut_table[1082] = 16'b0001001101101010; 
assign lut_table[1083] = 16'b0001001101101011; 
assign lut_table[1084] = 16'b0001001101101100; 
assign lut_table[1085] = 16'b0001001101101101; 
assign lut_table[1086] = 16'b0001001101101110; 
assign lut_table[1087] = 16'b0001001101101111; 
assign lut_table[1088] = 16'b0001001101110111; 
assign lut_table[1089] = 16'b0001001101111000; 
assign lut_table[1090] = 16'b0001001101111001; 
assign lut_table[1091] = 16'b0001001101111010; 
assign lut_table[1092] = 16'b0001001101111011; 
assign lut_table[1093] = 16'b0001001101111100; 
assign lut_table[1094] = 16'b0001001101111101; 
assign lut_table[1095] = 16'b0001001101111110; 
assign lut_table[1096] = 16'b0001001101111111; 
assign lut_table[1097] = 16'b0001001110001000; 
assign lut_table[1098] = 16'b0001001110001001; 
assign lut_table[1099] = 16'b0001001110001010; 
assign lut_table[1100] = 16'b0001001110001011; 
assign lut_table[1101] = 16'b0001001110001100; 
assign lut_table[1102] = 16'b0001001110001101; 
assign lut_table[1103] = 16'b0001001110001110; 
assign lut_table[1104] = 16'b0001001110001111; 
assign lut_table[1105] = 16'b0001001110011001; 
assign lut_table[1106] = 16'b0001001110011010; 
assign lut_table[1107] = 16'b0001001110011011; 
assign lut_table[1108] = 16'b0001001110011100; 
assign lut_table[1109] = 16'b0001001110011101; 
assign lut_table[1110] = 16'b0001001110011110; 
assign lut_table[1111] = 16'b0001001110011111; 
assign lut_table[1112] = 16'b0001001110101010; 
assign lut_table[1113] = 16'b0001001110101011; 
assign lut_table[1114] = 16'b0001001110101100; 
assign lut_table[1115] = 16'b0001001110101101; 
assign lut_table[1116] = 16'b0001001110101110; 
assign lut_table[1117] = 16'b0001001110101111; 
assign lut_table[1118] = 16'b0001001110111011; 
assign lut_table[1119] = 16'b0001001110111100; 
assign lut_table[1120] = 16'b0001001110111101; 
assign lut_table[1121] = 16'b0001001110111110; 
assign lut_table[1122] = 16'b0001001110111111; 
assign lut_table[1123] = 16'b0001001111001100; 
assign lut_table[1124] = 16'b0001001111001101; 
assign lut_table[1125] = 16'b0001001111001110; 
assign lut_table[1126] = 16'b0001001111001111; 
assign lut_table[1127] = 16'b0001001111011101; 
assign lut_table[1128] = 16'b0001001111011110; 
assign lut_table[1129] = 16'b0001001111011111; 
assign lut_table[1130] = 16'b0001001111101110; 
assign lut_table[1131] = 16'b0001001111101111; 
assign lut_table[1132] = 16'b0001001111111111; 
assign lut_table[1133] = 16'b0001010001000100; 
assign lut_table[1134] = 16'b0001010001000101; 
assign lut_table[1135] = 16'b0001010001000110; 
assign lut_table[1136] = 16'b0001010001000111; 
assign lut_table[1137] = 16'b0001010001001000; 
assign lut_table[1138] = 16'b0001010001001001; 
assign lut_table[1139] = 16'b0001010001001010; 
assign lut_table[1140] = 16'b0001010001001011; 
assign lut_table[1141] = 16'b0001010001001100; 
assign lut_table[1142] = 16'b0001010001001101; 
assign lut_table[1143] = 16'b0001010001001110; 
assign lut_table[1144] = 16'b0001010001001111; 
assign lut_table[1145] = 16'b0001010001010101; 
assign lut_table[1146] = 16'b0001010001010110; 
assign lut_table[1147] = 16'b0001010001010111; 
assign lut_table[1148] = 16'b0001010001011000; 
assign lut_table[1149] = 16'b0001010001011001; 
assign lut_table[1150] = 16'b0001010001011010; 
assign lut_table[1151] = 16'b0001010001011011; 
assign lut_table[1152] = 16'b0001010001011100; 
assign lut_table[1153] = 16'b0001010001011101; 
assign lut_table[1154] = 16'b0001010001011110; 
assign lut_table[1155] = 16'b0001010001011111; 
assign lut_table[1156] = 16'b0001010001100110; 
assign lut_table[1157] = 16'b0001010001100111; 
assign lut_table[1158] = 16'b0001010001101000; 
assign lut_table[1159] = 16'b0001010001101001; 
assign lut_table[1160] = 16'b0001010001101010; 
assign lut_table[1161] = 16'b0001010001101011; 
assign lut_table[1162] = 16'b0001010001101100; 
assign lut_table[1163] = 16'b0001010001101101; 
assign lut_table[1164] = 16'b0001010001101110; 
assign lut_table[1165] = 16'b0001010001101111; 
assign lut_table[1166] = 16'b0001010001110111; 
assign lut_table[1167] = 16'b0001010001111000; 
assign lut_table[1168] = 16'b0001010001111001; 
assign lut_table[1169] = 16'b0001010001111010; 
assign lut_table[1170] = 16'b0001010001111011; 
assign lut_table[1171] = 16'b0001010001111100; 
assign lut_table[1172] = 16'b0001010001111101; 
assign lut_table[1173] = 16'b0001010001111110; 
assign lut_table[1174] = 16'b0001010001111111; 
assign lut_table[1175] = 16'b0001010010001000; 
assign lut_table[1176] = 16'b0001010010001001; 
assign lut_table[1177] = 16'b0001010010001010; 
assign lut_table[1178] = 16'b0001010010001011; 
assign lut_table[1179] = 16'b0001010010001100; 
assign lut_table[1180] = 16'b0001010010001101; 
assign lut_table[1181] = 16'b0001010010001110; 
assign lut_table[1182] = 16'b0001010010001111; 
assign lut_table[1183] = 16'b0001010010011001; 
assign lut_table[1184] = 16'b0001010010011010; 
assign lut_table[1185] = 16'b0001010010011011; 
assign lut_table[1186] = 16'b0001010010011100; 
assign lut_table[1187] = 16'b0001010010011101; 
assign lut_table[1188] = 16'b0001010010011110; 
assign lut_table[1189] = 16'b0001010010011111; 
assign lut_table[1190] = 16'b0001010010101010; 
assign lut_table[1191] = 16'b0001010010101011; 
assign lut_table[1192] = 16'b0001010010101100; 
assign lut_table[1193] = 16'b0001010010101101; 
assign lut_table[1194] = 16'b0001010010101110; 
assign lut_table[1195] = 16'b0001010010101111; 
assign lut_table[1196] = 16'b0001010010111011; 
assign lut_table[1197] = 16'b0001010010111100; 
assign lut_table[1198] = 16'b0001010010111101; 
assign lut_table[1199] = 16'b0001010010111110; 
assign lut_table[1200] = 16'b0001010010111111; 
assign lut_table[1201] = 16'b0001010011001100; 
assign lut_table[1202] = 16'b0001010011001101; 
assign lut_table[1203] = 16'b0001010011001110; 
assign lut_table[1204] = 16'b0001010011001111; 
assign lut_table[1205] = 16'b0001010011011101; 
assign lut_table[1206] = 16'b0001010011011110; 
assign lut_table[1207] = 16'b0001010011011111; 
assign lut_table[1208] = 16'b0001010011101110; 
assign lut_table[1209] = 16'b0001010011101111; 
assign lut_table[1210] = 16'b0001010011111111; 
assign lut_table[1211] = 16'b0001010101010101; 
assign lut_table[1212] = 16'b0001010101010110; 
assign lut_table[1213] = 16'b0001010101010111; 
assign lut_table[1214] = 16'b0001010101011000; 
assign lut_table[1215] = 16'b0001010101011001; 
assign lut_table[1216] = 16'b0001010101011010; 
assign lut_table[1217] = 16'b0001010101011011; 
assign lut_table[1218] = 16'b0001010101011100; 
assign lut_table[1219] = 16'b0001010101011101; 
assign lut_table[1220] = 16'b0001010101011110; 
assign lut_table[1221] = 16'b0001010101011111; 
assign lut_table[1222] = 16'b0001010101100110; 
assign lut_table[1223] = 16'b0001010101100111; 
assign lut_table[1224] = 16'b0001010101101000; 
assign lut_table[1225] = 16'b0001010101101001; 
assign lut_table[1226] = 16'b0001010101101010; 
assign lut_table[1227] = 16'b0001010101101011; 
assign lut_table[1228] = 16'b0001010101101100; 
assign lut_table[1229] = 16'b0001010101101101; 
assign lut_table[1230] = 16'b0001010101101110; 
assign lut_table[1231] = 16'b0001010101101111; 
assign lut_table[1232] = 16'b0001010101110111; 
assign lut_table[1233] = 16'b0001010101111000; 
assign lut_table[1234] = 16'b0001010101111001; 
assign lut_table[1235] = 16'b0001010101111010; 
assign lut_table[1236] = 16'b0001010101111011; 
assign lut_table[1237] = 16'b0001010101111100; 
assign lut_table[1238] = 16'b0001010101111101; 
assign lut_table[1239] = 16'b0001010101111110; 
assign lut_table[1240] = 16'b0001010101111111; 
assign lut_table[1241] = 16'b0001010110001000; 
assign lut_table[1242] = 16'b0001010110001001; 
assign lut_table[1243] = 16'b0001010110001010; 
assign lut_table[1244] = 16'b0001010110001011; 
assign lut_table[1245] = 16'b0001010110001100; 
assign lut_table[1246] = 16'b0001010110001101; 
assign lut_table[1247] = 16'b0001010110001110; 
assign lut_table[1248] = 16'b0001010110001111; 
assign lut_table[1249] = 16'b0001010110011001; 
assign lut_table[1250] = 16'b0001010110011010; 
assign lut_table[1251] = 16'b0001010110011011; 
assign lut_table[1252] = 16'b0001010110011100; 
assign lut_table[1253] = 16'b0001010110011101; 
assign lut_table[1254] = 16'b0001010110011110; 
assign lut_table[1255] = 16'b0001010110011111; 
assign lut_table[1256] = 16'b0001010110101010; 
assign lut_table[1257] = 16'b0001010110101011; 
assign lut_table[1258] = 16'b0001010110101100; 
assign lut_table[1259] = 16'b0001010110101101; 
assign lut_table[1260] = 16'b0001010110101110; 
assign lut_table[1261] = 16'b0001010110101111; 
assign lut_table[1262] = 16'b0001010110111011; 
assign lut_table[1263] = 16'b0001010110111100; 
assign lut_table[1264] = 16'b0001010110111101; 
assign lut_table[1265] = 16'b0001010110111110; 
assign lut_table[1266] = 16'b0001010110111111; 
assign lut_table[1267] = 16'b0001010111001100; 
assign lut_table[1268] = 16'b0001010111001101; 
assign lut_table[1269] = 16'b0001010111001110; 
assign lut_table[1270] = 16'b0001010111001111; 
assign lut_table[1271] = 16'b0001010111011101; 
assign lut_table[1272] = 16'b0001010111011110; 
assign lut_table[1273] = 16'b0001010111011111; 
assign lut_table[1274] = 16'b0001010111101110; 
assign lut_table[1275] = 16'b0001010111101111; 
assign lut_table[1276] = 16'b0001010111111111; 
assign lut_table[1277] = 16'b0001011001100110; 
assign lut_table[1278] = 16'b0001011001100111; 
assign lut_table[1279] = 16'b0001011001101000; 
assign lut_table[1280] = 16'b0001011001101001; 
assign lut_table[1281] = 16'b0001011001101010; 
assign lut_table[1282] = 16'b0001011001101011; 
assign lut_table[1283] = 16'b0001011001101100; 
assign lut_table[1284] = 16'b0001011001101101; 
assign lut_table[1285] = 16'b0001011001101110; 
assign lut_table[1286] = 16'b0001011001101111; 
assign lut_table[1287] = 16'b0001011001110111; 
assign lut_table[1288] = 16'b0001011001111000; 
assign lut_table[1289] = 16'b0001011001111001; 
assign lut_table[1290] = 16'b0001011001111010; 
assign lut_table[1291] = 16'b0001011001111011; 
assign lut_table[1292] = 16'b0001011001111100; 
assign lut_table[1293] = 16'b0001011001111101; 
assign lut_table[1294] = 16'b0001011001111110; 
assign lut_table[1295] = 16'b0001011001111111; 
assign lut_table[1296] = 16'b0001011010001000; 
assign lut_table[1297] = 16'b0001011010001001; 
assign lut_table[1298] = 16'b0001011010001010; 
assign lut_table[1299] = 16'b0001011010001011; 
assign lut_table[1300] = 16'b0001011010001100; 
assign lut_table[1301] = 16'b0001011010001101; 
assign lut_table[1302] = 16'b0001011010001110; 
assign lut_table[1303] = 16'b0001011010001111; 
assign lut_table[1304] = 16'b0001011010011001; 
assign lut_table[1305] = 16'b0001011010011010; 
assign lut_table[1306] = 16'b0001011010011011; 
assign lut_table[1307] = 16'b0001011010011100; 
assign lut_table[1308] = 16'b0001011010011101; 
assign lut_table[1309] = 16'b0001011010011110; 
assign lut_table[1310] = 16'b0001011010011111; 
assign lut_table[1311] = 16'b0001011010101010; 
assign lut_table[1312] = 16'b0001011010101011; 
assign lut_table[1313] = 16'b0001011010101100; 
assign lut_table[1314] = 16'b0001011010101101; 
assign lut_table[1315] = 16'b0001011010101110; 
assign lut_table[1316] = 16'b0001011010101111; 
assign lut_table[1317] = 16'b0001011010111011; 
assign lut_table[1318] = 16'b0001011010111100; 
assign lut_table[1319] = 16'b0001011010111101; 
assign lut_table[1320] = 16'b0001011010111110; 
assign lut_table[1321] = 16'b0001011010111111; 
assign lut_table[1322] = 16'b0001011011001100; 
assign lut_table[1323] = 16'b0001011011001101; 
assign lut_table[1324] = 16'b0001011011001110; 
assign lut_table[1325] = 16'b0001011011001111; 
assign lut_table[1326] = 16'b0001011011011101; 
assign lut_table[1327] = 16'b0001011011011110; 
assign lut_table[1328] = 16'b0001011011011111; 
assign lut_table[1329] = 16'b0001011011101110; 
assign lut_table[1330] = 16'b0001011011101111; 
assign lut_table[1331] = 16'b0001011011111111; 
assign lut_table[1332] = 16'b0001011101110111; 
assign lut_table[1333] = 16'b0001011101111000; 
assign lut_table[1334] = 16'b0001011101111001; 
assign lut_table[1335] = 16'b0001011101111010; 
assign lut_table[1336] = 16'b0001011101111011; 
assign lut_table[1337] = 16'b0001011101111100; 
assign lut_table[1338] = 16'b0001011101111101; 
assign lut_table[1339] = 16'b0001011101111110; 
assign lut_table[1340] = 16'b0001011101111111; 
assign lut_table[1341] = 16'b0001011110001000; 
assign lut_table[1342] = 16'b0001011110001001; 
assign lut_table[1343] = 16'b0001011110001010; 
assign lut_table[1344] = 16'b0001011110001011; 
assign lut_table[1345] = 16'b0001011110001100; 
assign lut_table[1346] = 16'b0001011110001101; 
assign lut_table[1347] = 16'b0001011110001110; 
assign lut_table[1348] = 16'b0001011110001111; 
assign lut_table[1349] = 16'b0001011110011001; 
assign lut_table[1350] = 16'b0001011110011010; 
assign lut_table[1351] = 16'b0001011110011011; 
assign lut_table[1352] = 16'b0001011110011100; 
assign lut_table[1353] = 16'b0001011110011101; 
assign lut_table[1354] = 16'b0001011110011110; 
assign lut_table[1355] = 16'b0001011110011111; 
assign lut_table[1356] = 16'b0001011110101010; 
assign lut_table[1357] = 16'b0001011110101011; 
assign lut_table[1358] = 16'b0001011110101100; 
assign lut_table[1359] = 16'b0001011110101101; 
assign lut_table[1360] = 16'b0001011110101110; 
assign lut_table[1361] = 16'b0001011110101111; 
assign lut_table[1362] = 16'b0001011110111011; 
assign lut_table[1363] = 16'b0001011110111100; 
assign lut_table[1364] = 16'b0001011110111101; 
assign lut_table[1365] = 16'b0001011110111110; 
assign lut_table[1366] = 16'b0001011110111111; 
assign lut_table[1367] = 16'b0001011111001100; 
assign lut_table[1368] = 16'b0001011111001101; 
assign lut_table[1369] = 16'b0001011111001110; 
assign lut_table[1370] = 16'b0001011111001111; 
assign lut_table[1371] = 16'b0001011111011101; 
assign lut_table[1372] = 16'b0001011111011110; 
assign lut_table[1373] = 16'b0001011111011111; 
assign lut_table[1374] = 16'b0001011111101110; 
assign lut_table[1375] = 16'b0001011111101111; 
assign lut_table[1376] = 16'b0001011111111111; 
assign lut_table[1377] = 16'b0001100010001000; 
assign lut_table[1378] = 16'b0001100010001001; 
assign lut_table[1379] = 16'b0001100010001010; 
assign lut_table[1380] = 16'b0001100010001011; 
assign lut_table[1381] = 16'b0001100010001100; 
assign lut_table[1382] = 16'b0001100010001101; 
assign lut_table[1383] = 16'b0001100010001110; 
assign lut_table[1384] = 16'b0001100010001111; 
assign lut_table[1385] = 16'b0001100010011001; 
assign lut_table[1386] = 16'b0001100010011010; 
assign lut_table[1387] = 16'b0001100010011011; 
assign lut_table[1388] = 16'b0001100010011100; 
assign lut_table[1389] = 16'b0001100010011101; 
assign lut_table[1390] = 16'b0001100010011110; 
assign lut_table[1391] = 16'b0001100010011111; 
assign lut_table[1392] = 16'b0001100010101010; 
assign lut_table[1393] = 16'b0001100010101011; 
assign lut_table[1394] = 16'b0001100010101100; 
assign lut_table[1395] = 16'b0001100010101101; 
assign lut_table[1396] = 16'b0001100010101110; 
assign lut_table[1397] = 16'b0001100010101111; 
assign lut_table[1398] = 16'b0001100010111011; 
assign lut_table[1399] = 16'b0001100010111100; 
assign lut_table[1400] = 16'b0001100010111101; 
assign lut_table[1401] = 16'b0001100010111110; 
assign lut_table[1402] = 16'b0001100010111111; 
assign lut_table[1403] = 16'b0001100011001100; 
assign lut_table[1404] = 16'b0001100011001101; 
assign lut_table[1405] = 16'b0001100011001110; 
assign lut_table[1406] = 16'b0001100011001111; 
assign lut_table[1407] = 16'b0001100011011101; 
assign lut_table[1408] = 16'b0001100011011110; 
assign lut_table[1409] = 16'b0001100011011111; 
assign lut_table[1410] = 16'b0001100011101110; 
assign lut_table[1411] = 16'b0001100011101111; 
assign lut_table[1412] = 16'b0001100011111111; 
assign lut_table[1413] = 16'b0001100110011001; 
assign lut_table[1414] = 16'b0001100110011010; 
assign lut_table[1415] = 16'b0001100110011011; 
assign lut_table[1416] = 16'b0001100110011100; 
assign lut_table[1417] = 16'b0001100110011101; 
assign lut_table[1418] = 16'b0001100110011110; 
assign lut_table[1419] = 16'b0001100110011111; 
assign lut_table[1420] = 16'b0001100110101010; 
assign lut_table[1421] = 16'b0001100110101011; 
assign lut_table[1422] = 16'b0001100110101100; 
assign lut_table[1423] = 16'b0001100110101101; 
assign lut_table[1424] = 16'b0001100110101110; 
assign lut_table[1425] = 16'b0001100110101111; 
assign lut_table[1426] = 16'b0001100110111011; 
assign lut_table[1427] = 16'b0001100110111100; 
assign lut_table[1428] = 16'b0001100110111101; 
assign lut_table[1429] = 16'b0001100110111110; 
assign lut_table[1430] = 16'b0001100110111111; 
assign lut_table[1431] = 16'b0001100111001100; 
assign lut_table[1432] = 16'b0001100111001101; 
assign lut_table[1433] = 16'b0001100111001110; 
assign lut_table[1434] = 16'b0001100111001111; 
assign lut_table[1435] = 16'b0001100111011101; 
assign lut_table[1436] = 16'b0001100111011110; 
assign lut_table[1437] = 16'b0001100111011111; 
assign lut_table[1438] = 16'b0001100111101110; 
assign lut_table[1439] = 16'b0001100111101111; 
assign lut_table[1440] = 16'b0001100111111111; 
assign lut_table[1441] = 16'b0001101010101010; 
assign lut_table[1442] = 16'b0001101010101011; 
assign lut_table[1443] = 16'b0001101010101100; 
assign lut_table[1444] = 16'b0001101010101101; 
assign lut_table[1445] = 16'b0001101010101110; 
assign lut_table[1446] = 16'b0001101010101111; 
assign lut_table[1447] = 16'b0001101010111011; 
assign lut_table[1448] = 16'b0001101010111100; 
assign lut_table[1449] = 16'b0001101010111101; 
assign lut_table[1450] = 16'b0001101010111110; 
assign lut_table[1451] = 16'b0001101010111111; 
assign lut_table[1452] = 16'b0001101011001100; 
assign lut_table[1453] = 16'b0001101011001101; 
assign lut_table[1454] = 16'b0001101011001110; 
assign lut_table[1455] = 16'b0001101011001111; 
assign lut_table[1456] = 16'b0001101011011101; 
assign lut_table[1457] = 16'b0001101011011110; 
assign lut_table[1458] = 16'b0001101011011111; 
assign lut_table[1459] = 16'b0001101011101110; 
assign lut_table[1460] = 16'b0001101011101111; 
assign lut_table[1461] = 16'b0001101011111111; 
assign lut_table[1462] = 16'b0001101110111011; 
assign lut_table[1463] = 16'b0001101110111100; 
assign lut_table[1464] = 16'b0001101110111101; 
assign lut_table[1465] = 16'b0001101110111110; 
assign lut_table[1466] = 16'b0001101110111111; 
assign lut_table[1467] = 16'b0001101111001100; 
assign lut_table[1468] = 16'b0001101111001101; 
assign lut_table[1469] = 16'b0001101111001110; 
assign lut_table[1470] = 16'b0001101111001111; 
assign lut_table[1471] = 16'b0001101111011101; 
assign lut_table[1472] = 16'b0001101111011110; 
assign lut_table[1473] = 16'b0001101111011111; 
assign lut_table[1474] = 16'b0001101111101110; 
assign lut_table[1475] = 16'b0001101111101111; 
assign lut_table[1476] = 16'b0001101111111111; 
assign lut_table[1477] = 16'b0001110011001100; 
assign lut_table[1478] = 16'b0001110011001101; 
assign lut_table[1479] = 16'b0001110011001110; 
assign lut_table[1480] = 16'b0001110011001111; 
assign lut_table[1481] = 16'b0001110011011101; 
assign lut_table[1482] = 16'b0001110011011110; 
assign lut_table[1483] = 16'b0001110011011111; 
assign lut_table[1484] = 16'b0001110011101110; 
assign lut_table[1485] = 16'b0001110011101111; 
assign lut_table[1486] = 16'b0001110011111111; 
assign lut_table[1487] = 16'b0001110111011101; 
assign lut_table[1488] = 16'b0001110111011110; 
assign lut_table[1489] = 16'b0001110111011111; 
assign lut_table[1490] = 16'b0001110111101110; 
assign lut_table[1491] = 16'b0001110111101111; 
assign lut_table[1492] = 16'b0001110111111111; 
assign lut_table[1493] = 16'b0001111011101110; 
assign lut_table[1494] = 16'b0001111011101111; 
assign lut_table[1495] = 16'b0001111011111111; 
assign lut_table[1496] = 16'b0001111111111111; 
assign lut_table[1497] = 16'b0010001000100010; 
assign lut_table[1498] = 16'b0010001000100011; 
assign lut_table[1499] = 16'b0010001000100100; 
assign lut_table[1500] = 16'b0010001000100101; 
assign lut_table[1501] = 16'b0010001000100110; 
assign lut_table[1502] = 16'b0010001000100111; 
assign lut_table[1503] = 16'b0010001000101000; 
assign lut_table[1504] = 16'b0010001000101001; 
assign lut_table[1505] = 16'b0010001000101010; 
assign lut_table[1506] = 16'b0010001000101011; 
assign lut_table[1507] = 16'b0010001000101100; 
assign lut_table[1508] = 16'b0010001000101101; 
assign lut_table[1509] = 16'b0010001000101110; 
assign lut_table[1510] = 16'b0010001000101111; 
assign lut_table[1511] = 16'b0010001000110011; 
assign lut_table[1512] = 16'b0010001000110100; 
assign lut_table[1513] = 16'b0010001000110101; 
assign lut_table[1514] = 16'b0010001000110110; 
assign lut_table[1515] = 16'b0010001000110111; 
assign lut_table[1516] = 16'b0010001000111000; 
assign lut_table[1517] = 16'b0010001000111001; 
assign lut_table[1518] = 16'b0010001000111010; 
assign lut_table[1519] = 16'b0010001000111011; 
assign lut_table[1520] = 16'b0010001000111100; 
assign lut_table[1521] = 16'b0010001000111101; 
assign lut_table[1522] = 16'b0010001000111110; 
assign lut_table[1523] = 16'b0010001000111111; 
assign lut_table[1524] = 16'b0010001001000100; 
assign lut_table[1525] = 16'b0010001001000101; 
assign lut_table[1526] = 16'b0010001001000110; 
assign lut_table[1527] = 16'b0010001001000111; 
assign lut_table[1528] = 16'b0010001001001000; 
assign lut_table[1529] = 16'b0010001001001001; 
assign lut_table[1530] = 16'b0010001001001010; 
assign lut_table[1531] = 16'b0010001001001011; 
assign lut_table[1532] = 16'b0010001001001100; 
assign lut_table[1533] = 16'b0010001001001101; 
assign lut_table[1534] = 16'b0010001001001110; 
assign lut_table[1535] = 16'b0010001001001111; 
assign lut_table[1536] = 16'b0010001001010101; 
assign lut_table[1537] = 16'b0010001001010110; 
assign lut_table[1538] = 16'b0010001001010111; 
assign lut_table[1539] = 16'b0010001001011000; 
assign lut_table[1540] = 16'b0010001001011001; 
assign lut_table[1541] = 16'b0010001001011010; 
assign lut_table[1542] = 16'b0010001001011011; 
assign lut_table[1543] = 16'b0010001001011100; 
assign lut_table[1544] = 16'b0010001001011101; 
assign lut_table[1545] = 16'b0010001001011110; 
assign lut_table[1546] = 16'b0010001001011111; 
assign lut_table[1547] = 16'b0010001001100110; 
assign lut_table[1548] = 16'b0010001001100111; 
assign lut_table[1549] = 16'b0010001001101000; 
assign lut_table[1550] = 16'b0010001001101001; 
assign lut_table[1551] = 16'b0010001001101010; 
assign lut_table[1552] = 16'b0010001001101011; 
assign lut_table[1553] = 16'b0010001001101100; 
assign lut_table[1554] = 16'b0010001001101101; 
assign lut_table[1555] = 16'b0010001001101110; 
assign lut_table[1556] = 16'b0010001001101111; 
assign lut_table[1557] = 16'b0010001001110111; 
assign lut_table[1558] = 16'b0010001001111000; 
assign lut_table[1559] = 16'b0010001001111001; 
assign lut_table[1560] = 16'b0010001001111010; 
assign lut_table[1561] = 16'b0010001001111011; 
assign lut_table[1562] = 16'b0010001001111100; 
assign lut_table[1563] = 16'b0010001001111101; 
assign lut_table[1564] = 16'b0010001001111110; 
assign lut_table[1565] = 16'b0010001001111111; 
assign lut_table[1566] = 16'b0010001010001000; 
assign lut_table[1567] = 16'b0010001010001001; 
assign lut_table[1568] = 16'b0010001010001010; 
assign lut_table[1569] = 16'b0010001010001011; 
assign lut_table[1570] = 16'b0010001010001100; 
assign lut_table[1571] = 16'b0010001010001101; 
assign lut_table[1572] = 16'b0010001010001110; 
assign lut_table[1573] = 16'b0010001010001111; 
assign lut_table[1574] = 16'b0010001010011001; 
assign lut_table[1575] = 16'b0010001010011010; 
assign lut_table[1576] = 16'b0010001010011011; 
assign lut_table[1577] = 16'b0010001010011100; 
assign lut_table[1578] = 16'b0010001010011101; 
assign lut_table[1579] = 16'b0010001010011110; 
assign lut_table[1580] = 16'b0010001010011111; 
assign lut_table[1581] = 16'b0010001010101010; 
assign lut_table[1582] = 16'b0010001010101011; 
assign lut_table[1583] = 16'b0010001010101100; 
assign lut_table[1584] = 16'b0010001010101101; 
assign lut_table[1585] = 16'b0010001010101110; 
assign lut_table[1586] = 16'b0010001010101111; 
assign lut_table[1587] = 16'b0010001010111011; 
assign lut_table[1588] = 16'b0010001010111100; 
assign lut_table[1589] = 16'b0010001010111101; 
assign lut_table[1590] = 16'b0010001010111110; 
assign lut_table[1591] = 16'b0010001010111111; 
assign lut_table[1592] = 16'b0010001011001100; 
assign lut_table[1593] = 16'b0010001011001101; 
assign lut_table[1594] = 16'b0010001011001110; 
assign lut_table[1595] = 16'b0010001011001111; 
assign lut_table[1596] = 16'b0010001011011101; 
assign lut_table[1597] = 16'b0010001011011110; 
assign lut_table[1598] = 16'b0010001011011111; 
assign lut_table[1599] = 16'b0010001011101110; 
assign lut_table[1600] = 16'b0010001011101111; 
assign lut_table[1601] = 16'b0010001011111111; 
assign lut_table[1602] = 16'b0010001100110011; 
assign lut_table[1603] = 16'b0010001100110100; 
assign lut_table[1604] = 16'b0010001100110101; 
assign lut_table[1605] = 16'b0010001100110110; 
assign lut_table[1606] = 16'b0010001100110111; 
assign lut_table[1607] = 16'b0010001100111000; 
assign lut_table[1608] = 16'b0010001100111001; 
assign lut_table[1609] = 16'b0010001100111010; 
assign lut_table[1610] = 16'b0010001100111011; 
assign lut_table[1611] = 16'b0010001100111100; 
assign lut_table[1612] = 16'b0010001100111101; 
assign lut_table[1613] = 16'b0010001100111110; 
assign lut_table[1614] = 16'b0010001100111111; 
assign lut_table[1615] = 16'b0010001101000100; 
assign lut_table[1616] = 16'b0010001101000101; 
assign lut_table[1617] = 16'b0010001101000110; 
assign lut_table[1618] = 16'b0010001101000111; 
assign lut_table[1619] = 16'b0010001101001000; 
assign lut_table[1620] = 16'b0010001101001001; 
assign lut_table[1621] = 16'b0010001101001010; 
assign lut_table[1622] = 16'b0010001101001011; 
assign lut_table[1623] = 16'b0010001101001100; 
assign lut_table[1624] = 16'b0010001101001101; 
assign lut_table[1625] = 16'b0010001101001110; 
assign lut_table[1626] = 16'b0010001101001111; 
assign lut_table[1627] = 16'b0010001101010101; 
assign lut_table[1628] = 16'b0010001101010110; 
assign lut_table[1629] = 16'b0010001101010111; 
assign lut_table[1630] = 16'b0010001101011000; 
assign lut_table[1631] = 16'b0010001101011001; 
assign lut_table[1632] = 16'b0010001101011010; 
assign lut_table[1633] = 16'b0010001101011011; 
assign lut_table[1634] = 16'b0010001101011100; 
assign lut_table[1635] = 16'b0010001101011101; 
assign lut_table[1636] = 16'b0010001101011110; 
assign lut_table[1637] = 16'b0010001101011111; 
assign lut_table[1638] = 16'b0010001101100110; 
assign lut_table[1639] = 16'b0010001101100111; 
assign lut_table[1640] = 16'b0010001101101000; 
assign lut_table[1641] = 16'b0010001101101001; 
assign lut_table[1642] = 16'b0010001101101010; 
assign lut_table[1643] = 16'b0010001101101011; 
assign lut_table[1644] = 16'b0010001101101100; 
assign lut_table[1645] = 16'b0010001101101101; 
assign lut_table[1646] = 16'b0010001101101110; 
assign lut_table[1647] = 16'b0010001101101111; 
assign lut_table[1648] = 16'b0010001101110111; 
assign lut_table[1649] = 16'b0010001101111000; 
assign lut_table[1650] = 16'b0010001101111001; 
assign lut_table[1651] = 16'b0010001101111010; 
assign lut_table[1652] = 16'b0010001101111011; 
assign lut_table[1653] = 16'b0010001101111100; 
assign lut_table[1654] = 16'b0010001101111101; 
assign lut_table[1655] = 16'b0010001101111110; 
assign lut_table[1656] = 16'b0010001101111111; 
assign lut_table[1657] = 16'b0010001110001000; 
assign lut_table[1658] = 16'b0010001110001001; 
assign lut_table[1659] = 16'b0010001110001010; 
assign lut_table[1660] = 16'b0010001110001011; 
assign lut_table[1661] = 16'b0010001110001100; 
assign lut_table[1662] = 16'b0010001110001101; 
assign lut_table[1663] = 16'b0010001110001110; 
assign lut_table[1664] = 16'b0010001110001111; 
assign lut_table[1665] = 16'b0010001110011001; 
assign lut_table[1666] = 16'b0010001110011010; 
assign lut_table[1667] = 16'b0010001110011011; 
assign lut_table[1668] = 16'b0010001110011100; 
assign lut_table[1669] = 16'b0010001110011101; 
assign lut_table[1670] = 16'b0010001110011110; 
assign lut_table[1671] = 16'b0010001110011111; 
assign lut_table[1672] = 16'b0010001110101010; 
assign lut_table[1673] = 16'b0010001110101011; 
assign lut_table[1674] = 16'b0010001110101100; 
assign lut_table[1675] = 16'b0010001110101101; 
assign lut_table[1676] = 16'b0010001110101110; 
assign lut_table[1677] = 16'b0010001110101111; 
assign lut_table[1678] = 16'b0010001110111011; 
assign lut_table[1679] = 16'b0010001110111100; 
assign lut_table[1680] = 16'b0010001110111101; 
assign lut_table[1681] = 16'b0010001110111110; 
assign lut_table[1682] = 16'b0010001110111111; 
assign lut_table[1683] = 16'b0010001111001100; 
assign lut_table[1684] = 16'b0010001111001101; 
assign lut_table[1685] = 16'b0010001111001110; 
assign lut_table[1686] = 16'b0010001111001111; 
assign lut_table[1687] = 16'b0010001111011101; 
assign lut_table[1688] = 16'b0010001111011110; 
assign lut_table[1689] = 16'b0010001111011111; 
assign lut_table[1690] = 16'b0010001111101110; 
assign lut_table[1691] = 16'b0010001111101111; 
assign lut_table[1692] = 16'b0010001111111111; 
assign lut_table[1693] = 16'b0010010001000100; 
assign lut_table[1694] = 16'b0010010001000101; 
assign lut_table[1695] = 16'b0010010001000110; 
assign lut_table[1696] = 16'b0010010001000111; 
assign lut_table[1697] = 16'b0010010001001000; 
assign lut_table[1698] = 16'b0010010001001001; 
assign lut_table[1699] = 16'b0010010001001010; 
assign lut_table[1700] = 16'b0010010001001011; 
assign lut_table[1701] = 16'b0010010001001100; 
assign lut_table[1702] = 16'b0010010001001101; 
assign lut_table[1703] = 16'b0010010001001110; 
assign lut_table[1704] = 16'b0010010001001111; 
assign lut_table[1705] = 16'b0010010001010101; 
assign lut_table[1706] = 16'b0010010001010110; 
assign lut_table[1707] = 16'b0010010001010111; 
assign lut_table[1708] = 16'b0010010001011000; 
assign lut_table[1709] = 16'b0010010001011001; 
assign lut_table[1710] = 16'b0010010001011010; 
assign lut_table[1711] = 16'b0010010001011011; 
assign lut_table[1712] = 16'b0010010001011100; 
assign lut_table[1713] = 16'b0010010001011101; 
assign lut_table[1714] = 16'b0010010001011110; 
assign lut_table[1715] = 16'b0010010001011111; 
assign lut_table[1716] = 16'b0010010001100110; 
assign lut_table[1717] = 16'b0010010001100111; 
assign lut_table[1718] = 16'b0010010001101000; 
assign lut_table[1719] = 16'b0010010001101001; 
assign lut_table[1720] = 16'b0010010001101010; 
assign lut_table[1721] = 16'b0010010001101011; 
assign lut_table[1722] = 16'b0010010001101100; 
assign lut_table[1723] = 16'b0010010001101101; 
assign lut_table[1724] = 16'b0010010001101110; 
assign lut_table[1725] = 16'b0010010001101111; 
assign lut_table[1726] = 16'b0010010001110111; 
assign lut_table[1727] = 16'b0010010001111000; 
assign lut_table[1728] = 16'b0010010001111001; 
assign lut_table[1729] = 16'b0010010001111010; 
assign lut_table[1730] = 16'b0010010001111011; 
assign lut_table[1731] = 16'b0010010001111100; 
assign lut_table[1732] = 16'b0010010001111101; 
assign lut_table[1733] = 16'b0010010001111110; 
assign lut_table[1734] = 16'b0010010001111111; 
assign lut_table[1735] = 16'b0010010010001000; 
assign lut_table[1736] = 16'b0010010010001001; 
assign lut_table[1737] = 16'b0010010010001010; 
assign lut_table[1738] = 16'b0010010010001011; 
assign lut_table[1739] = 16'b0010010010001100; 
assign lut_table[1740] = 16'b0010010010001101; 
assign lut_table[1741] = 16'b0010010010001110; 
assign lut_table[1742] = 16'b0010010010001111; 
assign lut_table[1743] = 16'b0010010010011001; 
assign lut_table[1744] = 16'b0010010010011010; 
assign lut_table[1745] = 16'b0010010010011011; 
assign lut_table[1746] = 16'b0010010010011100; 
assign lut_table[1747] = 16'b0010010010011101; 
assign lut_table[1748] = 16'b0010010010011110; 
assign lut_table[1749] = 16'b0010010010011111; 
assign lut_table[1750] = 16'b0010010010101010; 
assign lut_table[1751] = 16'b0010010010101011; 
assign lut_table[1752] = 16'b0010010010101100; 
assign lut_table[1753] = 16'b0010010010101101; 
assign lut_table[1754] = 16'b0010010010101110; 
assign lut_table[1755] = 16'b0010010010101111; 
assign lut_table[1756] = 16'b0010010010111011; 
assign lut_table[1757] = 16'b0010010010111100; 
assign lut_table[1758] = 16'b0010010010111101; 
assign lut_table[1759] = 16'b0010010010111110; 
assign lut_table[1760] = 16'b0010010010111111; 
assign lut_table[1761] = 16'b0010010011001100; 
assign lut_table[1762] = 16'b0010010011001101; 
assign lut_table[1763] = 16'b0010010011001110; 
assign lut_table[1764] = 16'b0010010011001111; 
assign lut_table[1765] = 16'b0010010011011101; 
assign lut_table[1766] = 16'b0010010011011110; 
assign lut_table[1767] = 16'b0010010011011111; 
assign lut_table[1768] = 16'b0010010011101110; 
assign lut_table[1769] = 16'b0010010011101111; 
assign lut_table[1770] = 16'b0010010011111111; 
assign lut_table[1771] = 16'b0010010101010101; 
assign lut_table[1772] = 16'b0010010101010110; 
assign lut_table[1773] = 16'b0010010101010111; 
assign lut_table[1774] = 16'b0010010101011000; 
assign lut_table[1775] = 16'b0010010101011001; 
assign lut_table[1776] = 16'b0010010101011010; 
assign lut_table[1777] = 16'b0010010101011011; 
assign lut_table[1778] = 16'b0010010101011100; 
assign lut_table[1779] = 16'b0010010101011101; 
assign lut_table[1780] = 16'b0010010101011110; 
assign lut_table[1781] = 16'b0010010101011111; 
assign lut_table[1782] = 16'b0010010101100110; 
assign lut_table[1783] = 16'b0010010101100111; 
assign lut_table[1784] = 16'b0010010101101000; 
assign lut_table[1785] = 16'b0010010101101001; 
assign lut_table[1786] = 16'b0010010101101010; 
assign lut_table[1787] = 16'b0010010101101011; 
assign lut_table[1788] = 16'b0010010101101100; 
assign lut_table[1789] = 16'b0010010101101101; 
assign lut_table[1790] = 16'b0010010101101110; 
assign lut_table[1791] = 16'b0010010101101111; 
assign lut_table[1792] = 16'b0010010101110111; 
assign lut_table[1793] = 16'b0010010101111000; 
assign lut_table[1794] = 16'b0010010101111001; 
assign lut_table[1795] = 16'b0010010101111010; 
assign lut_table[1796] = 16'b0010010101111011; 
assign lut_table[1797] = 16'b0010010101111100; 
assign lut_table[1798] = 16'b0010010101111101; 
assign lut_table[1799] = 16'b0010010101111110; 
assign lut_table[1800] = 16'b0010010101111111; 
assign lut_table[1801] = 16'b0010010110001000; 
assign lut_table[1802] = 16'b0010010110001001; 
assign lut_table[1803] = 16'b0010010110001010; 
assign lut_table[1804] = 16'b0010010110001011; 
assign lut_table[1805] = 16'b0010010110001100; 
assign lut_table[1806] = 16'b0010010110001101; 
assign lut_table[1807] = 16'b0010010110001110; 
assign lut_table[1808] = 16'b0010010110001111; 
assign lut_table[1809] = 16'b0010010110011001; 
assign lut_table[1810] = 16'b0010010110011010; 
assign lut_table[1811] = 16'b0010010110011011; 
assign lut_table[1812] = 16'b0010010110011100; 
assign lut_table[1813] = 16'b0010010110011101; 
assign lut_table[1814] = 16'b0010010110011110; 
assign lut_table[1815] = 16'b0010010110011111; 
assign lut_table[1816] = 16'b0010010110101010; 
assign lut_table[1817] = 16'b0010010110101011; 
assign lut_table[1818] = 16'b0010010110101100; 
assign lut_table[1819] = 16'b0010010110101101; 
assign lut_table[1820] = 16'b0010010110101110; 
assign lut_table[1821] = 16'b0010010110101111; 
assign lut_table[1822] = 16'b0010010110111011; 
assign lut_table[1823] = 16'b0010010110111100; 
assign lut_table[1824] = 16'b0010010110111101; 
assign lut_table[1825] = 16'b0010010110111110; 
assign lut_table[1826] = 16'b0010010110111111; 
assign lut_table[1827] = 16'b0010010111001100; 
assign lut_table[1828] = 16'b0010010111001101; 
assign lut_table[1829] = 16'b0010010111001110; 
assign lut_table[1830] = 16'b0010010111001111; 
assign lut_table[1831] = 16'b0010010111011101; 
assign lut_table[1832] = 16'b0010010111011110; 
assign lut_table[1833] = 16'b0010010111011111; 
assign lut_table[1834] = 16'b0010010111101110; 
assign lut_table[1835] = 16'b0010010111101111; 
assign lut_table[1836] = 16'b0010010111111111; 
assign lut_table[1837] = 16'b0010011001100110; 
assign lut_table[1838] = 16'b0010011001100111; 
assign lut_table[1839] = 16'b0010011001101000; 
assign lut_table[1840] = 16'b0010011001101001; 
assign lut_table[1841] = 16'b0010011001101010; 
assign lut_table[1842] = 16'b0010011001101011; 
assign lut_table[1843] = 16'b0010011001101100; 
assign lut_table[1844] = 16'b0010011001101101; 
assign lut_table[1845] = 16'b0010011001101110; 
assign lut_table[1846] = 16'b0010011001101111; 
assign lut_table[1847] = 16'b0010011001110111; 
assign lut_table[1848] = 16'b0010011001111000; 
assign lut_table[1849] = 16'b0010011001111001; 
assign lut_table[1850] = 16'b0010011001111010; 
assign lut_table[1851] = 16'b0010011001111011; 
assign lut_table[1852] = 16'b0010011001111100; 
assign lut_table[1853] = 16'b0010011001111101; 
assign lut_table[1854] = 16'b0010011001111110; 
assign lut_table[1855] = 16'b0010011001111111; 
assign lut_table[1856] = 16'b0010011010001000; 
assign lut_table[1857] = 16'b0010011010001001; 
assign lut_table[1858] = 16'b0010011010001010; 
assign lut_table[1859] = 16'b0010011010001011; 
assign lut_table[1860] = 16'b0010011010001100; 
assign lut_table[1861] = 16'b0010011010001101; 
assign lut_table[1862] = 16'b0010011010001110; 
assign lut_table[1863] = 16'b0010011010001111; 
assign lut_table[1864] = 16'b0010011010011001; 
assign lut_table[1865] = 16'b0010011010011010; 
assign lut_table[1866] = 16'b0010011010011011; 
assign lut_table[1867] = 16'b0010011010011100; 
assign lut_table[1868] = 16'b0010011010011101; 
assign lut_table[1869] = 16'b0010011010011110; 
assign lut_table[1870] = 16'b0010011010011111; 
assign lut_table[1871] = 16'b0010011010101010; 
assign lut_table[1872] = 16'b0010011010101011; 
assign lut_table[1873] = 16'b0010011010101100; 
assign lut_table[1874] = 16'b0010011010101101; 
assign lut_table[1875] = 16'b0010011010101110; 
assign lut_table[1876] = 16'b0010011010101111; 
assign lut_table[1877] = 16'b0010011010111011; 
assign lut_table[1878] = 16'b0010011010111100; 
assign lut_table[1879] = 16'b0010011010111101; 
assign lut_table[1880] = 16'b0010011010111110; 
assign lut_table[1881] = 16'b0010011010111111; 
assign lut_table[1882] = 16'b0010011011001100; 
assign lut_table[1883] = 16'b0010011011001101; 
assign lut_table[1884] = 16'b0010011011001110; 
assign lut_table[1885] = 16'b0010011011001111; 
assign lut_table[1886] = 16'b0010011011011101; 
assign lut_table[1887] = 16'b0010011011011110; 
assign lut_table[1888] = 16'b0010011011011111; 
assign lut_table[1889] = 16'b0010011011101110; 
assign lut_table[1890] = 16'b0010011011101111; 
assign lut_table[1891] = 16'b0010011011111111; 
assign lut_table[1892] = 16'b0010011101110111; 
assign lut_table[1893] = 16'b0010011101111000; 
assign lut_table[1894] = 16'b0010011101111001; 
assign lut_table[1895] = 16'b0010011101111010; 
assign lut_table[1896] = 16'b0010011101111011; 
assign lut_table[1897] = 16'b0010011101111100; 
assign lut_table[1898] = 16'b0010011101111101; 
assign lut_table[1899] = 16'b0010011101111110; 
assign lut_table[1900] = 16'b0010011101111111; 
assign lut_table[1901] = 16'b0010011110001000; 
assign lut_table[1902] = 16'b0010011110001001; 
assign lut_table[1903] = 16'b0010011110001010; 
assign lut_table[1904] = 16'b0010011110001011; 
assign lut_table[1905] = 16'b0010011110001100; 
assign lut_table[1906] = 16'b0010011110001101; 
assign lut_table[1907] = 16'b0010011110001110; 
assign lut_table[1908] = 16'b0010011110001111; 
assign lut_table[1909] = 16'b0010011110011001; 
assign lut_table[1910] = 16'b0010011110011010; 
assign lut_table[1911] = 16'b0010011110011011; 
assign lut_table[1912] = 16'b0010011110011100; 
assign lut_table[1913] = 16'b0010011110011101; 
assign lut_table[1914] = 16'b0010011110011110; 
assign lut_table[1915] = 16'b0010011110011111; 
assign lut_table[1916] = 16'b0010011110101010; 
assign lut_table[1917] = 16'b0010011110101011; 
assign lut_table[1918] = 16'b0010011110101100; 
assign lut_table[1919] = 16'b0010011110101101; 
assign lut_table[1920] = 16'b0010011110101110; 
assign lut_table[1921] = 16'b0010011110101111; 
assign lut_table[1922] = 16'b0010011110111011; 
assign lut_table[1923] = 16'b0010011110111100; 
assign lut_table[1924] = 16'b0010011110111101; 
assign lut_table[1925] = 16'b0010011110111110; 
assign lut_table[1926] = 16'b0010011110111111; 
assign lut_table[1927] = 16'b0010011111001100; 
assign lut_table[1928] = 16'b0010011111001101; 
assign lut_table[1929] = 16'b0010011111001110; 
assign lut_table[1930] = 16'b0010011111001111; 
assign lut_table[1931] = 16'b0010011111011101; 
assign lut_table[1932] = 16'b0010011111011110; 
assign lut_table[1933] = 16'b0010011111011111; 
assign lut_table[1934] = 16'b0010011111101110; 
assign lut_table[1935] = 16'b0010011111101111; 
assign lut_table[1936] = 16'b0010011111111111; 
assign lut_table[1937] = 16'b0010100010001000; 
assign lut_table[1938] = 16'b0010100010001001; 
assign lut_table[1939] = 16'b0010100010001010; 
assign lut_table[1940] = 16'b0010100010001011; 
assign lut_table[1941] = 16'b0010100010001100; 
assign lut_table[1942] = 16'b0010100010001101; 
assign lut_table[1943] = 16'b0010100010001110; 
assign lut_table[1944] = 16'b0010100010001111; 
assign lut_table[1945] = 16'b0010100010011001; 
assign lut_table[1946] = 16'b0010100010011010; 
assign lut_table[1947] = 16'b0010100010011011; 
assign lut_table[1948] = 16'b0010100010011100; 
assign lut_table[1949] = 16'b0010100010011101; 
assign lut_table[1950] = 16'b0010100010011110; 
assign lut_table[1951] = 16'b0010100010011111; 
assign lut_table[1952] = 16'b0010100010101010; 
assign lut_table[1953] = 16'b0010100010101011; 
assign lut_table[1954] = 16'b0010100010101100; 
assign lut_table[1955] = 16'b0010100010101101; 
assign lut_table[1956] = 16'b0010100010101110; 
assign lut_table[1957] = 16'b0010100010101111; 
assign lut_table[1958] = 16'b0010100010111011; 
assign lut_table[1959] = 16'b0010100010111100; 
assign lut_table[1960] = 16'b0010100010111101; 
assign lut_table[1961] = 16'b0010100010111110; 
assign lut_table[1962] = 16'b0010100010111111; 
assign lut_table[1963] = 16'b0010100011001100; 
assign lut_table[1964] = 16'b0010100011001101; 
assign lut_table[1965] = 16'b0010100011001110; 
assign lut_table[1966] = 16'b0010100011001111; 
assign lut_table[1967] = 16'b0010100011011101; 
assign lut_table[1968] = 16'b0010100011011110; 
assign lut_table[1969] = 16'b0010100011011111; 
assign lut_table[1970] = 16'b0010100011101110; 
assign lut_table[1971] = 16'b0010100011101111; 
assign lut_table[1972] = 16'b0010100011111111; 
assign lut_table[1973] = 16'b0010100110011001; 
assign lut_table[1974] = 16'b0010100110011010; 
assign lut_table[1975] = 16'b0010100110011011; 
assign lut_table[1976] = 16'b0010100110011100; 
assign lut_table[1977] = 16'b0010100110011101; 
assign lut_table[1978] = 16'b0010100110011110; 
assign lut_table[1979] = 16'b0010100110011111; 
assign lut_table[1980] = 16'b0010100110101010; 
assign lut_table[1981] = 16'b0010100110101011; 
assign lut_table[1982] = 16'b0010100110101100; 
assign lut_table[1983] = 16'b0010100110101101; 
assign lut_table[1984] = 16'b0010100110101110; 
assign lut_table[1985] = 16'b0010100110101111; 
assign lut_table[1986] = 16'b0010100110111011; 
assign lut_table[1987] = 16'b0010100110111100; 
assign lut_table[1988] = 16'b0010100110111101; 
assign lut_table[1989] = 16'b0010100110111110; 
assign lut_table[1990] = 16'b0010100110111111; 
assign lut_table[1991] = 16'b0010100111001100; 
assign lut_table[1992] = 16'b0010100111001101; 
assign lut_table[1993] = 16'b0010100111001110; 
assign lut_table[1994] = 16'b0010100111001111; 
assign lut_table[1995] = 16'b0010100111011101; 
assign lut_table[1996] = 16'b0010100111011110; 
assign lut_table[1997] = 16'b0010100111011111; 
assign lut_table[1998] = 16'b0010100111101110; 
assign lut_table[1999] = 16'b0010100111101111; 
assign lut_table[2000] = 16'b0010100111111111; 
assign lut_table[2001] = 16'b0010101010101010; 
assign lut_table[2002] = 16'b0010101010101011; 
assign lut_table[2003] = 16'b0010101010101100; 
assign lut_table[2004] = 16'b0010101010101101; 
assign lut_table[2005] = 16'b0010101010101110; 
assign lut_table[2006] = 16'b0010101010101111; 
assign lut_table[2007] = 16'b0010101010111011; 
assign lut_table[2008] = 16'b0010101010111100; 
assign lut_table[2009] = 16'b0010101010111101; 
assign lut_table[2010] = 16'b0010101010111110; 
assign lut_table[2011] = 16'b0010101010111111; 
assign lut_table[2012] = 16'b0010101011001100; 
assign lut_table[2013] = 16'b0010101011001101; 
assign lut_table[2014] = 16'b0010101011001110; 
assign lut_table[2015] = 16'b0010101011001111; 
assign lut_table[2016] = 16'b0010101011011101; 
assign lut_table[2017] = 16'b0010101011011110; 
assign lut_table[2018] = 16'b0010101011011111; 
assign lut_table[2019] = 16'b0010101011101110; 
assign lut_table[2020] = 16'b0010101011101111; 
assign lut_table[2021] = 16'b0010101011111111; 
assign lut_table[2022] = 16'b0010101110111011; 
assign lut_table[2023] = 16'b0010101110111100; 
assign lut_table[2024] = 16'b0010101110111101; 
assign lut_table[2025] = 16'b0010101110111110; 
assign lut_table[2026] = 16'b0010101110111111; 
assign lut_table[2027] = 16'b0010101111001100; 
assign lut_table[2028] = 16'b0010101111001101; 
assign lut_table[2029] = 16'b0010101111001110; 
assign lut_table[2030] = 16'b0010101111001111; 
assign lut_table[2031] = 16'b0010101111011101; 
assign lut_table[2032] = 16'b0010101111011110; 
assign lut_table[2033] = 16'b0010101111011111; 
assign lut_table[2034] = 16'b0010101111101110; 
assign lut_table[2035] = 16'b0010101111101111; 
assign lut_table[2036] = 16'b0010101111111111; 
assign lut_table[2037] = 16'b0010110011001100; 
assign lut_table[2038] = 16'b0010110011001101; 
assign lut_table[2039] = 16'b0010110011001110; 
assign lut_table[2040] = 16'b0010110011001111; 
assign lut_table[2041] = 16'b0010110011011101; 
assign lut_table[2042] = 16'b0010110011011110; 
assign lut_table[2043] = 16'b0010110011011111; 
assign lut_table[2044] = 16'b0010110011101110; 
assign lut_table[2045] = 16'b0010110011101111; 
assign lut_table[2046] = 16'b0010110011111111; 
assign lut_table[2047] = 16'b0010110111011101; 
assign lut_table[2048] = 16'b0010110111011110; 
assign lut_table[2049] = 16'b0010110111011111; 
assign lut_table[2050] = 16'b0010110111101110; 
assign lut_table[2051] = 16'b0010110111101111; 
assign lut_table[2052] = 16'b0010110111111111; 
assign lut_table[2053] = 16'b0010111011101110; 
assign lut_table[2054] = 16'b0010111011101111; 
assign lut_table[2055] = 16'b0010111011111111; 
assign lut_table[2056] = 16'b0010111111111111; 
assign lut_table[2057] = 16'b0011001100110011; 
assign lut_table[2058] = 16'b0011001100110100; 
assign lut_table[2059] = 16'b0011001100110101; 
assign lut_table[2060] = 16'b0011001100110110; 
assign lut_table[2061] = 16'b0011001100110111; 
assign lut_table[2062] = 16'b0011001100111000; 
assign lut_table[2063] = 16'b0011001100111001; 
assign lut_table[2064] = 16'b0011001100111010; 
assign lut_table[2065] = 16'b0011001100111011; 
assign lut_table[2066] = 16'b0011001100111100; 
assign lut_table[2067] = 16'b0011001100111101; 
assign lut_table[2068] = 16'b0011001100111110; 
assign lut_table[2069] = 16'b0011001100111111; 
assign lut_table[2070] = 16'b0011001101000100; 
assign lut_table[2071] = 16'b0011001101000101; 
assign lut_table[2072] = 16'b0011001101000110; 
assign lut_table[2073] = 16'b0011001101000111; 
assign lut_table[2074] = 16'b0011001101001000; 
assign lut_table[2075] = 16'b0011001101001001; 
assign lut_table[2076] = 16'b0011001101001010; 
assign lut_table[2077] = 16'b0011001101001011; 
assign lut_table[2078] = 16'b0011001101001100; 
assign lut_table[2079] = 16'b0011001101001101; 
assign lut_table[2080] = 16'b0011001101001110; 
assign lut_table[2081] = 16'b0011001101001111; 
assign lut_table[2082] = 16'b0011001101010101; 
assign lut_table[2083] = 16'b0011001101010110; 
assign lut_table[2084] = 16'b0011001101010111; 
assign lut_table[2085] = 16'b0011001101011000; 
assign lut_table[2086] = 16'b0011001101011001; 
assign lut_table[2087] = 16'b0011001101011010; 
assign lut_table[2088] = 16'b0011001101011011; 
assign lut_table[2089] = 16'b0011001101011100; 
assign lut_table[2090] = 16'b0011001101011101; 
assign lut_table[2091] = 16'b0011001101011110; 
assign lut_table[2092] = 16'b0011001101011111; 
assign lut_table[2093] = 16'b0011001101100110; 
assign lut_table[2094] = 16'b0011001101100111; 
assign lut_table[2095] = 16'b0011001101101000; 
assign lut_table[2096] = 16'b0011001101101001; 
assign lut_table[2097] = 16'b0011001101101010; 
assign lut_table[2098] = 16'b0011001101101011; 
assign lut_table[2099] = 16'b0011001101101100; 
assign lut_table[2100] = 16'b0011001101101101; 
assign lut_table[2101] = 16'b0011001101101110; 
assign lut_table[2102] = 16'b0011001101101111; 
assign lut_table[2103] = 16'b0011001101110111; 
assign lut_table[2104] = 16'b0011001101111000; 
assign lut_table[2105] = 16'b0011001101111001; 
assign lut_table[2106] = 16'b0011001101111010; 
assign lut_table[2107] = 16'b0011001101111011; 
assign lut_table[2108] = 16'b0011001101111100; 
assign lut_table[2109] = 16'b0011001101111101; 
assign lut_table[2110] = 16'b0011001101111110; 
assign lut_table[2111] = 16'b0011001101111111; 
assign lut_table[2112] = 16'b0011001110001000; 
assign lut_table[2113] = 16'b0011001110001001; 
assign lut_table[2114] = 16'b0011001110001010; 
assign lut_table[2115] = 16'b0011001110001011; 
assign lut_table[2116] = 16'b0011001110001100; 
assign lut_table[2117] = 16'b0011001110001101; 
assign lut_table[2118] = 16'b0011001110001110; 
assign lut_table[2119] = 16'b0011001110001111; 
assign lut_table[2120] = 16'b0011001110011001; 
assign lut_table[2121] = 16'b0011001110011010; 
assign lut_table[2122] = 16'b0011001110011011; 
assign lut_table[2123] = 16'b0011001110011100; 
assign lut_table[2124] = 16'b0011001110011101; 
assign lut_table[2125] = 16'b0011001110011110; 
assign lut_table[2126] = 16'b0011001110011111; 
assign lut_table[2127] = 16'b0011001110101010; 
assign lut_table[2128] = 16'b0011001110101011; 
assign lut_table[2129] = 16'b0011001110101100; 
assign lut_table[2130] = 16'b0011001110101101; 
assign lut_table[2131] = 16'b0011001110101110; 
assign lut_table[2132] = 16'b0011001110101111; 
assign lut_table[2133] = 16'b0011001110111011; 
assign lut_table[2134] = 16'b0011001110111100; 
assign lut_table[2135] = 16'b0011001110111101; 
assign lut_table[2136] = 16'b0011001110111110; 
assign lut_table[2137] = 16'b0011001110111111; 
assign lut_table[2138] = 16'b0011001111001100; 
assign lut_table[2139] = 16'b0011001111001101; 
assign lut_table[2140] = 16'b0011001111001110; 
assign lut_table[2141] = 16'b0011001111001111; 
assign lut_table[2142] = 16'b0011001111011101; 
assign lut_table[2143] = 16'b0011001111011110; 
assign lut_table[2144] = 16'b0011001111011111; 
assign lut_table[2145] = 16'b0011001111101110; 
assign lut_table[2146] = 16'b0011001111101111; 
assign lut_table[2147] = 16'b0011001111111111; 
assign lut_table[2148] = 16'b0011010001000100; 
assign lut_table[2149] = 16'b0011010001000101; 
assign lut_table[2150] = 16'b0011010001000110; 
assign lut_table[2151] = 16'b0011010001000111; 
assign lut_table[2152] = 16'b0011010001001000; 
assign lut_table[2153] = 16'b0011010001001001; 
assign lut_table[2154] = 16'b0011010001001010; 
assign lut_table[2155] = 16'b0011010001001011; 
assign lut_table[2156] = 16'b0011010001001100; 
assign lut_table[2157] = 16'b0011010001001101; 
assign lut_table[2158] = 16'b0011010001001110; 
assign lut_table[2159] = 16'b0011010001001111; 
assign lut_table[2160] = 16'b0011010001010101; 
assign lut_table[2161] = 16'b0011010001010110; 
assign lut_table[2162] = 16'b0011010001010111; 
assign lut_table[2163] = 16'b0011010001011000; 
assign lut_table[2164] = 16'b0011010001011001; 
assign lut_table[2165] = 16'b0011010001011010; 
assign lut_table[2166] = 16'b0011010001011011; 
assign lut_table[2167] = 16'b0011010001011100; 
assign lut_table[2168] = 16'b0011010001011101; 
assign lut_table[2169] = 16'b0011010001011110; 
assign lut_table[2170] = 16'b0011010001011111; 
assign lut_table[2171] = 16'b0011010001100110; 
assign lut_table[2172] = 16'b0011010001100111; 
assign lut_table[2173] = 16'b0011010001101000; 
assign lut_table[2174] = 16'b0011010001101001; 
assign lut_table[2175] = 16'b0011010001101010; 
assign lut_table[2176] = 16'b0011010001101011; 
assign lut_table[2177] = 16'b0011010001101100; 
assign lut_table[2178] = 16'b0011010001101101; 
assign lut_table[2179] = 16'b0011010001101110; 
assign lut_table[2180] = 16'b0011010001101111; 
assign lut_table[2181] = 16'b0011010001110111; 
assign lut_table[2182] = 16'b0011010001111000; 
assign lut_table[2183] = 16'b0011010001111001; 
assign lut_table[2184] = 16'b0011010001111010; 
assign lut_table[2185] = 16'b0011010001111011; 
assign lut_table[2186] = 16'b0011010001111100; 
assign lut_table[2187] = 16'b0011010001111101; 
assign lut_table[2188] = 16'b0011010001111110; 
assign lut_table[2189] = 16'b0011010001111111; 
assign lut_table[2190] = 16'b0011010010001000; 
assign lut_table[2191] = 16'b0011010010001001; 
assign lut_table[2192] = 16'b0011010010001010; 
assign lut_table[2193] = 16'b0011010010001011; 
assign lut_table[2194] = 16'b0011010010001100; 
assign lut_table[2195] = 16'b0011010010001101; 
assign lut_table[2196] = 16'b0011010010001110; 
assign lut_table[2197] = 16'b0011010010001111; 
assign lut_table[2198] = 16'b0011010010011001; 
assign lut_table[2199] = 16'b0011010010011010; 
assign lut_table[2200] = 16'b0011010010011011; 
assign lut_table[2201] = 16'b0011010010011100; 
assign lut_table[2202] = 16'b0011010010011101; 
assign lut_table[2203] = 16'b0011010010011110; 
assign lut_table[2204] = 16'b0011010010011111; 
assign lut_table[2205] = 16'b0011010010101010; 
assign lut_table[2206] = 16'b0011010010101011; 
assign lut_table[2207] = 16'b0011010010101100; 
assign lut_table[2208] = 16'b0011010010101101; 
assign lut_table[2209] = 16'b0011010010101110; 
assign lut_table[2210] = 16'b0011010010101111; 
assign lut_table[2211] = 16'b0011010010111011; 
assign lut_table[2212] = 16'b0011010010111100; 
assign lut_table[2213] = 16'b0011010010111101; 
assign lut_table[2214] = 16'b0011010010111110; 
assign lut_table[2215] = 16'b0011010010111111; 
assign lut_table[2216] = 16'b0011010011001100; 
assign lut_table[2217] = 16'b0011010011001101; 
assign lut_table[2218] = 16'b0011010011001110; 
assign lut_table[2219] = 16'b0011010011001111; 
assign lut_table[2220] = 16'b0011010011011101; 
assign lut_table[2221] = 16'b0011010011011110; 
assign lut_table[2222] = 16'b0011010011011111; 
assign lut_table[2223] = 16'b0011010011101110; 
assign lut_table[2224] = 16'b0011010011101111; 
assign lut_table[2225] = 16'b0011010011111111; 
assign lut_table[2226] = 16'b0011010101010101; 
assign lut_table[2227] = 16'b0011010101010110; 
assign lut_table[2228] = 16'b0011010101010111; 
assign lut_table[2229] = 16'b0011010101011000; 
assign lut_table[2230] = 16'b0011010101011001; 
assign lut_table[2231] = 16'b0011010101011010; 
assign lut_table[2232] = 16'b0011010101011011; 
assign lut_table[2233] = 16'b0011010101011100; 
assign lut_table[2234] = 16'b0011010101011101; 
assign lut_table[2235] = 16'b0011010101011110; 
assign lut_table[2236] = 16'b0011010101011111; 
assign lut_table[2237] = 16'b0011010101100110; 
assign lut_table[2238] = 16'b0011010101100111; 
assign lut_table[2239] = 16'b0011010101101000; 
assign lut_table[2240] = 16'b0011010101101001; 
assign lut_table[2241] = 16'b0011010101101010; 
assign lut_table[2242] = 16'b0011010101101011; 
assign lut_table[2243] = 16'b0011010101101100; 
assign lut_table[2244] = 16'b0011010101101101; 
assign lut_table[2245] = 16'b0011010101101110; 
assign lut_table[2246] = 16'b0011010101101111; 
assign lut_table[2247] = 16'b0011010101110111; 
assign lut_table[2248] = 16'b0011010101111000; 
assign lut_table[2249] = 16'b0011010101111001; 
assign lut_table[2250] = 16'b0011010101111010; 
assign lut_table[2251] = 16'b0011010101111011; 
assign lut_table[2252] = 16'b0011010101111100; 
assign lut_table[2253] = 16'b0011010101111101; 
assign lut_table[2254] = 16'b0011010101111110; 
assign lut_table[2255] = 16'b0011010101111111; 
assign lut_table[2256] = 16'b0011010110001000; 
assign lut_table[2257] = 16'b0011010110001001; 
assign lut_table[2258] = 16'b0011010110001010; 
assign lut_table[2259] = 16'b0011010110001011; 
assign lut_table[2260] = 16'b0011010110001100; 
assign lut_table[2261] = 16'b0011010110001101; 
assign lut_table[2262] = 16'b0011010110001110; 
assign lut_table[2263] = 16'b0011010110001111; 
assign lut_table[2264] = 16'b0011010110011001; 
assign lut_table[2265] = 16'b0011010110011010; 
assign lut_table[2266] = 16'b0011010110011011; 
assign lut_table[2267] = 16'b0011010110011100; 
assign lut_table[2268] = 16'b0011010110011101; 
assign lut_table[2269] = 16'b0011010110011110; 
assign lut_table[2270] = 16'b0011010110011111; 
assign lut_table[2271] = 16'b0011010110101010; 
assign lut_table[2272] = 16'b0011010110101011; 
assign lut_table[2273] = 16'b0011010110101100; 
assign lut_table[2274] = 16'b0011010110101101; 
assign lut_table[2275] = 16'b0011010110101110; 
assign lut_table[2276] = 16'b0011010110101111; 
assign lut_table[2277] = 16'b0011010110111011; 
assign lut_table[2278] = 16'b0011010110111100; 
assign lut_table[2279] = 16'b0011010110111101; 
assign lut_table[2280] = 16'b0011010110111110; 
assign lut_table[2281] = 16'b0011010110111111; 
assign lut_table[2282] = 16'b0011010111001100; 
assign lut_table[2283] = 16'b0011010111001101; 
assign lut_table[2284] = 16'b0011010111001110; 
assign lut_table[2285] = 16'b0011010111001111; 
assign lut_table[2286] = 16'b0011010111011101; 
assign lut_table[2287] = 16'b0011010111011110; 
assign lut_table[2288] = 16'b0011010111011111; 
assign lut_table[2289] = 16'b0011010111101110; 
assign lut_table[2290] = 16'b0011010111101111; 
assign lut_table[2291] = 16'b0011010111111111; 
assign lut_table[2292] = 16'b0011011001100110; 
assign lut_table[2293] = 16'b0011011001100111; 
assign lut_table[2294] = 16'b0011011001101000; 
assign lut_table[2295] = 16'b0011011001101001; 
assign lut_table[2296] = 16'b0011011001101010; 
assign lut_table[2297] = 16'b0011011001101011; 
assign lut_table[2298] = 16'b0011011001101100; 
assign lut_table[2299] = 16'b0011011001101101; 
assign lut_table[2300] = 16'b0011011001101110; 
assign lut_table[2301] = 16'b0011011001101111; 
assign lut_table[2302] = 16'b0011011001110111; 
assign lut_table[2303] = 16'b0011011001111000; 
assign lut_table[2304] = 16'b0011011001111001; 
assign lut_table[2305] = 16'b0011011001111010; 
assign lut_table[2306] = 16'b0011011001111011; 
assign lut_table[2307] = 16'b0011011001111100; 
assign lut_table[2308] = 16'b0011011001111101; 
assign lut_table[2309] = 16'b0011011001111110; 
assign lut_table[2310] = 16'b0011011001111111; 
assign lut_table[2311] = 16'b0011011010001000; 
assign lut_table[2312] = 16'b0011011010001001; 
assign lut_table[2313] = 16'b0011011010001010; 
assign lut_table[2314] = 16'b0011011010001011; 
assign lut_table[2315] = 16'b0011011010001100; 
assign lut_table[2316] = 16'b0011011010001101; 
assign lut_table[2317] = 16'b0011011010001110; 
assign lut_table[2318] = 16'b0011011010001111; 
assign lut_table[2319] = 16'b0011011010011001; 
assign lut_table[2320] = 16'b0011011010011010; 
assign lut_table[2321] = 16'b0011011010011011; 
assign lut_table[2322] = 16'b0011011010011100; 
assign lut_table[2323] = 16'b0011011010011101; 
assign lut_table[2324] = 16'b0011011010011110; 
assign lut_table[2325] = 16'b0011011010011111; 
assign lut_table[2326] = 16'b0011011010101010; 
assign lut_table[2327] = 16'b0011011010101011; 
assign lut_table[2328] = 16'b0011011010101100; 
assign lut_table[2329] = 16'b0011011010101101; 
assign lut_table[2330] = 16'b0011011010101110; 
assign lut_table[2331] = 16'b0011011010101111; 
assign lut_table[2332] = 16'b0011011010111011; 
assign lut_table[2333] = 16'b0011011010111100; 
assign lut_table[2334] = 16'b0011011010111101; 
assign lut_table[2335] = 16'b0011011010111110; 
assign lut_table[2336] = 16'b0011011010111111; 
assign lut_table[2337] = 16'b0011011011001100; 
assign lut_table[2338] = 16'b0011011011001101; 
assign lut_table[2339] = 16'b0011011011001110; 
assign lut_table[2340] = 16'b0011011011001111; 
assign lut_table[2341] = 16'b0011011011011101; 
assign lut_table[2342] = 16'b0011011011011110; 
assign lut_table[2343] = 16'b0011011011011111; 
assign lut_table[2344] = 16'b0011011011101110; 
assign lut_table[2345] = 16'b0011011011101111; 
assign lut_table[2346] = 16'b0011011011111111; 
assign lut_table[2347] = 16'b0011011101110111; 
assign lut_table[2348] = 16'b0011011101111000; 
assign lut_table[2349] = 16'b0011011101111001; 
assign lut_table[2350] = 16'b0011011101111010; 
assign lut_table[2351] = 16'b0011011101111011; 
assign lut_table[2352] = 16'b0011011101111100; 
assign lut_table[2353] = 16'b0011011101111101; 
assign lut_table[2354] = 16'b0011011101111110; 
assign lut_table[2355] = 16'b0011011101111111; 
assign lut_table[2356] = 16'b0011011110001000; 
assign lut_table[2357] = 16'b0011011110001001; 
assign lut_table[2358] = 16'b0011011110001010; 
assign lut_table[2359] = 16'b0011011110001011; 
assign lut_table[2360] = 16'b0011011110001100; 
assign lut_table[2361] = 16'b0011011110001101; 
assign lut_table[2362] = 16'b0011011110001110; 
assign lut_table[2363] = 16'b0011011110001111; 
assign lut_table[2364] = 16'b0011011110011001; 
assign lut_table[2365] = 16'b0011011110011010; 
assign lut_table[2366] = 16'b0011011110011011; 
assign lut_table[2367] = 16'b0011011110011100; 
assign lut_table[2368] = 16'b0011011110011101; 
assign lut_table[2369] = 16'b0011011110011110; 
assign lut_table[2370] = 16'b0011011110011111; 
assign lut_table[2371] = 16'b0011011110101010; 
assign lut_table[2372] = 16'b0011011110101011; 
assign lut_table[2373] = 16'b0011011110101100; 
assign lut_table[2374] = 16'b0011011110101101; 
assign lut_table[2375] = 16'b0011011110101110; 
assign lut_table[2376] = 16'b0011011110101111; 
assign lut_table[2377] = 16'b0011011110111011; 
assign lut_table[2378] = 16'b0011011110111100; 
assign lut_table[2379] = 16'b0011011110111101; 
assign lut_table[2380] = 16'b0011011110111110; 
assign lut_table[2381] = 16'b0011011110111111; 
assign lut_table[2382] = 16'b0011011111001100; 
assign lut_table[2383] = 16'b0011011111001101; 
assign lut_table[2384] = 16'b0011011111001110; 
assign lut_table[2385] = 16'b0011011111001111; 
assign lut_table[2386] = 16'b0011011111011101; 
assign lut_table[2387] = 16'b0011011111011110; 
assign lut_table[2388] = 16'b0011011111011111; 
assign lut_table[2389] = 16'b0011011111101110; 
assign lut_table[2390] = 16'b0011011111101111; 
assign lut_table[2391] = 16'b0011011111111111; 
assign lut_table[2392] = 16'b0011100010001000; 
assign lut_table[2393] = 16'b0011100010001001; 
assign lut_table[2394] = 16'b0011100010001010; 
assign lut_table[2395] = 16'b0011100010001011; 
assign lut_table[2396] = 16'b0011100010001100; 
assign lut_table[2397] = 16'b0011100010001101; 
assign lut_table[2398] = 16'b0011100010001110; 
assign lut_table[2399] = 16'b0011100010001111; 
assign lut_table[2400] = 16'b0011100010011001; 
assign lut_table[2401] = 16'b0011100010011010; 
assign lut_table[2402] = 16'b0011100010011011; 
assign lut_table[2403] = 16'b0011100010011100; 
assign lut_table[2404] = 16'b0011100010011101; 
assign lut_table[2405] = 16'b0011100010011110; 
assign lut_table[2406] = 16'b0011100010011111; 
assign lut_table[2407] = 16'b0011100010101010; 
assign lut_table[2408] = 16'b0011100010101011; 
assign lut_table[2409] = 16'b0011100010101100; 
assign lut_table[2410] = 16'b0011100010101101; 
assign lut_table[2411] = 16'b0011100010101110; 
assign lut_table[2412] = 16'b0011100010101111; 
assign lut_table[2413] = 16'b0011100010111011; 
assign lut_table[2414] = 16'b0011100010111100; 
assign lut_table[2415] = 16'b0011100010111101; 
assign lut_table[2416] = 16'b0011100010111110; 
assign lut_table[2417] = 16'b0011100010111111; 
assign lut_table[2418] = 16'b0011100011001100; 
assign lut_table[2419] = 16'b0011100011001101; 
assign lut_table[2420] = 16'b0011100011001110; 
assign lut_table[2421] = 16'b0011100011001111; 
assign lut_table[2422] = 16'b0011100011011101; 
assign lut_table[2423] = 16'b0011100011011110; 
assign lut_table[2424] = 16'b0011100011011111; 
assign lut_table[2425] = 16'b0011100011101110; 
assign lut_table[2426] = 16'b0011100011101111; 
assign lut_table[2427] = 16'b0011100011111111; 
assign lut_table[2428] = 16'b0011100110011001; 
assign lut_table[2429] = 16'b0011100110011010; 
assign lut_table[2430] = 16'b0011100110011011; 
assign lut_table[2431] = 16'b0011100110011100; 
assign lut_table[2432] = 16'b0011100110011101; 
assign lut_table[2433] = 16'b0011100110011110; 
assign lut_table[2434] = 16'b0011100110011111; 
assign lut_table[2435] = 16'b0011100110101010; 
assign lut_table[2436] = 16'b0011100110101011; 
assign lut_table[2437] = 16'b0011100110101100; 
assign lut_table[2438] = 16'b0011100110101101; 
assign lut_table[2439] = 16'b0011100110101110; 
assign lut_table[2440] = 16'b0011100110101111; 
assign lut_table[2441] = 16'b0011100110111011; 
assign lut_table[2442] = 16'b0011100110111100; 
assign lut_table[2443] = 16'b0011100110111101; 
assign lut_table[2444] = 16'b0011100110111110; 
assign lut_table[2445] = 16'b0011100110111111; 
assign lut_table[2446] = 16'b0011100111001100; 
assign lut_table[2447] = 16'b0011100111001101; 
assign lut_table[2448] = 16'b0011100111001110; 
assign lut_table[2449] = 16'b0011100111001111; 
assign lut_table[2450] = 16'b0011100111011101; 
assign lut_table[2451] = 16'b0011100111011110; 
assign lut_table[2452] = 16'b0011100111011111; 
assign lut_table[2453] = 16'b0011100111101110; 
assign lut_table[2454] = 16'b0011100111101111; 
assign lut_table[2455] = 16'b0011100111111111; 
assign lut_table[2456] = 16'b0011101010101010; 
assign lut_table[2457] = 16'b0011101010101011; 
assign lut_table[2458] = 16'b0011101010101100; 
assign lut_table[2459] = 16'b0011101010101101; 
assign lut_table[2460] = 16'b0011101010101110; 
assign lut_table[2461] = 16'b0011101010101111; 
assign lut_table[2462] = 16'b0011101010111011; 
assign lut_table[2463] = 16'b0011101010111100; 
assign lut_table[2464] = 16'b0011101010111101; 
assign lut_table[2465] = 16'b0011101010111110; 
assign lut_table[2466] = 16'b0011101010111111; 
assign lut_table[2467] = 16'b0011101011001100; 
assign lut_table[2468] = 16'b0011101011001101; 
assign lut_table[2469] = 16'b0011101011001110; 
assign lut_table[2470] = 16'b0011101011001111; 
assign lut_table[2471] = 16'b0011101011011101; 
assign lut_table[2472] = 16'b0011101011011110; 
assign lut_table[2473] = 16'b0011101011011111; 
assign lut_table[2474] = 16'b0011101011101110; 
assign lut_table[2475] = 16'b0011101011101111; 
assign lut_table[2476] = 16'b0011101011111111; 
assign lut_table[2477] = 16'b0011101110111011; 
assign lut_table[2478] = 16'b0011101110111100; 
assign lut_table[2479] = 16'b0011101110111101; 
assign lut_table[2480] = 16'b0011101110111110; 
assign lut_table[2481] = 16'b0011101110111111; 
assign lut_table[2482] = 16'b0011101111001100; 
assign lut_table[2483] = 16'b0011101111001101; 
assign lut_table[2484] = 16'b0011101111001110; 
assign lut_table[2485] = 16'b0011101111001111; 
assign lut_table[2486] = 16'b0011101111011101; 
assign lut_table[2487] = 16'b0011101111011110; 
assign lut_table[2488] = 16'b0011101111011111; 
assign lut_table[2489] = 16'b0011101111101110; 
assign lut_table[2490] = 16'b0011101111101111; 
assign lut_table[2491] = 16'b0011101111111111; 
assign lut_table[2492] = 16'b0011110011001100; 
assign lut_table[2493] = 16'b0011110011001101; 
assign lut_table[2494] = 16'b0011110011001110; 
assign lut_table[2495] = 16'b0011110011001111; 
assign lut_table[2496] = 16'b0011110011011101; 
assign lut_table[2497] = 16'b0011110011011110; 
assign lut_table[2498] = 16'b0011110011011111; 
assign lut_table[2499] = 16'b0011110011101110; 
assign lut_table[2500] = 16'b0011110011101111; 
assign lut_table[2501] = 16'b0011110011111111; 
assign lut_table[2502] = 16'b0011110111011101; 
assign lut_table[2503] = 16'b0011110111011110; 
assign lut_table[2504] = 16'b0011110111011111; 
assign lut_table[2505] = 16'b0011110111101110; 
assign lut_table[2506] = 16'b0011110111101111; 
assign lut_table[2507] = 16'b0011110111111111; 
assign lut_table[2508] = 16'b0011111011101110; 
assign lut_table[2509] = 16'b0011111011101111; 
assign lut_table[2510] = 16'b0011111011111111; 
assign lut_table[2511] = 16'b0011111111111111; 
assign lut_table[2512] = 16'b0100010001000100; 
assign lut_table[2513] = 16'b0100010001000101; 
assign lut_table[2514] = 16'b0100010001000110; 
assign lut_table[2515] = 16'b0100010001000111; 
assign lut_table[2516] = 16'b0100010001001000; 
assign lut_table[2517] = 16'b0100010001001001; 
assign lut_table[2518] = 16'b0100010001001010; 
assign lut_table[2519] = 16'b0100010001001011; 
assign lut_table[2520] = 16'b0100010001001100; 
assign lut_table[2521] = 16'b0100010001001101; 
assign lut_table[2522] = 16'b0100010001001110; 
assign lut_table[2523] = 16'b0100010001001111; 
assign lut_table[2524] = 16'b0100010001010101; 
assign lut_table[2525] = 16'b0100010001010110; 
assign lut_table[2526] = 16'b0100010001010111; 
assign lut_table[2527] = 16'b0100010001011000; 
assign lut_table[2528] = 16'b0100010001011001; 
assign lut_table[2529] = 16'b0100010001011010; 
assign lut_table[2530] = 16'b0100010001011011; 
assign lut_table[2531] = 16'b0100010001011100; 
assign lut_table[2532] = 16'b0100010001011101; 
assign lut_table[2533] = 16'b0100010001011110; 
assign lut_table[2534] = 16'b0100010001011111; 
assign lut_table[2535] = 16'b0100010001100110; 
assign lut_table[2536] = 16'b0100010001100111; 
assign lut_table[2537] = 16'b0100010001101000; 
assign lut_table[2538] = 16'b0100010001101001; 
assign lut_table[2539] = 16'b0100010001101010; 
assign lut_table[2540] = 16'b0100010001101011; 
assign lut_table[2541] = 16'b0100010001101100; 
assign lut_table[2542] = 16'b0100010001101101; 
assign lut_table[2543] = 16'b0100010001101110; 
assign lut_table[2544] = 16'b0100010001101111; 
assign lut_table[2545] = 16'b0100010001110111; 
assign lut_table[2546] = 16'b0100010001111000; 
assign lut_table[2547] = 16'b0100010001111001; 
assign lut_table[2548] = 16'b0100010001111010; 
assign lut_table[2549] = 16'b0100010001111011; 
assign lut_table[2550] = 16'b0100010001111100; 
assign lut_table[2551] = 16'b0100010001111101; 
assign lut_table[2552] = 16'b0100010001111110; 
assign lut_table[2553] = 16'b0100010001111111; 
assign lut_table[2554] = 16'b0100010010001000; 
assign lut_table[2555] = 16'b0100010010001001; 
assign lut_table[2556] = 16'b0100010010001010; 
assign lut_table[2557] = 16'b0100010010001011; 
assign lut_table[2558] = 16'b0100010010001100; 
assign lut_table[2559] = 16'b0100010010001101; 
assign lut_table[2560] = 16'b0100010010001110; 
assign lut_table[2561] = 16'b0100010010001111; 
assign lut_table[2562] = 16'b0100010010011001; 
assign lut_table[2563] = 16'b0100010010011010; 
assign lut_table[2564] = 16'b0100010010011011; 
assign lut_table[2565] = 16'b0100010010011100; 
assign lut_table[2566] = 16'b0100010010011101; 
assign lut_table[2567] = 16'b0100010010011110; 
assign lut_table[2568] = 16'b0100010010011111; 
assign lut_table[2569] = 16'b0100010010101010; 
assign lut_table[2570] = 16'b0100010010101011; 
assign lut_table[2571] = 16'b0100010010101100; 
assign lut_table[2572] = 16'b0100010010101101; 
assign lut_table[2573] = 16'b0100010010101110; 
assign lut_table[2574] = 16'b0100010010101111; 
assign lut_table[2575] = 16'b0100010010111011; 
assign lut_table[2576] = 16'b0100010010111100; 
assign lut_table[2577] = 16'b0100010010111101; 
assign lut_table[2578] = 16'b0100010010111110; 
assign lut_table[2579] = 16'b0100010010111111; 
assign lut_table[2580] = 16'b0100010011001100; 
assign lut_table[2581] = 16'b0100010011001101; 
assign lut_table[2582] = 16'b0100010011001110; 
assign lut_table[2583] = 16'b0100010011001111; 
assign lut_table[2584] = 16'b0100010011011101; 
assign lut_table[2585] = 16'b0100010011011110; 
assign lut_table[2586] = 16'b0100010011011111; 
assign lut_table[2587] = 16'b0100010011101110; 
assign lut_table[2588] = 16'b0100010011101111; 
assign lut_table[2589] = 16'b0100010011111111; 
assign lut_table[2590] = 16'b0100010101010101; 
assign lut_table[2591] = 16'b0100010101010110; 
assign lut_table[2592] = 16'b0100010101010111; 
assign lut_table[2593] = 16'b0100010101011000; 
assign lut_table[2594] = 16'b0100010101011001; 
assign lut_table[2595] = 16'b0100010101011010; 
assign lut_table[2596] = 16'b0100010101011011; 
assign lut_table[2597] = 16'b0100010101011100; 
assign lut_table[2598] = 16'b0100010101011101; 
assign lut_table[2599] = 16'b0100010101011110; 
assign lut_table[2600] = 16'b0100010101011111; 
assign lut_table[2601] = 16'b0100010101100110; 
assign lut_table[2602] = 16'b0100010101100111; 
assign lut_table[2603] = 16'b0100010101101000; 
assign lut_table[2604] = 16'b0100010101101001; 
assign lut_table[2605] = 16'b0100010101101010; 
assign lut_table[2606] = 16'b0100010101101011; 
assign lut_table[2607] = 16'b0100010101101100; 
assign lut_table[2608] = 16'b0100010101101101; 
assign lut_table[2609] = 16'b0100010101101110; 
assign lut_table[2610] = 16'b0100010101101111; 
assign lut_table[2611] = 16'b0100010101110111; 
assign lut_table[2612] = 16'b0100010101111000; 
assign lut_table[2613] = 16'b0100010101111001; 
assign lut_table[2614] = 16'b0100010101111010; 
assign lut_table[2615] = 16'b0100010101111011; 
assign lut_table[2616] = 16'b0100010101111100; 
assign lut_table[2617] = 16'b0100010101111101; 
assign lut_table[2618] = 16'b0100010101111110; 
assign lut_table[2619] = 16'b0100010101111111; 
assign lut_table[2620] = 16'b0100010110001000; 
assign lut_table[2621] = 16'b0100010110001001; 
assign lut_table[2622] = 16'b0100010110001010; 
assign lut_table[2623] = 16'b0100010110001011; 
assign lut_table[2624] = 16'b0100010110001100; 
assign lut_table[2625] = 16'b0100010110001101; 
assign lut_table[2626] = 16'b0100010110001110; 
assign lut_table[2627] = 16'b0100010110001111; 
assign lut_table[2628] = 16'b0100010110011001; 
assign lut_table[2629] = 16'b0100010110011010; 
assign lut_table[2630] = 16'b0100010110011011; 
assign lut_table[2631] = 16'b0100010110011100; 
assign lut_table[2632] = 16'b0100010110011101; 
assign lut_table[2633] = 16'b0100010110011110; 
assign lut_table[2634] = 16'b0100010110011111; 
assign lut_table[2635] = 16'b0100010110101010; 
assign lut_table[2636] = 16'b0100010110101011; 
assign lut_table[2637] = 16'b0100010110101100; 
assign lut_table[2638] = 16'b0100010110101101; 
assign lut_table[2639] = 16'b0100010110101110; 
assign lut_table[2640] = 16'b0100010110101111; 
assign lut_table[2641] = 16'b0100010110111011; 
assign lut_table[2642] = 16'b0100010110111100; 
assign lut_table[2643] = 16'b0100010110111101; 
assign lut_table[2644] = 16'b0100010110111110; 
assign lut_table[2645] = 16'b0100010110111111; 
assign lut_table[2646] = 16'b0100010111001100; 
assign lut_table[2647] = 16'b0100010111001101; 
assign lut_table[2648] = 16'b0100010111001110; 
assign lut_table[2649] = 16'b0100010111001111; 
assign lut_table[2650] = 16'b0100010111011101; 
assign lut_table[2651] = 16'b0100010111011110; 
assign lut_table[2652] = 16'b0100010111011111; 
assign lut_table[2653] = 16'b0100010111101110; 
assign lut_table[2654] = 16'b0100010111101111; 
assign lut_table[2655] = 16'b0100010111111111; 
assign lut_table[2656] = 16'b0100011001100110; 
assign lut_table[2657] = 16'b0100011001100111; 
assign lut_table[2658] = 16'b0100011001101000; 
assign lut_table[2659] = 16'b0100011001101001; 
assign lut_table[2660] = 16'b0100011001101010; 
assign lut_table[2661] = 16'b0100011001101011; 
assign lut_table[2662] = 16'b0100011001101100; 
assign lut_table[2663] = 16'b0100011001101101; 
assign lut_table[2664] = 16'b0100011001101110; 
assign lut_table[2665] = 16'b0100011001101111; 
assign lut_table[2666] = 16'b0100011001110111; 
assign lut_table[2667] = 16'b0100011001111000; 
assign lut_table[2668] = 16'b0100011001111001; 
assign lut_table[2669] = 16'b0100011001111010; 
assign lut_table[2670] = 16'b0100011001111011; 
assign lut_table[2671] = 16'b0100011001111100; 
assign lut_table[2672] = 16'b0100011001111101; 
assign lut_table[2673] = 16'b0100011001111110; 
assign lut_table[2674] = 16'b0100011001111111; 
assign lut_table[2675] = 16'b0100011010001000; 
assign lut_table[2676] = 16'b0100011010001001; 
assign lut_table[2677] = 16'b0100011010001010; 
assign lut_table[2678] = 16'b0100011010001011; 
assign lut_table[2679] = 16'b0100011010001100; 
assign lut_table[2680] = 16'b0100011010001101; 
assign lut_table[2681] = 16'b0100011010001110; 
assign lut_table[2682] = 16'b0100011010001111; 
assign lut_table[2683] = 16'b0100011010011001; 
assign lut_table[2684] = 16'b0100011010011010; 
assign lut_table[2685] = 16'b0100011010011011; 
assign lut_table[2686] = 16'b0100011010011100; 
assign lut_table[2687] = 16'b0100011010011101; 
assign lut_table[2688] = 16'b0100011010011110; 
assign lut_table[2689] = 16'b0100011010011111; 
assign lut_table[2690] = 16'b0100011010101010; 
assign lut_table[2691] = 16'b0100011010101011; 
assign lut_table[2692] = 16'b0100011010101100; 
assign lut_table[2693] = 16'b0100011010101101; 
assign lut_table[2694] = 16'b0100011010101110; 
assign lut_table[2695] = 16'b0100011010101111; 
assign lut_table[2696] = 16'b0100011010111011; 
assign lut_table[2697] = 16'b0100011010111100; 
assign lut_table[2698] = 16'b0100011010111101; 
assign lut_table[2699] = 16'b0100011010111110; 
assign lut_table[2700] = 16'b0100011010111111; 
assign lut_table[2701] = 16'b0100011011001100; 
assign lut_table[2702] = 16'b0100011011001101; 
assign lut_table[2703] = 16'b0100011011001110; 
assign lut_table[2704] = 16'b0100011011001111; 
assign lut_table[2705] = 16'b0100011011011101; 
assign lut_table[2706] = 16'b0100011011011110; 
assign lut_table[2707] = 16'b0100011011011111; 
assign lut_table[2708] = 16'b0100011011101110; 
assign lut_table[2709] = 16'b0100011011101111; 
assign lut_table[2710] = 16'b0100011011111111; 
assign lut_table[2711] = 16'b0100011101110111; 
assign lut_table[2712] = 16'b0100011101111000; 
assign lut_table[2713] = 16'b0100011101111001; 
assign lut_table[2714] = 16'b0100011101111010; 
assign lut_table[2715] = 16'b0100011101111011; 
assign lut_table[2716] = 16'b0100011101111100; 
assign lut_table[2717] = 16'b0100011101111101; 
assign lut_table[2718] = 16'b0100011101111110; 
assign lut_table[2719] = 16'b0100011101111111; 
assign lut_table[2720] = 16'b0100011110001000; 
assign lut_table[2721] = 16'b0100011110001001; 
assign lut_table[2722] = 16'b0100011110001010; 
assign lut_table[2723] = 16'b0100011110001011; 
assign lut_table[2724] = 16'b0100011110001100; 
assign lut_table[2725] = 16'b0100011110001101; 
assign lut_table[2726] = 16'b0100011110001110; 
assign lut_table[2727] = 16'b0100011110001111; 
assign lut_table[2728] = 16'b0100011110011001; 
assign lut_table[2729] = 16'b0100011110011010; 
assign lut_table[2730] = 16'b0100011110011011; 
assign lut_table[2731] = 16'b0100011110011100; 
assign lut_table[2732] = 16'b0100011110011101; 
assign lut_table[2733] = 16'b0100011110011110; 
assign lut_table[2734] = 16'b0100011110011111; 
assign lut_table[2735] = 16'b0100011110101010; 
assign lut_table[2736] = 16'b0100011110101011; 
assign lut_table[2737] = 16'b0100011110101100; 
assign lut_table[2738] = 16'b0100011110101101; 
assign lut_table[2739] = 16'b0100011110101110; 
assign lut_table[2740] = 16'b0100011110101111; 
assign lut_table[2741] = 16'b0100011110111011; 
assign lut_table[2742] = 16'b0100011110111100; 
assign lut_table[2743] = 16'b0100011110111101; 
assign lut_table[2744] = 16'b0100011110111110; 
assign lut_table[2745] = 16'b0100011110111111; 
assign lut_table[2746] = 16'b0100011111001100; 
assign lut_table[2747] = 16'b0100011111001101; 
assign lut_table[2748] = 16'b0100011111001110; 
assign lut_table[2749] = 16'b0100011111001111; 
assign lut_table[2750] = 16'b0100011111011101; 
assign lut_table[2751] = 16'b0100011111011110; 
assign lut_table[2752] = 16'b0100011111011111; 
assign lut_table[2753] = 16'b0100011111101110; 
assign lut_table[2754] = 16'b0100011111101111; 
assign lut_table[2755] = 16'b0100011111111111; 
assign lut_table[2756] = 16'b0100100010001000; 
assign lut_table[2757] = 16'b0100100010001001; 
assign lut_table[2758] = 16'b0100100010001010; 
assign lut_table[2759] = 16'b0100100010001011; 
assign lut_table[2760] = 16'b0100100010001100; 
assign lut_table[2761] = 16'b0100100010001101; 
assign lut_table[2762] = 16'b0100100010001110; 
assign lut_table[2763] = 16'b0100100010001111; 
assign lut_table[2764] = 16'b0100100010011001; 
assign lut_table[2765] = 16'b0100100010011010; 
assign lut_table[2766] = 16'b0100100010011011; 
assign lut_table[2767] = 16'b0100100010011100; 
assign lut_table[2768] = 16'b0100100010011101; 
assign lut_table[2769] = 16'b0100100010011110; 
assign lut_table[2770] = 16'b0100100010011111; 
assign lut_table[2771] = 16'b0100100010101010; 
assign lut_table[2772] = 16'b0100100010101011; 
assign lut_table[2773] = 16'b0100100010101100; 
assign lut_table[2774] = 16'b0100100010101101; 
assign lut_table[2775] = 16'b0100100010101110; 
assign lut_table[2776] = 16'b0100100010101111; 
assign lut_table[2777] = 16'b0100100010111011; 
assign lut_table[2778] = 16'b0100100010111100; 
assign lut_table[2779] = 16'b0100100010111101; 
assign lut_table[2780] = 16'b0100100010111110; 
assign lut_table[2781] = 16'b0100100010111111; 
assign lut_table[2782] = 16'b0100100011001100; 
assign lut_table[2783] = 16'b0100100011001101; 
assign lut_table[2784] = 16'b0100100011001110; 
assign lut_table[2785] = 16'b0100100011001111; 
assign lut_table[2786] = 16'b0100100011011101; 
assign lut_table[2787] = 16'b0100100011011110; 
assign lut_table[2788] = 16'b0100100011011111; 
assign lut_table[2789] = 16'b0100100011101110; 
assign lut_table[2790] = 16'b0100100011101111; 
assign lut_table[2791] = 16'b0100100011111111; 
assign lut_table[2792] = 16'b0100100110011001; 
assign lut_table[2793] = 16'b0100100110011010; 
assign lut_table[2794] = 16'b0100100110011011; 
assign lut_table[2795] = 16'b0100100110011100; 
assign lut_table[2796] = 16'b0100100110011101; 
assign lut_table[2797] = 16'b0100100110011110; 
assign lut_table[2798] = 16'b0100100110011111; 
assign lut_table[2799] = 16'b0100100110101010; 
assign lut_table[2800] = 16'b0100100110101011; 
assign lut_table[2801] = 16'b0100100110101100; 
assign lut_table[2802] = 16'b0100100110101101; 
assign lut_table[2803] = 16'b0100100110101110; 
assign lut_table[2804] = 16'b0100100110101111; 
assign lut_table[2805] = 16'b0100100110111011; 
assign lut_table[2806] = 16'b0100100110111100; 
assign lut_table[2807] = 16'b0100100110111101; 
assign lut_table[2808] = 16'b0100100110111110; 
assign lut_table[2809] = 16'b0100100110111111; 
assign lut_table[2810] = 16'b0100100111001100; 
assign lut_table[2811] = 16'b0100100111001101; 
assign lut_table[2812] = 16'b0100100111001110; 
assign lut_table[2813] = 16'b0100100111001111; 
assign lut_table[2814] = 16'b0100100111011101; 
assign lut_table[2815] = 16'b0100100111011110; 
assign lut_table[2816] = 16'b0100100111011111; 
assign lut_table[2817] = 16'b0100100111101110; 
assign lut_table[2818] = 16'b0100100111101111; 
assign lut_table[2819] = 16'b0100100111111111; 
assign lut_table[2820] = 16'b0100101010101010; 
assign lut_table[2821] = 16'b0100101010101011; 
assign lut_table[2822] = 16'b0100101010101100; 
assign lut_table[2823] = 16'b0100101010101101; 
assign lut_table[2824] = 16'b0100101010101110; 
assign lut_table[2825] = 16'b0100101010101111; 
assign lut_table[2826] = 16'b0100101010111011; 
assign lut_table[2827] = 16'b0100101010111100; 
assign lut_table[2828] = 16'b0100101010111101; 
assign lut_table[2829] = 16'b0100101010111110; 
assign lut_table[2830] = 16'b0100101010111111; 
assign lut_table[2831] = 16'b0100101011001100; 
assign lut_table[2832] = 16'b0100101011001101; 
assign lut_table[2833] = 16'b0100101011001110; 
assign lut_table[2834] = 16'b0100101011001111; 
assign lut_table[2835] = 16'b0100101011011101; 
assign lut_table[2836] = 16'b0100101011011110; 
assign lut_table[2837] = 16'b0100101011011111; 
assign lut_table[2838] = 16'b0100101011101110; 
assign lut_table[2839] = 16'b0100101011101111; 
assign lut_table[2840] = 16'b0100101011111111; 
assign lut_table[2841] = 16'b0100101110111011; 
assign lut_table[2842] = 16'b0100101110111100; 
assign lut_table[2843] = 16'b0100101110111101; 
assign lut_table[2844] = 16'b0100101110111110; 
assign lut_table[2845] = 16'b0100101110111111; 
assign lut_table[2846] = 16'b0100101111001100; 
assign lut_table[2847] = 16'b0100101111001101; 
assign lut_table[2848] = 16'b0100101111001110; 
assign lut_table[2849] = 16'b0100101111001111; 
assign lut_table[2850] = 16'b0100101111011101; 
assign lut_table[2851] = 16'b0100101111011110; 
assign lut_table[2852] = 16'b0100101111011111; 
assign lut_table[2853] = 16'b0100101111101110; 
assign lut_table[2854] = 16'b0100101111101111; 
assign lut_table[2855] = 16'b0100101111111111; 
assign lut_table[2856] = 16'b0100110011001100; 
assign lut_table[2857] = 16'b0100110011001101; 
assign lut_table[2858] = 16'b0100110011001110; 
assign lut_table[2859] = 16'b0100110011001111; 
assign lut_table[2860] = 16'b0100110011011101; 
assign lut_table[2861] = 16'b0100110011011110; 
assign lut_table[2862] = 16'b0100110011011111; 
assign lut_table[2863] = 16'b0100110011101110; 
assign lut_table[2864] = 16'b0100110011101111; 
assign lut_table[2865] = 16'b0100110011111111; 
assign lut_table[2866] = 16'b0100110111011101; 
assign lut_table[2867] = 16'b0100110111011110; 
assign lut_table[2868] = 16'b0100110111011111; 
assign lut_table[2869] = 16'b0100110111101110; 
assign lut_table[2870] = 16'b0100110111101111; 
assign lut_table[2871] = 16'b0100110111111111; 
assign lut_table[2872] = 16'b0100111011101110; 
assign lut_table[2873] = 16'b0100111011101111; 
assign lut_table[2874] = 16'b0100111011111111; 
assign lut_table[2875] = 16'b0100111111111111; 
assign lut_table[2876] = 16'b0101010101010101; 
assign lut_table[2877] = 16'b0101010101010110; 
assign lut_table[2878] = 16'b0101010101010111; 
assign lut_table[2879] = 16'b0101010101011000; 
assign lut_table[2880] = 16'b0101010101011001; 
assign lut_table[2881] = 16'b0101010101011010; 
assign lut_table[2882] = 16'b0101010101011011; 
assign lut_table[2883] = 16'b0101010101011100; 
assign lut_table[2884] = 16'b0101010101011101; 
assign lut_table[2885] = 16'b0101010101011110; 
assign lut_table[2886] = 16'b0101010101011111; 
assign lut_table[2887] = 16'b0101010101100110; 
assign lut_table[2888] = 16'b0101010101100111; 
assign lut_table[2889] = 16'b0101010101101000; 
assign lut_table[2890] = 16'b0101010101101001; 
assign lut_table[2891] = 16'b0101010101101010; 
assign lut_table[2892] = 16'b0101010101101011; 
assign lut_table[2893] = 16'b0101010101101100; 
assign lut_table[2894] = 16'b0101010101101101; 
assign lut_table[2895] = 16'b0101010101101110; 
assign lut_table[2896] = 16'b0101010101101111; 
assign lut_table[2897] = 16'b0101010101110111; 
assign lut_table[2898] = 16'b0101010101111000; 
assign lut_table[2899] = 16'b0101010101111001; 
assign lut_table[2900] = 16'b0101010101111010; 
assign lut_table[2901] = 16'b0101010101111011; 
assign lut_table[2902] = 16'b0101010101111100; 
assign lut_table[2903] = 16'b0101010101111101; 
assign lut_table[2904] = 16'b0101010101111110; 
assign lut_table[2905] = 16'b0101010101111111; 
assign lut_table[2906] = 16'b0101010110001000; 
assign lut_table[2907] = 16'b0101010110001001; 
assign lut_table[2908] = 16'b0101010110001010; 
assign lut_table[2909] = 16'b0101010110001011; 
assign lut_table[2910] = 16'b0101010110001100; 
assign lut_table[2911] = 16'b0101010110001101; 
assign lut_table[2912] = 16'b0101010110001110; 
assign lut_table[2913] = 16'b0101010110001111; 
assign lut_table[2914] = 16'b0101010110011001; 
assign lut_table[2915] = 16'b0101010110011010; 
assign lut_table[2916] = 16'b0101010110011011; 
assign lut_table[2917] = 16'b0101010110011100; 
assign lut_table[2918] = 16'b0101010110011101; 
assign lut_table[2919] = 16'b0101010110011110; 
assign lut_table[2920] = 16'b0101010110011111; 
assign lut_table[2921] = 16'b0101010110101010; 
assign lut_table[2922] = 16'b0101010110101011; 
assign lut_table[2923] = 16'b0101010110101100; 
assign lut_table[2924] = 16'b0101010110101101; 
assign lut_table[2925] = 16'b0101010110101110; 
assign lut_table[2926] = 16'b0101010110101111; 
assign lut_table[2927] = 16'b0101010110111011; 
assign lut_table[2928] = 16'b0101010110111100; 
assign lut_table[2929] = 16'b0101010110111101; 
assign lut_table[2930] = 16'b0101010110111110; 
assign lut_table[2931] = 16'b0101010110111111; 
assign lut_table[2932] = 16'b0101010111001100; 
assign lut_table[2933] = 16'b0101010111001101; 
assign lut_table[2934] = 16'b0101010111001110; 
assign lut_table[2935] = 16'b0101010111001111; 
assign lut_table[2936] = 16'b0101010111011101; 
assign lut_table[2937] = 16'b0101010111011110; 
assign lut_table[2938] = 16'b0101010111011111; 
assign lut_table[2939] = 16'b0101010111101110; 
assign lut_table[2940] = 16'b0101010111101111; 
assign lut_table[2941] = 16'b0101010111111111; 
assign lut_table[2942] = 16'b0101011001100110; 
assign lut_table[2943] = 16'b0101011001100111; 
assign lut_table[2944] = 16'b0101011001101000; 
assign lut_table[2945] = 16'b0101011001101001; 
assign lut_table[2946] = 16'b0101011001101010; 
assign lut_table[2947] = 16'b0101011001101011; 
assign lut_table[2948] = 16'b0101011001101100; 
assign lut_table[2949] = 16'b0101011001101101; 
assign lut_table[2950] = 16'b0101011001101110; 
assign lut_table[2951] = 16'b0101011001101111; 
assign lut_table[2952] = 16'b0101011001110111; 
assign lut_table[2953] = 16'b0101011001111000; 
assign lut_table[2954] = 16'b0101011001111001; 
assign lut_table[2955] = 16'b0101011001111010; 
assign lut_table[2956] = 16'b0101011001111011; 
assign lut_table[2957] = 16'b0101011001111100; 
assign lut_table[2958] = 16'b0101011001111101; 
assign lut_table[2959] = 16'b0101011001111110; 
assign lut_table[2960] = 16'b0101011001111111; 
assign lut_table[2961] = 16'b0101011010001000; 
assign lut_table[2962] = 16'b0101011010001001; 
assign lut_table[2963] = 16'b0101011010001010; 
assign lut_table[2964] = 16'b0101011010001011; 
assign lut_table[2965] = 16'b0101011010001100; 
assign lut_table[2966] = 16'b0101011010001101; 
assign lut_table[2967] = 16'b0101011010001110; 
assign lut_table[2968] = 16'b0101011010001111; 
assign lut_table[2969] = 16'b0101011010011001; 
assign lut_table[2970] = 16'b0101011010011010; 
assign lut_table[2971] = 16'b0101011010011011; 
assign lut_table[2972] = 16'b0101011010011100; 
assign lut_table[2973] = 16'b0101011010011101; 
assign lut_table[2974] = 16'b0101011010011110; 
assign lut_table[2975] = 16'b0101011010011111; 
assign lut_table[2976] = 16'b0101011010101010; 
assign lut_table[2977] = 16'b0101011010101011; 
assign lut_table[2978] = 16'b0101011010101100; 
assign lut_table[2979] = 16'b0101011010101101; 
assign lut_table[2980] = 16'b0101011010101110; 
assign lut_table[2981] = 16'b0101011010101111; 
assign lut_table[2982] = 16'b0101011010111011; 
assign lut_table[2983] = 16'b0101011010111100; 
assign lut_table[2984] = 16'b0101011010111101; 
assign lut_table[2985] = 16'b0101011010111110; 
assign lut_table[2986] = 16'b0101011010111111; 
assign lut_table[2987] = 16'b0101011011001100; 
assign lut_table[2988] = 16'b0101011011001101; 
assign lut_table[2989] = 16'b0101011011001110; 
assign lut_table[2990] = 16'b0101011011001111; 
assign lut_table[2991] = 16'b0101011011011101; 
assign lut_table[2992] = 16'b0101011011011110; 
assign lut_table[2993] = 16'b0101011011011111; 
assign lut_table[2994] = 16'b0101011011101110; 
assign lut_table[2995] = 16'b0101011011101111; 
assign lut_table[2996] = 16'b0101011011111111; 
assign lut_table[2997] = 16'b0101011101110111; 
assign lut_table[2998] = 16'b0101011101111000; 
assign lut_table[2999] = 16'b0101011101111001; 
assign lut_table[3000] = 16'b0101011101111010; 
assign lut_table[3001] = 16'b0101011101111011; 
assign lut_table[3002] = 16'b0101011101111100; 
assign lut_table[3003] = 16'b0101011101111101; 
assign lut_table[3004] = 16'b0101011101111110; 
assign lut_table[3005] = 16'b0101011101111111; 
assign lut_table[3006] = 16'b0101011110001000; 
assign lut_table[3007] = 16'b0101011110001001; 
assign lut_table[3008] = 16'b0101011110001010; 
assign lut_table[3009] = 16'b0101011110001011; 
assign lut_table[3010] = 16'b0101011110001100; 
assign lut_table[3011] = 16'b0101011110001101; 
assign lut_table[3012] = 16'b0101011110001110; 
assign lut_table[3013] = 16'b0101011110001111; 
assign lut_table[3014] = 16'b0101011110011001; 
assign lut_table[3015] = 16'b0101011110011010; 
assign lut_table[3016] = 16'b0101011110011011; 
assign lut_table[3017] = 16'b0101011110011100; 
assign lut_table[3018] = 16'b0101011110011101; 
assign lut_table[3019] = 16'b0101011110011110; 
assign lut_table[3020] = 16'b0101011110011111; 
assign lut_table[3021] = 16'b0101011110101010; 
assign lut_table[3022] = 16'b0101011110101011; 
assign lut_table[3023] = 16'b0101011110101100; 
assign lut_table[3024] = 16'b0101011110101101; 
assign lut_table[3025] = 16'b0101011110101110; 
assign lut_table[3026] = 16'b0101011110101111; 
assign lut_table[3027] = 16'b0101011110111011; 
assign lut_table[3028] = 16'b0101011110111100; 
assign lut_table[3029] = 16'b0101011110111101; 
assign lut_table[3030] = 16'b0101011110111110; 
assign lut_table[3031] = 16'b0101011110111111; 
assign lut_table[3032] = 16'b0101011111001100; 
assign lut_table[3033] = 16'b0101011111001101; 
assign lut_table[3034] = 16'b0101011111001110; 
assign lut_table[3035] = 16'b0101011111001111; 
assign lut_table[3036] = 16'b0101011111011101; 
assign lut_table[3037] = 16'b0101011111011110; 
assign lut_table[3038] = 16'b0101011111011111; 
assign lut_table[3039] = 16'b0101011111101110; 
assign lut_table[3040] = 16'b0101011111101111; 
assign lut_table[3041] = 16'b0101011111111111; 
assign lut_table[3042] = 16'b0101100010001000; 
assign lut_table[3043] = 16'b0101100010001001; 
assign lut_table[3044] = 16'b0101100010001010; 
assign lut_table[3045] = 16'b0101100010001011; 
assign lut_table[3046] = 16'b0101100010001100; 
assign lut_table[3047] = 16'b0101100010001101; 
assign lut_table[3048] = 16'b0101100010001110; 
assign lut_table[3049] = 16'b0101100010001111; 
assign lut_table[3050] = 16'b0101100010011001; 
assign lut_table[3051] = 16'b0101100010011010; 
assign lut_table[3052] = 16'b0101100010011011; 
assign lut_table[3053] = 16'b0101100010011100; 
assign lut_table[3054] = 16'b0101100010011101; 
assign lut_table[3055] = 16'b0101100010011110; 
assign lut_table[3056] = 16'b0101100010011111; 
assign lut_table[3057] = 16'b0101100010101010; 
assign lut_table[3058] = 16'b0101100010101011; 
assign lut_table[3059] = 16'b0101100010101100; 
assign lut_table[3060] = 16'b0101100010101101; 
assign lut_table[3061] = 16'b0101100010101110; 
assign lut_table[3062] = 16'b0101100010101111; 
assign lut_table[3063] = 16'b0101100010111011; 
assign lut_table[3064] = 16'b0101100010111100; 
assign lut_table[3065] = 16'b0101100010111101; 
assign lut_table[3066] = 16'b0101100010111110; 
assign lut_table[3067] = 16'b0101100010111111; 
assign lut_table[3068] = 16'b0101100011001100; 
assign lut_table[3069] = 16'b0101100011001101; 
assign lut_table[3070] = 16'b0101100011001110; 
assign lut_table[3071] = 16'b0101100011001111; 
assign lut_table[3072] = 16'b0101100011011101; 
assign lut_table[3073] = 16'b0101100011011110; 
assign lut_table[3074] = 16'b0101100011011111; 
assign lut_table[3075] = 16'b0101100011101110; 
assign lut_table[3076] = 16'b0101100011101111; 
assign lut_table[3077] = 16'b0101100011111111; 
assign lut_table[3078] = 16'b0101100110011001; 
assign lut_table[3079] = 16'b0101100110011010; 
assign lut_table[3080] = 16'b0101100110011011; 
assign lut_table[3081] = 16'b0101100110011100; 
assign lut_table[3082] = 16'b0101100110011101; 
assign lut_table[3083] = 16'b0101100110011110; 
assign lut_table[3084] = 16'b0101100110011111; 
assign lut_table[3085] = 16'b0101100110101010; 
assign lut_table[3086] = 16'b0101100110101011; 
assign lut_table[3087] = 16'b0101100110101100; 
assign lut_table[3088] = 16'b0101100110101101; 
assign lut_table[3089] = 16'b0101100110101110; 
assign lut_table[3090] = 16'b0101100110101111; 
assign lut_table[3091] = 16'b0101100110111011; 
assign lut_table[3092] = 16'b0101100110111100; 
assign lut_table[3093] = 16'b0101100110111101; 
assign lut_table[3094] = 16'b0101100110111110; 
assign lut_table[3095] = 16'b0101100110111111; 
assign lut_table[3096] = 16'b0101100111001100; 
assign lut_table[3097] = 16'b0101100111001101; 
assign lut_table[3098] = 16'b0101100111001110; 
assign lut_table[3099] = 16'b0101100111001111; 
assign lut_table[3100] = 16'b0101100111011101; 
assign lut_table[3101] = 16'b0101100111011110; 
assign lut_table[3102] = 16'b0101100111011111; 
assign lut_table[3103] = 16'b0101100111101110; 
assign lut_table[3104] = 16'b0101100111101111; 
assign lut_table[3105] = 16'b0101100111111111; 
assign lut_table[3106] = 16'b0101101010101010; 
assign lut_table[3107] = 16'b0101101010101011; 
assign lut_table[3108] = 16'b0101101010101100; 
assign lut_table[3109] = 16'b0101101010101101; 
assign lut_table[3110] = 16'b0101101010101110; 
assign lut_table[3111] = 16'b0101101010101111; 
assign lut_table[3112] = 16'b0101101010111011; 
assign lut_table[3113] = 16'b0101101010111100; 
assign lut_table[3114] = 16'b0101101010111101; 
assign lut_table[3115] = 16'b0101101010111110; 
assign lut_table[3116] = 16'b0101101010111111; 
assign lut_table[3117] = 16'b0101101011001100; 
assign lut_table[3118] = 16'b0101101011001101; 
assign lut_table[3119] = 16'b0101101011001110; 
assign lut_table[3120] = 16'b0101101011001111; 
assign lut_table[3121] = 16'b0101101011011101; 
assign lut_table[3122] = 16'b0101101011011110; 
assign lut_table[3123] = 16'b0101101011011111; 
assign lut_table[3124] = 16'b0101101011101110; 
assign lut_table[3125] = 16'b0101101011101111; 
assign lut_table[3126] = 16'b0101101011111111; 
assign lut_table[3127] = 16'b0101101110111011; 
assign lut_table[3128] = 16'b0101101110111100; 
assign lut_table[3129] = 16'b0101101110111101; 
assign lut_table[3130] = 16'b0101101110111110; 
assign lut_table[3131] = 16'b0101101110111111; 
assign lut_table[3132] = 16'b0101101111001100; 
assign lut_table[3133] = 16'b0101101111001101; 
assign lut_table[3134] = 16'b0101101111001110; 
assign lut_table[3135] = 16'b0101101111001111; 
assign lut_table[3136] = 16'b0101101111011101; 
assign lut_table[3137] = 16'b0101101111011110; 
assign lut_table[3138] = 16'b0101101111011111; 
assign lut_table[3139] = 16'b0101101111101110; 
assign lut_table[3140] = 16'b0101101111101111; 
assign lut_table[3141] = 16'b0101101111111111; 
assign lut_table[3142] = 16'b0101110011001100; 
assign lut_table[3143] = 16'b0101110011001101; 
assign lut_table[3144] = 16'b0101110011001110; 
assign lut_table[3145] = 16'b0101110011001111; 
assign lut_table[3146] = 16'b0101110011011101; 
assign lut_table[3147] = 16'b0101110011011110; 
assign lut_table[3148] = 16'b0101110011011111; 
assign lut_table[3149] = 16'b0101110011101110; 
assign lut_table[3150] = 16'b0101110011101111; 
assign lut_table[3151] = 16'b0101110011111111; 
assign lut_table[3152] = 16'b0101110111011101; 
assign lut_table[3153] = 16'b0101110111011110; 
assign lut_table[3154] = 16'b0101110111011111; 
assign lut_table[3155] = 16'b0101110111101110; 
assign lut_table[3156] = 16'b0101110111101111; 
assign lut_table[3157] = 16'b0101110111111111; 
assign lut_table[3158] = 16'b0101111011101110; 
assign lut_table[3159] = 16'b0101111011101111; 
assign lut_table[3160] = 16'b0101111011111111; 
assign lut_table[3161] = 16'b0101111111111111; 
assign lut_table[3162] = 16'b0110011001100110; 
assign lut_table[3163] = 16'b0110011001100111; 
assign lut_table[3164] = 16'b0110011001101000; 
assign lut_table[3165] = 16'b0110011001101001; 
assign lut_table[3166] = 16'b0110011001101010; 
assign lut_table[3167] = 16'b0110011001101011; 
assign lut_table[3168] = 16'b0110011001101100; 
assign lut_table[3169] = 16'b0110011001101101; 
assign lut_table[3170] = 16'b0110011001101110; 
assign lut_table[3171] = 16'b0110011001101111; 
assign lut_table[3172] = 16'b0110011001110111; 
assign lut_table[3173] = 16'b0110011001111000; 
assign lut_table[3174] = 16'b0110011001111001; 
assign lut_table[3175] = 16'b0110011001111010; 
assign lut_table[3176] = 16'b0110011001111011; 
assign lut_table[3177] = 16'b0110011001111100; 
assign lut_table[3178] = 16'b0110011001111101; 
assign lut_table[3179] = 16'b0110011001111110; 
assign lut_table[3180] = 16'b0110011001111111; 
assign lut_table[3181] = 16'b0110011010001000; 
assign lut_table[3182] = 16'b0110011010001001; 
assign lut_table[3183] = 16'b0110011010001010; 
assign lut_table[3184] = 16'b0110011010001011; 
assign lut_table[3185] = 16'b0110011010001100; 
assign lut_table[3186] = 16'b0110011010001101; 
assign lut_table[3187] = 16'b0110011010001110; 
assign lut_table[3188] = 16'b0110011010001111; 
assign lut_table[3189] = 16'b0110011010011001; 
assign lut_table[3190] = 16'b0110011010011010; 
assign lut_table[3191] = 16'b0110011010011011; 
assign lut_table[3192] = 16'b0110011010011100; 
assign lut_table[3193] = 16'b0110011010011101; 
assign lut_table[3194] = 16'b0110011010011110; 
assign lut_table[3195] = 16'b0110011010011111; 
assign lut_table[3196] = 16'b0110011010101010; 
assign lut_table[3197] = 16'b0110011010101011; 
assign lut_table[3198] = 16'b0110011010101100; 
assign lut_table[3199] = 16'b0110011010101101; 
assign lut_table[3200] = 16'b0110011010101110; 
assign lut_table[3201] = 16'b0110011010101111; 
assign lut_table[3202] = 16'b0110011010111011; 
assign lut_table[3203] = 16'b0110011010111100; 
assign lut_table[3204] = 16'b0110011010111101; 
assign lut_table[3205] = 16'b0110011010111110; 
assign lut_table[3206] = 16'b0110011010111111; 
assign lut_table[3207] = 16'b0110011011001100; 
assign lut_table[3208] = 16'b0110011011001101; 
assign lut_table[3209] = 16'b0110011011001110; 
assign lut_table[3210] = 16'b0110011011001111; 
assign lut_table[3211] = 16'b0110011011011101; 
assign lut_table[3212] = 16'b0110011011011110; 
assign lut_table[3213] = 16'b0110011011011111; 
assign lut_table[3214] = 16'b0110011011101110; 
assign lut_table[3215] = 16'b0110011011101111; 
assign lut_table[3216] = 16'b0110011011111111; 
assign lut_table[3217] = 16'b0110011101110111; 
assign lut_table[3218] = 16'b0110011101111000; 
assign lut_table[3219] = 16'b0110011101111001; 
assign lut_table[3220] = 16'b0110011101111010; 
assign lut_table[3221] = 16'b0110011101111011; 
assign lut_table[3222] = 16'b0110011101111100; 
assign lut_table[3223] = 16'b0110011101111101; 
assign lut_table[3224] = 16'b0110011101111110; 
assign lut_table[3225] = 16'b0110011101111111; 
assign lut_table[3226] = 16'b0110011110001000; 
assign lut_table[3227] = 16'b0110011110001001; 
assign lut_table[3228] = 16'b0110011110001010; 
assign lut_table[3229] = 16'b0110011110001011; 
assign lut_table[3230] = 16'b0110011110001100; 
assign lut_table[3231] = 16'b0110011110001101; 
assign lut_table[3232] = 16'b0110011110001110; 
assign lut_table[3233] = 16'b0110011110001111; 
assign lut_table[3234] = 16'b0110011110011001; 
assign lut_table[3235] = 16'b0110011110011010; 
assign lut_table[3236] = 16'b0110011110011011; 
assign lut_table[3237] = 16'b0110011110011100; 
assign lut_table[3238] = 16'b0110011110011101; 
assign lut_table[3239] = 16'b0110011110011110; 
assign lut_table[3240] = 16'b0110011110011111; 
assign lut_table[3241] = 16'b0110011110101010; 
assign lut_table[3242] = 16'b0110011110101011; 
assign lut_table[3243] = 16'b0110011110101100; 
assign lut_table[3244] = 16'b0110011110101101; 
assign lut_table[3245] = 16'b0110011110101110; 
assign lut_table[3246] = 16'b0110011110101111; 
assign lut_table[3247] = 16'b0110011110111011; 
assign lut_table[3248] = 16'b0110011110111100; 
assign lut_table[3249] = 16'b0110011110111101; 
assign lut_table[3250] = 16'b0110011110111110; 
assign lut_table[3251] = 16'b0110011110111111; 
assign lut_table[3252] = 16'b0110011111001100; 
assign lut_table[3253] = 16'b0110011111001101; 
assign lut_table[3254] = 16'b0110011111001110; 
assign lut_table[3255] = 16'b0110011111001111; 
assign lut_table[3256] = 16'b0110011111011101; 
assign lut_table[3257] = 16'b0110011111011110; 
assign lut_table[3258] = 16'b0110011111011111; 
assign lut_table[3259] = 16'b0110011111101110; 
assign lut_table[3260] = 16'b0110011111101111; 
assign lut_table[3261] = 16'b0110011111111111; 
assign lut_table[3262] = 16'b0110100010001000; 
assign lut_table[3263] = 16'b0110100010001001; 
assign lut_table[3264] = 16'b0110100010001010; 
assign lut_table[3265] = 16'b0110100010001011; 
assign lut_table[3266] = 16'b0110100010001100; 
assign lut_table[3267] = 16'b0110100010001101; 
assign lut_table[3268] = 16'b0110100010001110; 
assign lut_table[3269] = 16'b0110100010001111; 
assign lut_table[3270] = 16'b0110100010011001; 
assign lut_table[3271] = 16'b0110100010011010; 
assign lut_table[3272] = 16'b0110100010011011; 
assign lut_table[3273] = 16'b0110100010011100; 
assign lut_table[3274] = 16'b0110100010011101; 
assign lut_table[3275] = 16'b0110100010011110; 
assign lut_table[3276] = 16'b0110100010011111; 
assign lut_table[3277] = 16'b0110100010101010; 
assign lut_table[3278] = 16'b0110100010101011; 
assign lut_table[3279] = 16'b0110100010101100; 
assign lut_table[3280] = 16'b0110100010101101; 
assign lut_table[3281] = 16'b0110100010101110; 
assign lut_table[3282] = 16'b0110100010101111; 
assign lut_table[3283] = 16'b0110100010111011; 
assign lut_table[3284] = 16'b0110100010111100; 
assign lut_table[3285] = 16'b0110100010111101; 
assign lut_table[3286] = 16'b0110100010111110; 
assign lut_table[3287] = 16'b0110100010111111; 
assign lut_table[3288] = 16'b0110100011001100; 
assign lut_table[3289] = 16'b0110100011001101; 
assign lut_table[3290] = 16'b0110100011001110; 
assign lut_table[3291] = 16'b0110100011001111; 
assign lut_table[3292] = 16'b0110100011011101; 
assign lut_table[3293] = 16'b0110100011011110; 
assign lut_table[3294] = 16'b0110100011011111; 
assign lut_table[3295] = 16'b0110100011101110; 
assign lut_table[3296] = 16'b0110100011101111; 
assign lut_table[3297] = 16'b0110100011111111; 
assign lut_table[3298] = 16'b0110100110011001; 
assign lut_table[3299] = 16'b0110100110011010; 
assign lut_table[3300] = 16'b0110100110011011; 
assign lut_table[3301] = 16'b0110100110011100; 
assign lut_table[3302] = 16'b0110100110011101; 
assign lut_table[3303] = 16'b0110100110011110; 
assign lut_table[3304] = 16'b0110100110011111; 
assign lut_table[3305] = 16'b0110100110101010; 
assign lut_table[3306] = 16'b0110100110101011; 
assign lut_table[3307] = 16'b0110100110101100; 
assign lut_table[3308] = 16'b0110100110101101; 
assign lut_table[3309] = 16'b0110100110101110; 
assign lut_table[3310] = 16'b0110100110101111; 
assign lut_table[3311] = 16'b0110100110111011; 
assign lut_table[3312] = 16'b0110100110111100; 
assign lut_table[3313] = 16'b0110100110111101; 
assign lut_table[3314] = 16'b0110100110111110; 
assign lut_table[3315] = 16'b0110100110111111; 
assign lut_table[3316] = 16'b0110100111001100; 
assign lut_table[3317] = 16'b0110100111001101; 
assign lut_table[3318] = 16'b0110100111001110; 
assign lut_table[3319] = 16'b0110100111001111; 
assign lut_table[3320] = 16'b0110100111011101; 
assign lut_table[3321] = 16'b0110100111011110; 
assign lut_table[3322] = 16'b0110100111011111; 
assign lut_table[3323] = 16'b0110100111101110; 
assign lut_table[3324] = 16'b0110100111101111; 
assign lut_table[3325] = 16'b0110100111111111; 
assign lut_table[3326] = 16'b0110101010101010; 
assign lut_table[3327] = 16'b0110101010101011; 
assign lut_table[3328] = 16'b0110101010101100; 
assign lut_table[3329] = 16'b0110101010101101; 
assign lut_table[3330] = 16'b0110101010101110; 
assign lut_table[3331] = 16'b0110101010101111; 
assign lut_table[3332] = 16'b0110101010111011; 
assign lut_table[3333] = 16'b0110101010111100; 
assign lut_table[3334] = 16'b0110101010111101; 
assign lut_table[3335] = 16'b0110101010111110; 
assign lut_table[3336] = 16'b0110101010111111; 
assign lut_table[3337] = 16'b0110101011001100; 
assign lut_table[3338] = 16'b0110101011001101; 
assign lut_table[3339] = 16'b0110101011001110; 
assign lut_table[3340] = 16'b0110101011001111; 
assign lut_table[3341] = 16'b0110101011011101; 
assign lut_table[3342] = 16'b0110101011011110; 
assign lut_table[3343] = 16'b0110101011011111; 
assign lut_table[3344] = 16'b0110101011101110; 
assign lut_table[3345] = 16'b0110101011101111; 
assign lut_table[3346] = 16'b0110101011111111; 
assign lut_table[3347] = 16'b0110101110111011; 
assign lut_table[3348] = 16'b0110101110111100; 
assign lut_table[3349] = 16'b0110101110111101; 
assign lut_table[3350] = 16'b0110101110111110; 
assign lut_table[3351] = 16'b0110101110111111; 
assign lut_table[3352] = 16'b0110101111001100; 
assign lut_table[3353] = 16'b0110101111001101; 
assign lut_table[3354] = 16'b0110101111001110; 
assign lut_table[3355] = 16'b0110101111001111; 
assign lut_table[3356] = 16'b0110101111011101; 
assign lut_table[3357] = 16'b0110101111011110; 
assign lut_table[3358] = 16'b0110101111011111; 
assign lut_table[3359] = 16'b0110101111101110; 
assign lut_table[3360] = 16'b0110101111101111; 
assign lut_table[3361] = 16'b0110101111111111; 
assign lut_table[3362] = 16'b0110110011001100; 
assign lut_table[3363] = 16'b0110110011001101; 
assign lut_table[3364] = 16'b0110110011001110; 
assign lut_table[3365] = 16'b0110110011001111; 
assign lut_table[3366] = 16'b0110110011011101; 
assign lut_table[3367] = 16'b0110110011011110; 
assign lut_table[3368] = 16'b0110110011011111; 
assign lut_table[3369] = 16'b0110110011101110; 
assign lut_table[3370] = 16'b0110110011101111; 
assign lut_table[3371] = 16'b0110110011111111; 
assign lut_table[3372] = 16'b0110110111011101; 
assign lut_table[3373] = 16'b0110110111011110; 
assign lut_table[3374] = 16'b0110110111011111; 
assign lut_table[3375] = 16'b0110110111101110; 
assign lut_table[3376] = 16'b0110110111101111; 
assign lut_table[3377] = 16'b0110110111111111; 
assign lut_table[3378] = 16'b0110111011101110; 
assign lut_table[3379] = 16'b0110111011101111; 
assign lut_table[3380] = 16'b0110111011111111; 
assign lut_table[3381] = 16'b0110111111111111; 
assign lut_table[3382] = 16'b0111011101110111; 
assign lut_table[3383] = 16'b0111011101111000; 
assign lut_table[3384] = 16'b0111011101111001; 
assign lut_table[3385] = 16'b0111011101111010; 
assign lut_table[3386] = 16'b0111011101111011; 
assign lut_table[3387] = 16'b0111011101111100; 
assign lut_table[3388] = 16'b0111011101111101; 
assign lut_table[3389] = 16'b0111011101111110; 
assign lut_table[3390] = 16'b0111011101111111; 
assign lut_table[3391] = 16'b0111011110001000; 
assign lut_table[3392] = 16'b0111011110001001; 
assign lut_table[3393] = 16'b0111011110001010; 
assign lut_table[3394] = 16'b0111011110001011; 
assign lut_table[3395] = 16'b0111011110001100; 
assign lut_table[3396] = 16'b0111011110001101; 
assign lut_table[3397] = 16'b0111011110001110; 
assign lut_table[3398] = 16'b0111011110001111; 
assign lut_table[3399] = 16'b0111011110011001; 
assign lut_table[3400] = 16'b0111011110011010; 
assign lut_table[3401] = 16'b0111011110011011; 
assign lut_table[3402] = 16'b0111011110011100; 
assign lut_table[3403] = 16'b0111011110011101; 
assign lut_table[3404] = 16'b0111011110011110; 
assign lut_table[3405] = 16'b0111011110011111; 
assign lut_table[3406] = 16'b0111011110101010; 
assign lut_table[3407] = 16'b0111011110101011; 
assign lut_table[3408] = 16'b0111011110101100; 
assign lut_table[3409] = 16'b0111011110101101; 
assign lut_table[3410] = 16'b0111011110101110; 
assign lut_table[3411] = 16'b0111011110101111; 
assign lut_table[3412] = 16'b0111011110111011; 
assign lut_table[3413] = 16'b0111011110111100; 
assign lut_table[3414] = 16'b0111011110111101; 
assign lut_table[3415] = 16'b0111011110111110; 
assign lut_table[3416] = 16'b0111011110111111; 
assign lut_table[3417] = 16'b0111011111001100; 
assign lut_table[3418] = 16'b0111011111001101; 
assign lut_table[3419] = 16'b0111011111001110; 
assign lut_table[3420] = 16'b0111011111001111; 
assign lut_table[3421] = 16'b0111011111011101; 
assign lut_table[3422] = 16'b0111011111011110; 
assign lut_table[3423] = 16'b0111011111011111; 
assign lut_table[3424] = 16'b0111011111101110; 
assign lut_table[3425] = 16'b0111011111101111; 
assign lut_table[3426] = 16'b0111011111111111; 
assign lut_table[3427] = 16'b0111100010001000; 
assign lut_table[3428] = 16'b0111100010001001; 
assign lut_table[3429] = 16'b0111100010001010; 
assign lut_table[3430] = 16'b0111100010001011; 
assign lut_table[3431] = 16'b0111100010001100; 
assign lut_table[3432] = 16'b0111100010001101; 
assign lut_table[3433] = 16'b0111100010001110; 
assign lut_table[3434] = 16'b0111100010001111; 
assign lut_table[3435] = 16'b0111100010011001; 
assign lut_table[3436] = 16'b0111100010011010; 
assign lut_table[3437] = 16'b0111100010011011; 
assign lut_table[3438] = 16'b0111100010011100; 
assign lut_table[3439] = 16'b0111100010011101; 
assign lut_table[3440] = 16'b0111100010011110; 
assign lut_table[3441] = 16'b0111100010011111; 
assign lut_table[3442] = 16'b0111100010101010; 
assign lut_table[3443] = 16'b0111100010101011; 
assign lut_table[3444] = 16'b0111100010101100; 
assign lut_table[3445] = 16'b0111100010101101; 
assign lut_table[3446] = 16'b0111100010101110; 
assign lut_table[3447] = 16'b0111100010101111; 
assign lut_table[3448] = 16'b0111100010111011; 
assign lut_table[3449] = 16'b0111100010111100; 
assign lut_table[3450] = 16'b0111100010111101; 
assign lut_table[3451] = 16'b0111100010111110; 
assign lut_table[3452] = 16'b0111100010111111; 
assign lut_table[3453] = 16'b0111100011001100; 
assign lut_table[3454] = 16'b0111100011001101; 
assign lut_table[3455] = 16'b0111100011001110; 
assign lut_table[3456] = 16'b0111100011001111; 
assign lut_table[3457] = 16'b0111100011011101; 
assign lut_table[3458] = 16'b0111100011011110; 
assign lut_table[3459] = 16'b0111100011011111; 
assign lut_table[3460] = 16'b0111100011101110; 
assign lut_table[3461] = 16'b0111100011101111; 
assign lut_table[3462] = 16'b0111100011111111; 
assign lut_table[3463] = 16'b0111100110011001; 
assign lut_table[3464] = 16'b0111100110011010; 
assign lut_table[3465] = 16'b0111100110011011; 
assign lut_table[3466] = 16'b0111100110011100; 
assign lut_table[3467] = 16'b0111100110011101; 
assign lut_table[3468] = 16'b0111100110011110; 
assign lut_table[3469] = 16'b0111100110011111; 
assign lut_table[3470] = 16'b0111100110101010; 
assign lut_table[3471] = 16'b0111100110101011; 
assign lut_table[3472] = 16'b0111100110101100; 
assign lut_table[3473] = 16'b0111100110101101; 
assign lut_table[3474] = 16'b0111100110101110; 
assign lut_table[3475] = 16'b0111100110101111; 
assign lut_table[3476] = 16'b0111100110111011; 
assign lut_table[3477] = 16'b0111100110111100; 
assign lut_table[3478] = 16'b0111100110111101; 
assign lut_table[3479] = 16'b0111100110111110; 
assign lut_table[3480] = 16'b0111100110111111; 
assign lut_table[3481] = 16'b0111100111001100; 
assign lut_table[3482] = 16'b0111100111001101; 
assign lut_table[3483] = 16'b0111100111001110; 
assign lut_table[3484] = 16'b0111100111001111; 
assign lut_table[3485] = 16'b0111100111011101; 
assign lut_table[3486] = 16'b0111100111011110; 
assign lut_table[3487] = 16'b0111100111011111; 
assign lut_table[3488] = 16'b0111100111101110; 
assign lut_table[3489] = 16'b0111100111101111; 
assign lut_table[3490] = 16'b0111100111111111; 
assign lut_table[3491] = 16'b0111101010101010; 
assign lut_table[3492] = 16'b0111101010101011; 
assign lut_table[3493] = 16'b0111101010101100; 
assign lut_table[3494] = 16'b0111101010101101; 
assign lut_table[3495] = 16'b0111101010101110; 
assign lut_table[3496] = 16'b0111101010101111; 
assign lut_table[3497] = 16'b0111101010111011; 
assign lut_table[3498] = 16'b0111101010111100; 
assign lut_table[3499] = 16'b0111101010111101; 
assign lut_table[3500] = 16'b0111101010111110; 
assign lut_table[3501] = 16'b0111101010111111; 
assign lut_table[3502] = 16'b0111101011001100; 
assign lut_table[3503] = 16'b0111101011001101; 
assign lut_table[3504] = 16'b0111101011001110; 
assign lut_table[3505] = 16'b0111101011001111; 
assign lut_table[3506] = 16'b0111101011011101; 
assign lut_table[3507] = 16'b0111101011011110; 
assign lut_table[3508] = 16'b0111101011011111; 
assign lut_table[3509] = 16'b0111101011101110; 
assign lut_table[3510] = 16'b0111101011101111; 
assign lut_table[3511] = 16'b0111101011111111; 
assign lut_table[3512] = 16'b0111101110111011; 
assign lut_table[3513] = 16'b0111101110111100; 
assign lut_table[3514] = 16'b0111101110111101; 
assign lut_table[3515] = 16'b0111101110111110; 
assign lut_table[3516] = 16'b0111101110111111; 
assign lut_table[3517] = 16'b0111101111001100; 
assign lut_table[3518] = 16'b0111101111001101; 
assign lut_table[3519] = 16'b0111101111001110; 
assign lut_table[3520] = 16'b0111101111001111; 
assign lut_table[3521] = 16'b0111101111011101; 
assign lut_table[3522] = 16'b0111101111011110; 
assign lut_table[3523] = 16'b0111101111011111; 
assign lut_table[3524] = 16'b0111101111101110; 
assign lut_table[3525] = 16'b0111101111101111; 
assign lut_table[3526] = 16'b0111101111111111; 
assign lut_table[3527] = 16'b0111110011001100; 
assign lut_table[3528] = 16'b0111110011001101; 
assign lut_table[3529] = 16'b0111110011001110; 
assign lut_table[3530] = 16'b0111110011001111; 
assign lut_table[3531] = 16'b0111110011011101; 
assign lut_table[3532] = 16'b0111110011011110; 
assign lut_table[3533] = 16'b0111110011011111; 
assign lut_table[3534] = 16'b0111110011101110; 
assign lut_table[3535] = 16'b0111110011101111; 
assign lut_table[3536] = 16'b0111110011111111; 
assign lut_table[3537] = 16'b0111110111011101; 
assign lut_table[3538] = 16'b0111110111011110; 
assign lut_table[3539] = 16'b0111110111011111; 
assign lut_table[3540] = 16'b0111110111101110; 
assign lut_table[3541] = 16'b0111110111101111; 
assign lut_table[3542] = 16'b0111110111111111; 
assign lut_table[3543] = 16'b0111111011101110; 
assign lut_table[3544] = 16'b0111111011101111; 
assign lut_table[3545] = 16'b0111111011111111; 
assign lut_table[3546] = 16'b0111111111111111; 
assign lut_table[3547] = 16'b1000100010001000; 
assign lut_table[3548] = 16'b1000100010001001; 
assign lut_table[3549] = 16'b1000100010001010; 
assign lut_table[3550] = 16'b1000100010001011; 
assign lut_table[3551] = 16'b1000100010001100; 
assign lut_table[3552] = 16'b1000100010001101; 
assign lut_table[3553] = 16'b1000100010001110; 
assign lut_table[3554] = 16'b1000100010001111; 
assign lut_table[3555] = 16'b1000100010011001; 
assign lut_table[3556] = 16'b1000100010011010; 
assign lut_table[3557] = 16'b1000100010011011; 
assign lut_table[3558] = 16'b1000100010011100; 
assign lut_table[3559] = 16'b1000100010011101; 
assign lut_table[3560] = 16'b1000100010011110; 
assign lut_table[3561] = 16'b1000100010011111; 
assign lut_table[3562] = 16'b1000100010101010; 
assign lut_table[3563] = 16'b1000100010101011; 
assign lut_table[3564] = 16'b1000100010101100; 
assign lut_table[3565] = 16'b1000100010101101; 
assign lut_table[3566] = 16'b1000100010101110; 
assign lut_table[3567] = 16'b1000100010101111; 
assign lut_table[3568] = 16'b1000100010111011; 
assign lut_table[3569] = 16'b1000100010111100; 
assign lut_table[3570] = 16'b1000100010111101; 
assign lut_table[3571] = 16'b1000100010111110; 
assign lut_table[3572] = 16'b1000100010111111; 
assign lut_table[3573] = 16'b1000100011001100; 
assign lut_table[3574] = 16'b1000100011001101; 
assign lut_table[3575] = 16'b1000100011001110; 
assign lut_table[3576] = 16'b1000100011001111; 
assign lut_table[3577] = 16'b1000100011011101; 
assign lut_table[3578] = 16'b1000100011011110; 
assign lut_table[3579] = 16'b1000100011011111; 
assign lut_table[3580] = 16'b1000100011101110; 
assign lut_table[3581] = 16'b1000100011101111; 
assign lut_table[3582] = 16'b1000100011111111; 
assign lut_table[3583] = 16'b1000100110011001; 
assign lut_table[3584] = 16'b1000100110011010; 
assign lut_table[3585] = 16'b1000100110011011; 
assign lut_table[3586] = 16'b1000100110011100; 
assign lut_table[3587] = 16'b1000100110011101; 
assign lut_table[3588] = 16'b1000100110011110; 
assign lut_table[3589] = 16'b1000100110011111; 
assign lut_table[3590] = 16'b1000100110101010; 
assign lut_table[3591] = 16'b1000100110101011; 
assign lut_table[3592] = 16'b1000100110101100; 
assign lut_table[3593] = 16'b1000100110101101; 
assign lut_table[3594] = 16'b1000100110101110; 
assign lut_table[3595] = 16'b1000100110101111; 
assign lut_table[3596] = 16'b1000100110111011; 
assign lut_table[3597] = 16'b1000100110111100; 
assign lut_table[3598] = 16'b1000100110111101; 
assign lut_table[3599] = 16'b1000100110111110; 
assign lut_table[3600] = 16'b1000100110111111; 
assign lut_table[3601] = 16'b1000100111001100; 
assign lut_table[3602] = 16'b1000100111001101; 
assign lut_table[3603] = 16'b1000100111001110; 
assign lut_table[3604] = 16'b1000100111001111; 
assign lut_table[3605] = 16'b1000100111011101; 
assign lut_table[3606] = 16'b1000100111011110; 
assign lut_table[3607] = 16'b1000100111011111; 
assign lut_table[3608] = 16'b1000100111101110; 
assign lut_table[3609] = 16'b1000100111101111; 
assign lut_table[3610] = 16'b1000100111111111; 
assign lut_table[3611] = 16'b1000101010101010; 
assign lut_table[3612] = 16'b1000101010101011; 
assign lut_table[3613] = 16'b1000101010101100; 
assign lut_table[3614] = 16'b1000101010101101; 
assign lut_table[3615] = 16'b1000101010101110; 
assign lut_table[3616] = 16'b1000101010101111; 
assign lut_table[3617] = 16'b1000101010111011; 
assign lut_table[3618] = 16'b1000101010111100; 
assign lut_table[3619] = 16'b1000101010111101; 
assign lut_table[3620] = 16'b1000101010111110; 
assign lut_table[3621] = 16'b1000101010111111; 
assign lut_table[3622] = 16'b1000101011001100; 
assign lut_table[3623] = 16'b1000101011001101; 
assign lut_table[3624] = 16'b1000101011001110; 
assign lut_table[3625] = 16'b1000101011001111; 
assign lut_table[3626] = 16'b1000101011011101; 
assign lut_table[3627] = 16'b1000101011011110; 
assign lut_table[3628] = 16'b1000101011011111; 
assign lut_table[3629] = 16'b1000101011101110; 
assign lut_table[3630] = 16'b1000101011101111; 
assign lut_table[3631] = 16'b1000101011111111; 
assign lut_table[3632] = 16'b1000101110111011; 
assign lut_table[3633] = 16'b1000101110111100; 
assign lut_table[3634] = 16'b1000101110111101; 
assign lut_table[3635] = 16'b1000101110111110; 
assign lut_table[3636] = 16'b1000101110111111; 
assign lut_table[3637] = 16'b1000101111001100; 
assign lut_table[3638] = 16'b1000101111001101; 
assign lut_table[3639] = 16'b1000101111001110; 
assign lut_table[3640] = 16'b1000101111001111; 
assign lut_table[3641] = 16'b1000101111011101; 
assign lut_table[3642] = 16'b1000101111011110; 
assign lut_table[3643] = 16'b1000101111011111; 
assign lut_table[3644] = 16'b1000101111101110; 
assign lut_table[3645] = 16'b1000101111101111; 
assign lut_table[3646] = 16'b1000101111111111; 
assign lut_table[3647] = 16'b1000110011001100; 
assign lut_table[3648] = 16'b1000110011001101; 
assign lut_table[3649] = 16'b1000110011001110; 
assign lut_table[3650] = 16'b1000110011001111; 
assign lut_table[3651] = 16'b1000110011011101; 
assign lut_table[3652] = 16'b1000110011011110; 
assign lut_table[3653] = 16'b1000110011011111; 
assign lut_table[3654] = 16'b1000110011101110; 
assign lut_table[3655] = 16'b1000110011101111; 
assign lut_table[3656] = 16'b1000110011111111; 
assign lut_table[3657] = 16'b1000110111011101; 
assign lut_table[3658] = 16'b1000110111011110; 
assign lut_table[3659] = 16'b1000110111011111; 
assign lut_table[3660] = 16'b1000110111101110; 
assign lut_table[3661] = 16'b1000110111101111; 
assign lut_table[3662] = 16'b1000110111111111; 
assign lut_table[3663] = 16'b1000111011101110; 
assign lut_table[3664] = 16'b1000111011101111; 
assign lut_table[3665] = 16'b1000111011111111; 
assign lut_table[3666] = 16'b1000111111111111; 
assign lut_table[3667] = 16'b1001100110011001; 
assign lut_table[3668] = 16'b1001100110011010; 
assign lut_table[3669] = 16'b1001100110011011; 
assign lut_table[3670] = 16'b1001100110011100; 
assign lut_table[3671] = 16'b1001100110011101; 
assign lut_table[3672] = 16'b1001100110011110; 
assign lut_table[3673] = 16'b1001100110011111; 
assign lut_table[3674] = 16'b1001100110101010; 
assign lut_table[3675] = 16'b1001100110101011; 
assign lut_table[3676] = 16'b1001100110101100; 
assign lut_table[3677] = 16'b1001100110101101; 
assign lut_table[3678] = 16'b1001100110101110; 
assign lut_table[3679] = 16'b1001100110101111; 
assign lut_table[3680] = 16'b1001100110111011; 
assign lut_table[3681] = 16'b1001100110111100; 
assign lut_table[3682] = 16'b1001100110111101; 
assign lut_table[3683] = 16'b1001100110111110; 
assign lut_table[3684] = 16'b1001100110111111; 
assign lut_table[3685] = 16'b1001100111001100; 
assign lut_table[3686] = 16'b1001100111001101; 
assign lut_table[3687] = 16'b1001100111001110; 
assign lut_table[3688] = 16'b1001100111001111; 
assign lut_table[3689] = 16'b1001100111011101; 
assign lut_table[3690] = 16'b1001100111011110; 
assign lut_table[3691] = 16'b1001100111011111; 
assign lut_table[3692] = 16'b1001100111101110; 
assign lut_table[3693] = 16'b1001100111101111; 
assign lut_table[3694] = 16'b1001100111111111; 
assign lut_table[3695] = 16'b1001101010101010; 
assign lut_table[3696] = 16'b1001101010101011; 
assign lut_table[3697] = 16'b1001101010101100; 
assign lut_table[3698] = 16'b1001101010101101; 
assign lut_table[3699] = 16'b1001101010101110; 
assign lut_table[3700] = 16'b1001101010101111; 
assign lut_table[3701] = 16'b1001101010111011; 
assign lut_table[3702] = 16'b1001101010111100; 
assign lut_table[3703] = 16'b1001101010111101; 
assign lut_table[3704] = 16'b1001101010111110; 
assign lut_table[3705] = 16'b1001101010111111; 
assign lut_table[3706] = 16'b1001101011001100; 
assign lut_table[3707] = 16'b1001101011001101; 
assign lut_table[3708] = 16'b1001101011001110; 
assign lut_table[3709] = 16'b1001101011001111; 
assign lut_table[3710] = 16'b1001101011011101; 
assign lut_table[3711] = 16'b1001101011011110; 
assign lut_table[3712] = 16'b1001101011011111; 
assign lut_table[3713] = 16'b1001101011101110; 
assign lut_table[3714] = 16'b1001101011101111; 
assign lut_table[3715] = 16'b1001101011111111; 
assign lut_table[3716] = 16'b1001101110111011; 
assign lut_table[3717] = 16'b1001101110111100; 
assign lut_table[3718] = 16'b1001101110111101; 
assign lut_table[3719] = 16'b1001101110111110; 
assign lut_table[3720] = 16'b1001101110111111; 
assign lut_table[3721] = 16'b1001101111001100; 
assign lut_table[3722] = 16'b1001101111001101; 
assign lut_table[3723] = 16'b1001101111001110; 
assign lut_table[3724] = 16'b1001101111001111; 
assign lut_table[3725] = 16'b1001101111011101; 
assign lut_table[3726] = 16'b1001101111011110; 
assign lut_table[3727] = 16'b1001101111011111; 
assign lut_table[3728] = 16'b1001101111101110; 
assign lut_table[3729] = 16'b1001101111101111; 
assign lut_table[3730] = 16'b1001101111111111; 
assign lut_table[3731] = 16'b1001110011001100; 
assign lut_table[3732] = 16'b1001110011001101; 
assign lut_table[3733] = 16'b1001110011001110; 
assign lut_table[3734] = 16'b1001110011001111; 
assign lut_table[3735] = 16'b1001110011011101; 
assign lut_table[3736] = 16'b1001110011011110; 
assign lut_table[3737] = 16'b1001110011011111; 
assign lut_table[3738] = 16'b1001110011101110; 
assign lut_table[3739] = 16'b1001110011101111; 
assign lut_table[3740] = 16'b1001110011111111; 
assign lut_table[3741] = 16'b1001110111011101; 
assign lut_table[3742] = 16'b1001110111011110; 
assign lut_table[3743] = 16'b1001110111011111; 
assign lut_table[3744] = 16'b1001110111101110; 
assign lut_table[3745] = 16'b1001110111101111; 
assign lut_table[3746] = 16'b1001110111111111; 
assign lut_table[3747] = 16'b1001111011101110; 
assign lut_table[3748] = 16'b1001111011101111; 
assign lut_table[3749] = 16'b1001111011111111; 
assign lut_table[3750] = 16'b1001111111111111; 
assign lut_table[3751] = 16'b1010101010101010; 
assign lut_table[3752] = 16'b1010101010101011; 
assign lut_table[3753] = 16'b1010101010101100; 
assign lut_table[3754] = 16'b1010101010101101; 
assign lut_table[3755] = 16'b1010101010101110; 
assign lut_table[3756] = 16'b1010101010101111; 
assign lut_table[3757] = 16'b1010101010111011; 
assign lut_table[3758] = 16'b1010101010111100; 
assign lut_table[3759] = 16'b1010101010111101; 
assign lut_table[3760] = 16'b1010101010111110; 
assign lut_table[3761] = 16'b1010101010111111; 
assign lut_table[3762] = 16'b1010101011001100; 
assign lut_table[3763] = 16'b1010101011001101; 
assign lut_table[3764] = 16'b1010101011001110; 
assign lut_table[3765] = 16'b1010101011001111; 
assign lut_table[3766] = 16'b1010101011011101; 
assign lut_table[3767] = 16'b1010101011011110; 
assign lut_table[3768] = 16'b1010101011011111; 
assign lut_table[3769] = 16'b1010101011101110; 
assign lut_table[3770] = 16'b1010101011101111; 
assign lut_table[3771] = 16'b1010101011111111; 
assign lut_table[3772] = 16'b1010101110111011; 
assign lut_table[3773] = 16'b1010101110111100; 
assign lut_table[3774] = 16'b1010101110111101; 
assign lut_table[3775] = 16'b1010101110111110; 
assign lut_table[3776] = 16'b1010101110111111; 
assign lut_table[3777] = 16'b1010101111001100; 
assign lut_table[3778] = 16'b1010101111001101; 
assign lut_table[3779] = 16'b1010101111001110; 
assign lut_table[3780] = 16'b1010101111001111; 
assign lut_table[3781] = 16'b1010101111011101; 
assign lut_table[3782] = 16'b1010101111011110; 
assign lut_table[3783] = 16'b1010101111011111; 
assign lut_table[3784] = 16'b1010101111101110; 
assign lut_table[3785] = 16'b1010101111101111; 
assign lut_table[3786] = 16'b1010101111111111; 
assign lut_table[3787] = 16'b1010110011001100; 
assign lut_table[3788] = 16'b1010110011001101; 
assign lut_table[3789] = 16'b1010110011001110; 
assign lut_table[3790] = 16'b1010110011001111; 
assign lut_table[3791] = 16'b1010110011011101; 
assign lut_table[3792] = 16'b1010110011011110; 
assign lut_table[3793] = 16'b1010110011011111; 
assign lut_table[3794] = 16'b1010110011101110; 
assign lut_table[3795] = 16'b1010110011101111; 
assign lut_table[3796] = 16'b1010110011111111; 
assign lut_table[3797] = 16'b1010110111011101; 
assign lut_table[3798] = 16'b1010110111011110; 
assign lut_table[3799] = 16'b1010110111011111; 
assign lut_table[3800] = 16'b1010110111101110; 
assign lut_table[3801] = 16'b1010110111101111; 
assign lut_table[3802] = 16'b1010110111111111; 
assign lut_table[3803] = 16'b1010111011101110; 
assign lut_table[3804] = 16'b1010111011101111; 
assign lut_table[3805] = 16'b1010111011111111; 
assign lut_table[3806] = 16'b1010111111111111; 
assign lut_table[3807] = 16'b1011101110111011; 
assign lut_table[3808] = 16'b1011101110111100; 
assign lut_table[3809] = 16'b1011101110111101; 
assign lut_table[3810] = 16'b1011101110111110; 
assign lut_table[3811] = 16'b1011101110111111; 
assign lut_table[3812] = 16'b1011101111001100; 
assign lut_table[3813] = 16'b1011101111001101; 
assign lut_table[3814] = 16'b1011101111001110; 
assign lut_table[3815] = 16'b1011101111001111; 
assign lut_table[3816] = 16'b1011101111011101; 
assign lut_table[3817] = 16'b1011101111011110; 
assign lut_table[3818] = 16'b1011101111011111; 
assign lut_table[3819] = 16'b1011101111101110; 
assign lut_table[3820] = 16'b1011101111101111; 
assign lut_table[3821] = 16'b1011101111111111; 
assign lut_table[3822] = 16'b1011110011001100; 
assign lut_table[3823] = 16'b1011110011001101; 
assign lut_table[3824] = 16'b1011110011001110; 
assign lut_table[3825] = 16'b1011110011001111; 
assign lut_table[3826] = 16'b1011110011011101; 
assign lut_table[3827] = 16'b1011110011011110; 
assign lut_table[3828] = 16'b1011110011011111; 
assign lut_table[3829] = 16'b1011110011101110; 
assign lut_table[3830] = 16'b1011110011101111; 
assign lut_table[3831] = 16'b1011110011111111; 
assign lut_table[3832] = 16'b1011110111011101; 
assign lut_table[3833] = 16'b1011110111011110; 
assign lut_table[3834] = 16'b1011110111011111; 
assign lut_table[3835] = 16'b1011110111101110; 
assign lut_table[3836] = 16'b1011110111101111; 
assign lut_table[3837] = 16'b1011110111111111; 
assign lut_table[3838] = 16'b1011111011101110; 
assign lut_table[3839] = 16'b1011111011101111; 
assign lut_table[3840] = 16'b1011111011111111; 
assign lut_table[3841] = 16'b1011111111111111; 
assign lut_table[3842] = 16'b1100110011001100; 
assign lut_table[3843] = 16'b1100110011001101; 
assign lut_table[3844] = 16'b1100110011001110; 
assign lut_table[3845] = 16'b1100110011001111; 
assign lut_table[3846] = 16'b1100110011011101; 
assign lut_table[3847] = 16'b1100110011011110; 
assign lut_table[3848] = 16'b1100110011011111; 
assign lut_table[3849] = 16'b1100110011101110; 
assign lut_table[3850] = 16'b1100110011101111; 
assign lut_table[3851] = 16'b1100110011111111; 
assign lut_table[3852] = 16'b1100110111011101; 
assign lut_table[3853] = 16'b1100110111011110; 
assign lut_table[3854] = 16'b1100110111011111; 
assign lut_table[3855] = 16'b1100110111101110; 
assign lut_table[3856] = 16'b1100110111101111; 
assign lut_table[3857] = 16'b1100110111111111; 
assign lut_table[3858] = 16'b1100111011101110; 
assign lut_table[3859] = 16'b1100111011101111; 
assign lut_table[3860] = 16'b1100111011111111; 
assign lut_table[3861] = 16'b1100111111111111; 
assign lut_table[3862] = 16'b1101110111011101; 
assign lut_table[3863] = 16'b1101110111011110; 
assign lut_table[3864] = 16'b1101110111011111; 
assign lut_table[3865] = 16'b1101110111101110; 
assign lut_table[3866] = 16'b1101110111101111; 
assign lut_table[3867] = 16'b1101110111111111; 
assign lut_table[3868] = 16'b1101111011101110; 
assign lut_table[3869] = 16'b1101111011101111; 
assign lut_table[3870] = 16'b1101111011111111; 
assign lut_table[3871] = 16'b1101111111111111; 
assign lut_table[3872] = 16'b1110111011101110; 
assign lut_table[3873] = 16'b1110111011101111; 
assign lut_table[3874] = 16'b1110111011111111; 
assign lut_table[3875] = 16'b1110111111111111; 
assign lut_table[3876] = 16'b1111111111111111; 

/*ENCODING*/
generate
  always@(msbs_i or msbs_j or msbs_k or msbs_w or encoding) begin
    for(int b = 0 ; b  < 8; b = b+1) begin
        code[b][0][11 : 0] = 12'b0;
        code[b][1][11 : 0] = 12'b0;
        code[b][2][11 : 0] = 12'b0;
        code[b][3][11 : 0] = 12'b0;
        if (encoding[b] == 1'b1)  begin
          for (int i = 0 ; i < 3877; i = i + 1) begin
            if (((lut_table[i][15 : 12]==msbs_i[b][0][3 : 0])&&(lut_table[i][11 : 8]==msbs_j[b][0][3 : 0]) && (lut_table[i][7 : 4] == msbs_k[b][0][3 : 0]) && (lut_table[i][3 : 0] == msbs_w[b][0][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_i[b][0][3 : 0])&&(lut_table[i][11 : 8]==msbs_j[b][0][3 : 0]) && (lut_table[i][7 : 4] == msbs_w[b][0][3 : 0]) && (lut_table[i][3 : 0] == msbs_k[b][0][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_i[b][0][3 : 0])&&(lut_table[i][11 : 8]==msbs_k[b][0][3 : 0]) && (lut_table[i][7 : 4] == msbs_j[b][0][3 : 0]) && (lut_table[i][3 : 0] == msbs_w[b][0][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_i[b][0][3 : 0])&&(lut_table[i][11 : 8]==msbs_k[b][0][3 : 0]) && (lut_table[i][7 : 4] == msbs_w[b][0][3 : 0]) && (lut_table[i][3 : 0] == msbs_j[b][0][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_i[b][0][3 : 0])&&(lut_table[i][11 : 8]==msbs_w[b][0][3 : 0]) && (lut_table[i][7 : 4] == msbs_j[b][0][3 : 0]) && (lut_table[i][3 : 0] == msbs_k[b][0][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_i[b][0][3 : 0])&&(lut_table[i][11 : 8]==msbs_w[b][0][3 : 0]) && (lut_table[i][7 : 4] == msbs_k[b][0][3 : 0]) && (lut_table[i][3 : 0] == msbs_j[b][0][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_j[b][0][3 : 0])&&(lut_table[i][11 : 8]==msbs_i[b][0][3 : 0]) && (lut_table[i][7 : 4] == msbs_k[b][0][3 : 0]) && (lut_table[i][3 : 0] == msbs_w[b][0][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_j[b][0][3 : 0])&&(lut_table[i][11 : 8]==msbs_i[b][0][3 : 0]) && (lut_table[i][7 : 4] == msbs_w[b][0][3 : 0]) && (lut_table[i][3 : 0] == msbs_k[b][0][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_j[b][0][3 : 0])&&(lut_table[i][11 : 8]==msbs_k[b][0][3 : 0]) && (lut_table[i][7 : 4] == msbs_i[b][0][3 : 0]) && (lut_table[i][3 : 0] == msbs_w[b][0][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_j[b][0][3 : 0])&&(lut_table[i][11 : 8]==msbs_k[b][0][3 : 0]) && (lut_table[i][7 : 4] == msbs_w[b][0][3 : 0]) && (lut_table[i][3 : 0] == msbs_i[b][0][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_j[b][0][3 : 0])&&(lut_table[i][11 : 8]==msbs_w[b][0][3 : 0]) && (lut_table[i][7 : 4] == msbs_i[b][0][3 : 0]) && (lut_table[i][3 : 0] == msbs_k[b][0][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_j[b][0][3 : 0])&&(lut_table[i][11 : 8]==msbs_w[b][0][3 : 0]) && (lut_table[i][7 : 4] == msbs_k[b][0][3 : 0]) && (lut_table[i][3 : 0] == msbs_i[b][0][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_k[b][0][3 : 0])&&(lut_table[i][11 : 8]==msbs_i[b][0][3 : 0]) && (lut_table[i][7 : 4] == msbs_j[b][0][3 : 0]) && (lut_table[i][3 : 0] == msbs_w[b][0][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_k[b][0][3 : 0])&&(lut_table[i][11 : 8]==msbs_i[b][0][3 : 0]) && (lut_table[i][7 : 4] == msbs_w[b][0][3 : 0]) && (lut_table[i][3 : 0] == msbs_j[b][0][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_k[b][0][3 : 0])&&(lut_table[i][11 : 8]==msbs_j[b][0][3 : 0]) && (lut_table[i][7 : 4] == msbs_i[b][0][3 : 0]) && (lut_table[i][3 : 0] == msbs_w[b][0][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_k[b][0][3 : 0])&&(lut_table[i][11 : 8]==msbs_j[b][0][3 : 0]) && (lut_table[i][7 : 4] == msbs_w[b][0][3 : 0]) && (lut_table[i][3 : 0] == msbs_i[b][0][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_k[b][0][3 : 0])&&(lut_table[i][11 : 8]==msbs_w[b][0][3 : 0]) && (lut_table[i][7 : 4] == msbs_i[b][0][3 : 0]) && (lut_table[i][3 : 0] == msbs_j[b][0][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_k[b][0][3 : 0])&&(lut_table[i][11 : 8]==msbs_w[b][0][3 : 0]) && (lut_table[i][7 : 4] == msbs_j[b][0][3 : 0]) && (lut_table[i][3 : 0] == msbs_i[b][0][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_w[b][0][3 : 0])&&(lut_table[i][11 : 8]==msbs_i[b][0][3 : 0]) && (lut_table[i][7 : 4] == msbs_j[b][0][3 : 0]) && (lut_table[i][3 : 0] == msbs_k[b][0][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_w[b][0][3 : 0])&&(lut_table[i][11 : 8]==msbs_i[b][0][3 : 0]) && (lut_table[i][7 : 4] == msbs_k[b][0][3 : 0]) && (lut_table[i][3 : 0] == msbs_j[b][0][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_w[b][0][3 : 0])&&(lut_table[i][11 : 8]==msbs_j[b][0][3 : 0]) && (lut_table[i][7 : 4] == msbs_i[b][0][3 : 0]) && (lut_table[i][3 : 0] == msbs_k[b][0][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_w[b][0][3 : 0])&&(lut_table[i][11 : 8]==msbs_j[b][0][3 : 0]) && (lut_table[i][7 : 4] == msbs_k[b][0][3 : 0]) && (lut_table[i][3 : 0] == msbs_i[b][0][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_w[b][0][3 : 0])&&(lut_table[i][11 : 8]==msbs_k[b][0][3 : 0]) && (lut_table[i][7 : 4] == msbs_i[b][0][3 : 0]) && (lut_table[i][3 : 0] == msbs_j[b][0][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_w[b][0][3 : 0])&&(lut_table[i][11 : 8]==msbs_k[b][0][3 : 0]) && (lut_table[i][7 : 4] == msbs_j[b][0][3 : 0]) && (lut_table[i][3 : 0] == msbs_i[b][0][3 : 0])) 
              ) begin
            code[b][0] = i[11 : 0];
            end 

            if (((lut_table[i][15 : 12]==msbs_i[b][1][3 : 0])&&(lut_table[i][11 : 8]==msbs_j[b][1][3 : 0]) && (lut_table[i][7 : 4] == msbs_k[b][1][3 : 0]) && (lut_table[i][3 : 0] == msbs_w[b][1][3 : 0])) ||
                  ((lut_table[i][15 : 12]==msbs_i[b][1][3 : 0])&&(lut_table[i][11 : 8]==msbs_j[b][1][3 : 0]) && (lut_table[i][7 : 4] == msbs_w[b][1][3 : 0]) && (lut_table[i][3 : 0] == msbs_k[b][1][3 : 0])) ||
                  ((lut_table[i][15 : 12]==msbs_i[b][1][3 : 0])&&(lut_table[i][11 : 8]==msbs_k[b][1][3 : 0]) && (lut_table[i][7 : 4] == msbs_j[b][1][3 : 0]) && (lut_table[i][3 : 0] == msbs_w[b][1][3 : 0])) ||
                  ((lut_table[i][15 : 12]==msbs_i[b][1][3 : 0])&&(lut_table[i][11 : 8]==msbs_k[b][1][3 : 0]) && (lut_table[i][7 : 4] == msbs_w[b][1][3 : 0]) && (lut_table[i][3 : 0] == msbs_j[b][1][3 : 0])) ||
                  ((lut_table[i][15 : 12]==msbs_i[b][1][3 : 0])&&(lut_table[i][11 : 8]==msbs_w[b][1][3 : 0]) && (lut_table[i][7 : 4] == msbs_j[b][1][3 : 0]) && (lut_table[i][3 : 0] == msbs_k[b][1][3 : 0])) ||
                  ((lut_table[i][15 : 12]==msbs_i[b][1][3 : 0])&&(lut_table[i][11 : 8]==msbs_w[b][1][3 : 0]) && (lut_table[i][7 : 4] == msbs_k[b][1][3 : 0]) && (lut_table[i][3 : 0] == msbs_j[b][1][3 : 0])) ||
                  ((lut_table[i][15 : 12]==msbs_j[b][1][3 : 0])&&(lut_table[i][11 : 8]==msbs_i[b][1][3 : 0]) && (lut_table[i][7 : 4] == msbs_k[b][1][3 : 0]) && (lut_table[i][3 : 0] == msbs_w[b][1][3 : 0])) ||
                  ((lut_table[i][15 : 12]==msbs_j[b][1][3 : 0])&&(lut_table[i][11 : 8]==msbs_i[b][1][3 : 0]) && (lut_table[i][7 : 4] == msbs_w[b][1][3 : 0]) && (lut_table[i][3 : 0] == msbs_k[b][1][3 : 0])) ||
                  ((lut_table[i][15 : 12]==msbs_j[b][1][3 : 0])&&(lut_table[i][11 : 8]==msbs_k[b][1][3 : 0]) && (lut_table[i][7 : 4] == msbs_i[b][1][3 : 0]) && (lut_table[i][3 : 0] == msbs_w[b][1][3 : 0])) ||
                  ((lut_table[i][15 : 12]==msbs_j[b][1][3 : 0])&&(lut_table[i][11 : 8]==msbs_k[b][1][3 : 0]) && (lut_table[i][7 : 4] == msbs_w[b][1][3 : 0]) && (lut_table[i][3 : 0] == msbs_i[b][1][3 : 0])) ||
                  ((lut_table[i][15 : 12]==msbs_j[b][1][3 : 0])&&(lut_table[i][11 : 8]==msbs_w[b][1][3 : 0]) && (lut_table[i][7 : 4] == msbs_i[b][1][3 : 0]) && (lut_table[i][3 : 0] == msbs_k[b][1][3 : 0])) ||
                  ((lut_table[i][15 : 12]==msbs_j[b][1][3 : 0])&&(lut_table[i][11 : 8]==msbs_w[b][1][3 : 0]) && (lut_table[i][7 : 4] == msbs_k[b][1][3 : 0]) && (lut_table[i][3 : 0] == msbs_i[b][1][3 : 0])) ||
                  ((lut_table[i][15 : 12]==msbs_k[b][1][3 : 0])&&(lut_table[i][11 : 8]==msbs_i[b][1][3 : 0]) && (lut_table[i][7 : 4] == msbs_j[b][1][3 : 0]) && (lut_table[i][3 : 0] == msbs_w[b][1][3 : 0])) ||
                  ((lut_table[i][15 : 12]==msbs_k[b][1][3 : 0])&&(lut_table[i][11 : 8]==msbs_i[b][1][3 : 0]) && (lut_table[i][7 : 4] == msbs_w[b][1][3 : 0]) && (lut_table[i][3 : 0] == msbs_j[b][1][3 : 0])) ||
                  ((lut_table[i][15 : 12]==msbs_k[b][1][3 : 0])&&(lut_table[i][11 : 8]==msbs_j[b][1][3 : 0]) && (lut_table[i][7 : 4] == msbs_i[b][1][3 : 0]) && (lut_table[i][3 : 0] == msbs_w[b][1][3 : 0])) ||
                  ((lut_table[i][15 : 12]==msbs_k[b][1][3 : 0])&&(lut_table[i][11 : 8]==msbs_j[b][1][3 : 0]) && (lut_table[i][7 : 4] == msbs_w[b][1][3 : 0]) && (lut_table[i][3 : 0] == msbs_i[b][1][3 : 0])) ||
                  ((lut_table[i][15 : 12]==msbs_k[b][1][3 : 0])&&(lut_table[i][11 : 8]==msbs_w[b][1][3 : 0]) && (lut_table[i][7 : 4] == msbs_i[b][1][3 : 0]) && (lut_table[i][3 : 0] == msbs_j[b][1][3 : 0])) ||
                  ((lut_table[i][15 : 12]==msbs_k[b][1][3 : 0])&&(lut_table[i][11 : 8]==msbs_w[b][1][3 : 0]) && (lut_table[i][7 : 4] == msbs_j[b][1][3 : 0]) && (lut_table[i][3 : 0] == msbs_i[b][1][3 : 0])) ||
                  ((lut_table[i][15 : 12]==msbs_w[b][1][3 : 0])&&(lut_table[i][11 : 8]==msbs_i[b][1][3 : 0]) && (lut_table[i][7 : 4] == msbs_j[b][1][3 : 0]) && (lut_table[i][3 : 0] == msbs_k[b][1][3 : 0])) ||
                  ((lut_table[i][15 : 12]==msbs_w[b][1][3 : 0])&&(lut_table[i][11 : 8]==msbs_i[b][1][3 : 0]) && (lut_table[i][7 : 4] == msbs_k[b][1][3 : 0]) && (lut_table[i][3 : 0] == msbs_j[b][1][3 : 0])) ||
                  ((lut_table[i][15 : 12]==msbs_w[b][1][3 : 0])&&(lut_table[i][11 : 8]==msbs_j[b][1][3 : 0]) && (lut_table[i][7 : 4] == msbs_i[b][1][3 : 0]) && (lut_table[i][3 : 0] == msbs_k[b][1][3 : 0])) ||
                  ((lut_table[i][15 : 12]==msbs_w[b][1][3 : 0])&&(lut_table[i][11 : 8]==msbs_j[b][1][3 : 0]) && (lut_table[i][7 : 4] == msbs_k[b][1][3 : 0]) && (lut_table[i][3 : 0] == msbs_i[b][1][3 : 0])) ||
                  ((lut_table[i][15 : 12]==msbs_w[b][1][3 : 0])&&(lut_table[i][11 : 8]==msbs_k[b][1][3 : 0]) && (lut_table[i][7 : 4] == msbs_i[b][1][3 : 0]) && (lut_table[i][3 : 0] == msbs_j[b][1][3 : 0])) ||
                  ((lut_table[i][15 : 12]==msbs_w[b][1][3 : 0])&&(lut_table[i][11 : 8]==msbs_k[b][1][3 : 0]) && (lut_table[i][7 : 4] == msbs_j[b][1][3 : 0]) && (lut_table[i][3 : 0] == msbs_i[b][1][3 : 0])) 
                ) begin
              code[b][1] = i[11 : 0];
              end 

            if (((lut_table[i][15 : 12]==msbs_i[b][2][3 : 0])&&(lut_table[i][11 : 8]==msbs_j[b][2][3 : 0]) && (lut_table[i][7 : 4] == msbs_k[b][2][3 : 0]) && (lut_table[i][3 : 0] == msbs_w[b][2][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_i[b][2][3 : 0])&&(lut_table[i][11 : 8]==msbs_j[b][2][3 : 0]) && (lut_table[i][7 : 4] == msbs_w[b][2][3 : 0]) && (lut_table[i][3 : 0] == msbs_k[b][2][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_i[b][2][3 : 0])&&(lut_table[i][11 : 8]==msbs_k[b][2][3 : 0]) && (lut_table[i][7 : 4] == msbs_j[b][2][3 : 0]) && (lut_table[i][3 : 0] == msbs_w[b][2][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_i[b][2][3 : 0])&&(lut_table[i][11 : 8]==msbs_k[b][2][3 : 0]) && (lut_table[i][7 : 4] == msbs_w[b][2][3 : 0]) && (lut_table[i][3 : 0] == msbs_j[b][2][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_i[b][2][3 : 0])&&(lut_table[i][11 : 8]==msbs_w[b][2][3 : 0]) && (lut_table[i][7 : 4] == msbs_j[b][2][3 : 0]) && (lut_table[i][3 : 0] == msbs_k[b][2][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_i[b][2][3 : 0])&&(lut_table[i][11 : 8]==msbs_w[b][2][3 : 0]) && (lut_table[i][7 : 4] == msbs_k[b][2][3 : 0]) && (lut_table[i][3 : 0] == msbs_j[b][2][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_j[b][2][3 : 0])&&(lut_table[i][11 : 8]==msbs_i[b][2][3 : 0]) && (lut_table[i][7 : 4] == msbs_k[b][2][3 : 0]) && (lut_table[i][3 : 0] == msbs_w[b][2][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_j[b][2][3 : 0])&&(lut_table[i][11 : 8]==msbs_i[b][2][3 : 0]) && (lut_table[i][7 : 4] == msbs_w[b][2][3 : 0]) && (lut_table[i][3 : 0] == msbs_k[b][2][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_j[b][2][3 : 0])&&(lut_table[i][11 : 8]==msbs_k[b][2][3 : 0]) && (lut_table[i][7 : 4] == msbs_i[b][2][3 : 0]) && (lut_table[i][3 : 0] == msbs_w[b][2][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_j[b][2][3 : 0])&&(lut_table[i][11 : 8]==msbs_k[b][2][3 : 0]) && (lut_table[i][7 : 4] == msbs_w[b][2][3 : 0]) && (lut_table[i][3 : 0] == msbs_i[b][2][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_j[b][2][3 : 0])&&(lut_table[i][11 : 8]==msbs_w[b][2][3 : 0]) && (lut_table[i][7 : 4] == msbs_i[b][2][3 : 0]) && (lut_table[i][3 : 0] == msbs_k[b][2][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_j[b][2][3 : 0])&&(lut_table[i][11 : 8]==msbs_w[b][2][3 : 0]) && (lut_table[i][7 : 4] == msbs_k[b][2][3 : 0]) && (lut_table[i][3 : 0] == msbs_i[b][2][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_k[b][2][3 : 0])&&(lut_table[i][11 : 8]==msbs_i[b][2][3 : 0]) && (lut_table[i][7 : 4] == msbs_j[b][2][3 : 0]) && (lut_table[i][3 : 0] == msbs_w[b][2][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_k[b][2][3 : 0])&&(lut_table[i][11 : 8]==msbs_i[b][2][3 : 0]) && (lut_table[i][7 : 4] == msbs_w[b][2][3 : 0]) && (lut_table[i][3 : 0] == msbs_j[b][2][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_k[b][2][3 : 0])&&(lut_table[i][11 : 8]==msbs_j[b][2][3 : 0]) && (lut_table[i][7 : 4] == msbs_i[b][2][3 : 0]) && (lut_table[i][3 : 0] == msbs_w[b][2][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_k[b][2][3 : 0])&&(lut_table[i][11 : 8]==msbs_j[b][2][3 : 0]) && (lut_table[i][7 : 4] == msbs_w[b][2][3 : 0]) && (lut_table[i][3 : 0] == msbs_i[b][2][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_k[b][2][3 : 0])&&(lut_table[i][11 : 8]==msbs_w[b][2][3 : 0]) && (lut_table[i][7 : 4] == msbs_i[b][2][3 : 0]) && (lut_table[i][3 : 0] == msbs_j[b][2][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_k[b][2][3 : 0])&&(lut_table[i][11 : 8]==msbs_w[b][2][3 : 0]) && (lut_table[i][7 : 4] == msbs_j[b][2][3 : 0]) && (lut_table[i][3 : 0] == msbs_i[b][2][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_w[b][2][3 : 0])&&(lut_table[i][11 : 8]==msbs_i[b][2][3 : 0]) && (lut_table[i][7 : 4] == msbs_j[b][2][3 : 0]) && (lut_table[i][3 : 0] == msbs_k[b][2][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_w[b][2][3 : 0])&&(lut_table[i][11 : 8]==msbs_i[b][2][3 : 0]) && (lut_table[i][7 : 4] == msbs_k[b][2][3 : 0]) && (lut_table[i][3 : 0] == msbs_j[b][2][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_w[b][2][3 : 0])&&(lut_table[i][11 : 8]==msbs_j[b][2][3 : 0]) && (lut_table[i][7 : 4] == msbs_i[b][2][3 : 0]) && (lut_table[i][3 : 0] == msbs_k[b][2][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_w[b][2][3 : 0])&&(lut_table[i][11 : 8]==msbs_j[b][2][3 : 0]) && (lut_table[i][7 : 4] == msbs_k[b][2][3 : 0]) && (lut_table[i][3 : 0] == msbs_i[b][2][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_w[b][2][3 : 0])&&(lut_table[i][11 : 8]==msbs_k[b][2][3 : 0]) && (lut_table[i][7 : 4] == msbs_i[b][2][3 : 0]) && (lut_table[i][3 : 0] == msbs_j[b][2][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_w[b][2][3 : 0])&&(lut_table[i][11 : 8]==msbs_k[b][2][3 : 0]) && (lut_table[i][7 : 4] == msbs_j[b][2][3 : 0]) && (lut_table[i][3 : 0] == msbs_i[b][2][3 : 0])) 
              ) begin
            code[b][2] = i[11 : 0];
            end 


          if (((lut_table[i][15 : 12]==msbs_i[b][3][3 : 0])&&(lut_table[i][11 : 8]==msbs_j[b][3][3 : 0]) && (lut_table[i][7 : 4] == msbs_k[b][3][3 : 0]) && (lut_table[i][3 : 0] == msbs_w[b][3][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_i[b][3][3 : 0])&&(lut_table[i][11 : 8]==msbs_j[b][3][3 : 0]) && (lut_table[i][7 : 4] == msbs_w[b][3][3 : 0]) && (lut_table[i][3 : 0] == msbs_k[b][3][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_i[b][3][3 : 0])&&(lut_table[i][11 : 8]==msbs_k[b][3][3 : 0]) && (lut_table[i][7 : 4] == msbs_j[b][3][3 : 0]) && (lut_table[i][3 : 0] == msbs_w[b][3][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_i[b][3][3 : 0])&&(lut_table[i][11 : 8]==msbs_k[b][3][3 : 0]) && (lut_table[i][7 : 4] == msbs_w[b][3][3 : 0]) && (lut_table[i][3 : 0] == msbs_j[b][3][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_i[b][3][3 : 0])&&(lut_table[i][11 : 8]==msbs_w[b][3][3 : 0]) && (lut_table[i][7 : 4] == msbs_j[b][3][3 : 0]) && (lut_table[i][3 : 0] == msbs_k[b][3][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_i[b][3][3 : 0])&&(lut_table[i][11 : 8]==msbs_w[b][3][3 : 0]) && (lut_table[i][7 : 4] == msbs_k[b][3][3 : 0]) && (lut_table[i][3 : 0] == msbs_j[b][3][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_j[b][3][3 : 0])&&(lut_table[i][11 : 8]==msbs_i[b][3][3 : 0]) && (lut_table[i][7 : 4] == msbs_k[b][3][3 : 0]) && (lut_table[i][3 : 0] == msbs_w[b][3][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_j[b][3][3 : 0])&&(lut_table[i][11 : 8]==msbs_i[b][3][3 : 0]) && (lut_table[i][7 : 4] == msbs_w[b][3][3 : 0]) && (lut_table[i][3 : 0] == msbs_k[b][3][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_j[b][3][3 : 0])&&(lut_table[i][11 : 8]==msbs_k[b][3][3 : 0]) && (lut_table[i][7 : 4] == msbs_i[b][3][3 : 0]) && (lut_table[i][3 : 0] == msbs_w[b][3][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_j[b][3][3 : 0])&&(lut_table[i][11 : 8]==msbs_k[b][3][3 : 0]) && (lut_table[i][7 : 4] == msbs_w[b][3][3 : 0]) && (lut_table[i][3 : 0] == msbs_i[b][3][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_j[b][3][3 : 0])&&(lut_table[i][11 : 8]==msbs_w[b][3][3 : 0]) && (lut_table[i][7 : 4] == msbs_i[b][3][3 : 0]) && (lut_table[i][3 : 0] == msbs_k[b][3][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_j[b][3][3 : 0])&&(lut_table[i][11 : 8]==msbs_w[b][3][3 : 0]) && (lut_table[i][7 : 4] == msbs_k[b][3][3 : 0]) && (lut_table[i][3 : 0] == msbs_i[b][3][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_k[b][3][3 : 0])&&(lut_table[i][11 : 8]==msbs_i[b][3][3 : 0]) && (lut_table[i][7 : 4] == msbs_j[b][3][3 : 0]) && (lut_table[i][3 : 0] == msbs_w[b][3][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_k[b][3][3 : 0])&&(lut_table[i][11 : 8]==msbs_i[b][3][3 : 0]) && (lut_table[i][7 : 4] == msbs_w[b][3][3 : 0]) && (lut_table[i][3 : 0] == msbs_j[b][3][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_k[b][3][3 : 0])&&(lut_table[i][11 : 8]==msbs_j[b][3][3 : 0]) && (lut_table[i][7 : 4] == msbs_i[b][3][3 : 0]) && (lut_table[i][3 : 0] == msbs_w[b][3][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_k[b][3][3 : 0])&&(lut_table[i][11 : 8]==msbs_j[b][3][3 : 0]) && (lut_table[i][7 : 4] == msbs_w[b][3][3 : 0]) && (lut_table[i][3 : 0] == msbs_i[b][3][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_k[b][3][3 : 0])&&(lut_table[i][11 : 8]==msbs_w[b][3][3 : 0]) && (lut_table[i][7 : 4] == msbs_i[b][3][3 : 0]) && (lut_table[i][3 : 0] == msbs_j[b][3][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_k[b][3][3 : 0])&&(lut_table[i][11 : 8]==msbs_w[b][3][3 : 0]) && (lut_table[i][7 : 4] == msbs_j[b][3][3 : 0]) && (lut_table[i][3 : 0] == msbs_i[b][3][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_w[b][3][3 : 0])&&(lut_table[i][11 : 8]==msbs_i[b][3][3 : 0]) && (lut_table[i][7 : 4] == msbs_j[b][3][3 : 0]) && (lut_table[i][3 : 0] == msbs_k[b][3][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_w[b][3][3 : 0])&&(lut_table[i][11 : 8]==msbs_i[b][3][3 : 0]) && (lut_table[i][7 : 4] == msbs_k[b][3][3 : 0]) && (lut_table[i][3 : 0] == msbs_j[b][3][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_w[b][3][3 : 0])&&(lut_table[i][11 : 8]==msbs_j[b][3][3 : 0]) && (lut_table[i][7 : 4] == msbs_i[b][3][3 : 0]) && (lut_table[i][3 : 0] == msbs_k[b][3][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_w[b][3][3 : 0])&&(lut_table[i][11 : 8]==msbs_j[b][3][3 : 0]) && (lut_table[i][7 : 4] == msbs_k[b][3][3 : 0]) && (lut_table[i][3 : 0] == msbs_i[b][3][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_w[b][3][3 : 0])&&(lut_table[i][11 : 8]==msbs_k[b][3][3 : 0]) && (lut_table[i][7 : 4] == msbs_i[b][3][3 : 0]) && (lut_table[i][3 : 0] == msbs_j[b][3][3 : 0])) ||
                ((lut_table[i][15 : 12]==msbs_w[b][3][3 : 0])&&(lut_table[i][11 : 8]==msbs_k[b][3][3 : 0]) && (lut_table[i][7 : 4] == msbs_j[b][3][3 : 0]) && (lut_table[i][3 : 0] == msbs_i[b][3][3 : 0])) 
              ) begin
            code[b][3] = i[11 : 0];
            end 
        end
      end 
    end
  end
endgenerate


/*DECODING*/
always @(to_decode or decoding) begin
  for(int b = 0; b  < 8 ; b = b +1) begin
    for (int p = 0 ; p  < 4 ; p = p+1)begin
      if (decoding[b] == 1'b1) begin
        decoded_msbs_i_reg[b][p][3 : 0] = lut_table[to_decode[b][p]][3 : 0];
        decoded_msbs_j_reg[b][p][3 : 0] = lut_table[to_decode[b][p]][7 : 4];
        decoded_msbs_k_reg[b][p][3 : 0] = lut_table[to_decode[b][p]][11 : 8];
        decoded_msbs_w_reg[b][p][3 : 0] = lut_table[to_decode[b][p]][15 : 12];
      end else begin
        decoded_msbs_i_reg[b][p] = 4'b0000;
        decoded_msbs_j_reg[b][p] = 4'b0000;
        decoded_msbs_k_reg[b][p] = 4'b0000;
        decoded_msbs_w_reg[b][p] = 4'b0000;
      end
    end
  end
end

assign code_o = code;
assign decoded_msbs_i = decoded_msbs_i_reg;
assign decoded_msbs_j = decoded_msbs_j_reg;
assign decoded_msbs_k = decoded_msbs_k_reg;
assign decoded_msbs_w = decoded_msbs_w_reg;


endmodule
