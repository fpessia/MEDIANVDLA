// ================================================================
// NVDLA Open Source Project
//
// Copyright(c) 2016 - 2017 NVIDIA Corporation. Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with
// this distribution for more information.
// ================================================================
// File Name: NV_BLKBOX_BUFFER.v
`timescale 10ps/1ps
module NV_BLKBOX_BUFFER (
  Y
 ,A
 );
output Y ;
input A ;
assign Y = A;
endmodule
