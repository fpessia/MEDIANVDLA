// ================================================================
// NVDLA Open Source Project
// 
// Copyright(c) 2016 - 2017 NVIDIA Corporation.  Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with 
// this distribution for more information.
// ================================================================

// File Name: NV_BLKBOX_SINK.v
`timescale 10ps/1ps
module  NV_BLKBOX_SINK (
	 A
	);

input	 A ;

endmodule

