// ================================================================
// NVDLA Open Source Project
//
// Copyright(c) 2016 - 2017 NVIDIA Corporation. Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with
// this distribution for more information.
// ================================================================
// File Name: NV_NVDLA_SDP_CORE_c.v
`timescale 10ps/1ps
module SDP_C_mgc_in_wire_wait_v1 (ld, vd, d, lz, vz, z);
  parameter integer rscid = 1;
  parameter integer width = 8;
  input ld;
  output vd;
  output [width-1:0] d;
  output lz;
  input vz;
  input [width-1:0] z;
  wire vd;
  wire [width-1:0] d;
  wire lz;
  assign d = z;
  assign lz = ld;
  assign vd = vz;
endmodule
//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/SDP_C_mgc_out_stdreg_wait_v1.v
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
// All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------
module SDP_C_mgc_out_stdreg_wait_v1 (ld, vd, d, lz, vz, z);
  parameter integer rscid = 1;
  parameter integer width = 8;
  input ld;
  output vd;
  input [width-1:0] d;
  output lz;
  input vz;
  output [width-1:0] z;
  wire vd;
  wire lz;
  wire [width-1:0] z;
  assign z = d;
  assign lz = ld;
  assign vd = vz;
endmodule
//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/SDP_C_mgc_in_wire_v1.v
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
// All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------
module SDP_C_mgc_in_wire_v1 (d, z);
  parameter integer rscid = 1;
  parameter integer width = 8;
  output [width-1:0] d;
  input [width-1:0] z;
  wire [width-1:0] d;
  assign d = z;
endmodule
//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/mgc_shift_r_beh_v4.v
module SDP_C_mgc_shift_r_v4(a,s,z);
   parameter width_a = 4;
   parameter signd_a = 1;
   parameter width_s = 2;
   parameter width_z = 8;
   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;
   generate
     if (signd_a)
     begin: SIGNED
       assign z = fshr_u(a,s,a[width_a-1]);
     end
     else
     begin: UNSIGNED
       assign z = fshr_u(a,s,1'b0);
     end
   endgenerate
//Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      int olen = width_z;
      int ilen = signd_a ? width_a : width_a+1;
      int len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u = result[olen-1:0];
      end
   endfunction // fshl_u
endmodule
//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/mgc_shift_br_beh_v4.v
module SDP_C_mgc_shift_br_v4(a,s,z);
   parameter width_a = 4;
   parameter signd_a = 1;
   parameter width_s = 2;
   parameter width_z = 8;
   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;
   generate
     if (signd_a)
     begin: SIGNED
       assign z = fshr_s(a,s,a[width_a-1]);
     end
     else
     begin: UNSIGNED
       assign z = fshr_s(a,s,1'b0);
     end
   endgenerate
//Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      int olen = width_z;
      int ilen = width_a+1;
      int len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 = result[olen-1:0];
      end
   endfunction // fshl_u
//Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      int olen = width_z;
      int ilen = signd_a ? width_a : width_a+1;
      int len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u = result[olen-1:0];
      end
   endfunction // fshr_u
//Shift right - signed shift argument
   function [width_z-1:0] fshr_s;
     input [width_a-1:0] arg1;
     input [width_s-1:0] arg2;
     input sbit;
     begin
       if ( arg2[width_s-1] == 1'b0 )
       begin
         fshr_s = fshr_u(arg1, arg2, sbit);
       end
       else
       begin
         fshr_s = fshl_u_1({arg1, 1'b0},~arg2, sbit);
       end
     end
   endfunction
endmodule
//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v4.v
module SDP_C_mgc_shift_l_v4(a,s,z);
   parameter width_a = 4;
   parameter signd_a = 1;
   parameter width_s = 2;
   parameter width_z = 8;
   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;
   generate
   if (signd_a)
   begin: SIGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSIGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate
//Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      int olen = width_z;
      int ilen = width_a+1;
      int len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 = result[olen-1:0];
      end
   endfunction // fshl_u
//Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u
endmodule
//------> ../td_ccore_solutions/leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_0/rtl.v
// ----------------------------------------------------------------------
// HLS HDL: Verilog Netlister
// HLS Version: 10.0/264918 Production Release
// HLS Date: Mon Aug 8 13:35:54 PDT 2016
//
// Generated by: ezhang@hk-sim-11-129
// Generated date: Thu May 4 10:35:41 2017
// ----------------------------------------------------------------------
//
// ------------------------------------------------------------------
// Design Unit: SDP_C_leading_sign_17_0
// ------------------------------------------------------------------
module SDP_C_leading_sign_17_0 (
  mantissa, rtn
);
  input [16:0] mantissa;
  output [4:0] rtn;
// Interconnect Declarations
  wire IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_6_2_sdt_2;
  wire IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_18_3_sdt_3;
  wire IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_26_2_sdt_2;
  wire IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_42_4_sdt_4;
  wire IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_6_2_sdt_1;
  wire IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_14_2_sdt_1;
  wire IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_26_2_sdt_1;
  wire IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_34_2_sdt_1;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_7;
  wire[0:0] IntLeadZero_17U_leading_sign_17_0_rtn_and_63_nl;
  wire[0:0] IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_nor_nl;
  wire[0:0] IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_nor_10_nl;
  wire[0:0] IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_or_nl;
// Interconnect Declarations for Component Instantiations
  assign IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_6_2_sdt_2 = ~((mantissa[14:13]!=2'b00));
  assign IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_6_2_sdt_1 = ~((mantissa[16:15]!=2'b00));
  assign IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_14_2_sdt_1 = ~((mantissa[12:11]!=2'b00));
  assign c_h_1_2 = IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_6_2_sdt_1 & IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_6_2_sdt_2;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_18_3_sdt_3 = (mantissa[10:9]==2'b00)
      & IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_14_2_sdt_1;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_26_2_sdt_2 = ~((mantissa[6:5]!=2'b00));
  assign IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_26_2_sdt_1 = ~((mantissa[8:7]!=2'b00));
  assign IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_34_2_sdt_1 = ~((mantissa[4:3]!=2'b00));
  assign c_h_1_5 = IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_26_2_sdt_1 & IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_18_3_sdt_3;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_42_4_sdt_4 = (mantissa[2:1]==2'b00)
      & IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_34_2_sdt_1 & c_h_1_5;
  assign c_h_1_7 = c_h_1_6 & IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_42_4_sdt_4;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_and_63_nl = c_h_1_6 & (~ IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_42_4_sdt_4);
  assign IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_nor_nl
      = ~((~(c_h_1_2 & (c_h_1_5 | (~ IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_18_3_sdt_3))))
      | c_h_1_7);
  assign IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_nor_10_nl
      = ~((~(IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_6_2_sdt_1 & (IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_14_2_sdt_1
      | (~ IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_6_2_sdt_2)) & (~((~(IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_26_2_sdt_1
      & (IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_34_2_sdt_1 | (~ IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_26_2_sdt_2))))
      & c_h_1_6)))) | c_h_1_7);
  assign IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_or_nl
      = (~((~((~((mantissa[16]) | (~((mantissa[15:14]!=2'b01))))) & (~(((mantissa[12])
      | (~((mantissa[11:10]!=2'b01)))) & c_h_1_2)) & (~((~((~((mantissa[8]) | (~((mantissa[7:6]!=2'b01)))))
      & (~(((mantissa[4]) | (~((mantissa[3:2]!=2'b01)))) & c_h_1_5)))) & c_h_1_6))))
      | c_h_1_7)) | ((~ (mantissa[0])) & c_h_1_7);
  assign rtn = {c_h_1_7 , (IntLeadZero_17U_leading_sign_17_0_rtn_and_63_nl) , (IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_nor_nl)
      , (IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_nor_10_nl)
      , (IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_or_nl)};
endmodule
//------> ./rtl.v
// ----------------------------------------------------------------------
// HLS HDL: Verilog Netlister
// HLS Version: 10.0/264918 Production Release
// HLS Date: Mon Aug 8 13:35:54 PDT 2016
//
// Generated by: ezhang@hk-sim-10-055
// Generated date: Thu Jul 6 14:02:16 2017
// ----------------------------------------------------------------------
//
// ------------------------------------------------------------------
// Design Unit: SDP_C_chn_out_rsci_unreg
// ------------------------------------------------------------------
module SDP_C_chn_out_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: SDP_C_chn_in_rsci_unreg
// ------------------------------------------------------------------
module SDP_C_chn_in_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;
// Interconnect Declarations for Component Instantiations
  assign outsig = in_0;
endmodule
// ------------------------------------------------------------------
// Design Unit: NV_NVDLA_SDP_CORE_c_core_core_fsm
// FSM Module
// ------------------------------------------------------------------
module NV_NVDLA_SDP_CORE_c_core_core_fsm (
  nvdla_core_clk, nvdla_core_rstn, core_wen, fsm_output
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;
// FSM State Type Declaration for NV_NVDLA_SDP_CORE_c_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;
  reg [0:0] state_var;
  reg [0:0] state_var_NS;
// Interconnect Declarations for Component Instantiations
  always @(*)
  begin : NV_NVDLA_SDP_CORE_c_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
// core_rlp_C_0
      default : begin
        fsm_output = 2'b1;
        state_var_NS = main_C_0;
      end
    endcase
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: NV_NVDLA_SDP_CORE_c_core_staller
// ------------------------------------------------------------------
module NV_NVDLA_SDP_CORE_c_core_staller (
  nvdla_core_clk, nvdla_core_rstn, core_wen, chn_in_rsci_wen_comp, core_wten, chn_out_rsci_wen_comp
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output core_wen;
  input chn_in_rsci_wen_comp;
  output core_wten;
  reg core_wten;
  input chn_out_rsci_wen_comp;
// Interconnect Declarations for Component Instantiations
  assign core_wen = chn_in_rsci_wen_comp & chn_out_rsci_wen_comp;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      core_wten <= 1'b0;
    end
    else begin
      core_wten <= ~ core_wen;
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: NV_NVDLA_SDP_CORE_c_core_chn_out_rsci_chn_out_wait_dp
// ------------------------------------------------------------------
module NV_NVDLA_SDP_CORE_c_core_chn_out_rsci_chn_out_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_out_rsci_oswt, chn_out_rsci_bawt, chn_out_rsci_wen_comp,
      chn_out_rsci_biwt, chn_out_rsci_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_out_rsci_oswt;
  output chn_out_rsci_bawt;
  output chn_out_rsci_wen_comp;
  input chn_out_rsci_biwt;
  input chn_out_rsci_bdwt;
// Interconnect Declarations
  reg chn_out_rsci_bcwt;
// Interconnect Declarations for Component Instantiations
  assign chn_out_rsci_bawt = chn_out_rsci_biwt | chn_out_rsci_bcwt;
  assign chn_out_rsci_wen_comp = (~ chn_out_rsci_oswt) | chn_out_rsci_bawt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_out_rsci_bcwt <= 1'b0;
    end
    else begin
      chn_out_rsci_bcwt <= ~((~(chn_out_rsci_bcwt | chn_out_rsci_biwt)) | chn_out_rsci_bdwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: NV_NVDLA_SDP_CORE_c_core_chn_out_rsci_chn_out_wait_ctrl
// ------------------------------------------------------------------
module NV_NVDLA_SDP_CORE_c_core_chn_out_rsci_chn_out_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_out_rsci_oswt, core_wen, core_wten, chn_out_rsci_iswt0,
      chn_out_rsci_ld_core_psct, chn_out_rsci_biwt, chn_out_rsci_bdwt, chn_out_rsci_ld_core_sct,
      chn_out_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_out_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_out_rsci_iswt0;
  input chn_out_rsci_ld_core_psct;
  output chn_out_rsci_biwt;
  output chn_out_rsci_bdwt;
  output chn_out_rsci_ld_core_sct;
  input chn_out_rsci_vd;
// Interconnect Declarations
  wire chn_out_rsci_ogwt;
  wire chn_out_rsci_pdswt0;
  reg chn_out_rsci_icwt;
// Interconnect Declarations for Component Instantiations
  assign chn_out_rsci_pdswt0 = (~ core_wten) & chn_out_rsci_iswt0;
  assign chn_out_rsci_biwt = chn_out_rsci_ogwt & chn_out_rsci_vd;
  assign chn_out_rsci_ogwt = chn_out_rsci_pdswt0 | chn_out_rsci_icwt;
  assign chn_out_rsci_bdwt = chn_out_rsci_oswt & core_wen;
  assign chn_out_rsci_ld_core_sct = chn_out_rsci_ld_core_psct & chn_out_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_out_rsci_icwt <= 1'b0;
    end
    else begin
      chn_out_rsci_icwt <= ~((~(chn_out_rsci_icwt | chn_out_rsci_pdswt0)) | chn_out_rsci_biwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: NV_NVDLA_SDP_CORE_c_core_chn_in_rsci_chn_in_wait_dp
// ------------------------------------------------------------------
module NV_NVDLA_SDP_CORE_c_core_chn_in_rsci_chn_in_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_in_rsci_oswt, chn_in_rsci_bawt, chn_in_rsci_wen_comp,
      chn_in_rsci_d_mxwt, chn_in_rsci_biwt, chn_in_rsci_bdwt, chn_in_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_in_rsci_oswt;
  output chn_in_rsci_bawt;
  output chn_in_rsci_wen_comp;
  output [511:0] chn_in_rsci_d_mxwt;
  input chn_in_rsci_biwt;
  input chn_in_rsci_bdwt;
  input [511:0] chn_in_rsci_d;
// Interconnect Declarations
  reg chn_in_rsci_bcwt;
  reg [511:0] chn_in_rsci_d_bfwt;
// Interconnect Declarations for Component Instantiations
  assign chn_in_rsci_bawt = chn_in_rsci_biwt | chn_in_rsci_bcwt;
  assign chn_in_rsci_wen_comp = (~ chn_in_rsci_oswt) | chn_in_rsci_bawt;
  assign chn_in_rsci_d_mxwt = MUX_v_512_2_2(chn_in_rsci_d, chn_in_rsci_d_bfwt, chn_in_rsci_bcwt);
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_in_rsci_bcwt <= 1'b0;
      chn_in_rsci_d_bfwt <= 512'b0;
    end
    else begin
      chn_in_rsci_bcwt <= ~((~(chn_in_rsci_bcwt | chn_in_rsci_biwt)) | chn_in_rsci_bdwt);
      chn_in_rsci_d_bfwt <= chn_in_rsci_d_mxwt;
    end
  end
  function [511:0] MUX_v_512_2_2;
    input [511:0] input_0;
    input [511:0] input_1;
    input [0:0] sel;
    reg [511:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_512_2_2 = result;
  end
  endfunction
endmodule
// ------------------------------------------------------------------
// Design Unit: NV_NVDLA_SDP_CORE_c_core_chn_in_rsci_chn_in_wait_ctrl
// ------------------------------------------------------------------
module NV_NVDLA_SDP_CORE_c_core_chn_in_rsci_chn_in_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_in_rsci_oswt, core_wen, chn_in_rsci_iswt0,
      chn_in_rsci_ld_core_psct, core_wten, chn_in_rsci_biwt, chn_in_rsci_bdwt, chn_in_rsci_ld_core_sct,
      chn_in_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_in_rsci_oswt;
  input core_wen;
  input chn_in_rsci_iswt0;
  input chn_in_rsci_ld_core_psct;
  input core_wten;
  output chn_in_rsci_biwt;
  output chn_in_rsci_bdwt;
  output chn_in_rsci_ld_core_sct;
  input chn_in_rsci_vd;
// Interconnect Declarations
  wire chn_in_rsci_ogwt;
  wire chn_in_rsci_pdswt0;
  reg chn_in_rsci_icwt;
// Interconnect Declarations for Component Instantiations
  assign chn_in_rsci_pdswt0 = (~ core_wten) & chn_in_rsci_iswt0;
  assign chn_in_rsci_biwt = chn_in_rsci_ogwt & chn_in_rsci_vd;
  assign chn_in_rsci_ogwt = chn_in_rsci_pdswt0 | chn_in_rsci_icwt;
  assign chn_in_rsci_bdwt = chn_in_rsci_oswt & core_wen;
  assign chn_in_rsci_ld_core_sct = chn_in_rsci_ld_core_psct & chn_in_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_in_rsci_icwt <= 1'b0;
    end
    else begin
      chn_in_rsci_icwt <= ~((~(chn_in_rsci_icwt | chn_in_rsci_pdswt0)) | chn_in_rsci_biwt);
    end
  end
endmodule
// ------------------------------------------------------------------
// Design Unit: NV_NVDLA_SDP_CORE_c_core_chn_out_rsci
// ------------------------------------------------------------------
module NV_NVDLA_SDP_CORE_c_core_chn_out_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_out_rsc_z, chn_out_rsc_vz, chn_out_rsc_lz,
      chn_out_rsci_oswt, core_wen, core_wten, chn_out_rsci_iswt0, chn_out_rsci_bawt,
      chn_out_rsci_wen_comp, chn_out_rsci_ld_core_psct, chn_out_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output [271:0] chn_out_rsc_z;
  input chn_out_rsc_vz;
  output chn_out_rsc_lz;
  input chn_out_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_out_rsci_iswt0;
  output chn_out_rsci_bawt;
  output chn_out_rsci_wen_comp;
  input chn_out_rsci_ld_core_psct;
  input [271:0] chn_out_rsci_d;
// Interconnect Declarations
  wire chn_out_rsci_biwt;
  wire chn_out_rsci_bdwt;
  wire chn_out_rsci_ld_core_sct;
  wire chn_out_rsci_vd;
// Interconnect Declarations for Component Instantiations
  SDP_C_mgc_out_stdreg_wait_v1 #(.rscid(32'sd8),
  .width(32'sd272)) chn_out_rsci (
      .ld(chn_out_rsci_ld_core_sct),
      .vd(chn_out_rsci_vd),
      .d(chn_out_rsci_d),
      .lz(chn_out_rsc_lz),
      .vz(chn_out_rsc_vz),
      .z(chn_out_rsc_z)
    );
  NV_NVDLA_SDP_CORE_c_core_chn_out_rsci_chn_out_wait_ctrl NV_NVDLA_SDP_CORE_c_core_chn_out_rsci_chn_out_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_out_rsci_oswt(chn_out_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_out_rsci_iswt0(chn_out_rsci_iswt0),
      .chn_out_rsci_ld_core_psct(chn_out_rsci_ld_core_psct),
      .chn_out_rsci_biwt(chn_out_rsci_biwt),
      .chn_out_rsci_bdwt(chn_out_rsci_bdwt),
      .chn_out_rsci_ld_core_sct(chn_out_rsci_ld_core_sct),
      .chn_out_rsci_vd(chn_out_rsci_vd)
    );
  NV_NVDLA_SDP_CORE_c_core_chn_out_rsci_chn_out_wait_dp NV_NVDLA_SDP_CORE_c_core_chn_out_rsci_chn_out_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_out_rsci_oswt(chn_out_rsci_oswt),
      .chn_out_rsci_bawt(chn_out_rsci_bawt),
      .chn_out_rsci_wen_comp(chn_out_rsci_wen_comp),
      .chn_out_rsci_biwt(chn_out_rsci_biwt),
      .chn_out_rsci_bdwt(chn_out_rsci_bdwt)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: NV_NVDLA_SDP_CORE_c_core_chn_in_rsci
// ------------------------------------------------------------------
module NV_NVDLA_SDP_CORE_c_core_chn_in_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_in_rsc_z, chn_in_rsc_vz, chn_in_rsc_lz, chn_in_rsci_oswt,
      core_wen, chn_in_rsci_iswt0, chn_in_rsci_bawt, chn_in_rsci_wen_comp, chn_in_rsci_ld_core_psct,
      chn_in_rsci_d_mxwt, core_wten
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [511:0] chn_in_rsc_z;
  input chn_in_rsc_vz;
  output chn_in_rsc_lz;
  input chn_in_rsci_oswt;
  input core_wen;
  input chn_in_rsci_iswt0;
  output chn_in_rsci_bawt;
  output chn_in_rsci_wen_comp;
  input chn_in_rsci_ld_core_psct;
  output [511:0] chn_in_rsci_d_mxwt;
  input core_wten;
// Interconnect Declarations
  wire chn_in_rsci_biwt;
  wire chn_in_rsci_bdwt;
  wire chn_in_rsci_ld_core_sct;
  wire chn_in_rsci_vd;
  wire [511:0] chn_in_rsci_d;
// Interconnect Declarations for Component Instantiations
  SDP_C_mgc_in_wire_wait_v1 #(.rscid(32'sd1),
  .width(32'sd512)) chn_in_rsci (
      .ld(chn_in_rsci_ld_core_sct),
      .vd(chn_in_rsci_vd),
      .d(chn_in_rsci_d),
      .lz(chn_in_rsc_lz),
      .vz(chn_in_rsc_vz),
      .z(chn_in_rsc_z)
    );
  NV_NVDLA_SDP_CORE_c_core_chn_in_rsci_chn_in_wait_ctrl NV_NVDLA_SDP_CORE_c_core_chn_in_rsci_chn_in_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_in_rsci_oswt(chn_in_rsci_oswt),
      .core_wen(core_wen),
      .chn_in_rsci_iswt0(chn_in_rsci_iswt0),
      .chn_in_rsci_ld_core_psct(chn_in_rsci_ld_core_psct),
      .core_wten(core_wten),
      .chn_in_rsci_biwt(chn_in_rsci_biwt),
      .chn_in_rsci_bdwt(chn_in_rsci_bdwt),
      .chn_in_rsci_ld_core_sct(chn_in_rsci_ld_core_sct),
      .chn_in_rsci_vd(chn_in_rsci_vd)
    );
  NV_NVDLA_SDP_CORE_c_core_chn_in_rsci_chn_in_wait_dp NV_NVDLA_SDP_CORE_c_core_chn_in_rsci_chn_in_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_in_rsci_oswt(chn_in_rsci_oswt),
      .chn_in_rsci_bawt(chn_in_rsci_bawt),
      .chn_in_rsci_wen_comp(chn_in_rsci_wen_comp),
      .chn_in_rsci_d_mxwt(chn_in_rsci_d_mxwt),
      .chn_in_rsci_biwt(chn_in_rsci_biwt),
      .chn_in_rsci_bdwt(chn_in_rsci_bdwt),
      .chn_in_rsci_d(chn_in_rsci_d)
    );
endmodule
// ------------------------------------------------------------------
// Design Unit: NV_NVDLA_SDP_CORE_c_core
// ------------------------------------------------------------------
module NV_NVDLA_SDP_CORE_c_core (
  nvdla_core_clk, nvdla_core_rstn, chn_in_rsc_z, chn_in_rsc_vz, chn_in_rsc_lz, cfg_offset_rsc_z,
      cfg_scale_rsc_z, cfg_truncate_rsc_z, cfg_proc_precision_rsc_z, cfg_out_precision_rsc_z,
      cfg_mode_eql_rsc_z, chn_out_rsc_z, chn_out_rsc_vz, chn_out_rsc_lz, chn_in_rsci_oswt,
      chn_in_rsci_oswt_unreg, chn_out_rsci_oswt, chn_out_rsci_oswt_unreg
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [511:0] chn_in_rsc_z;
  input chn_in_rsc_vz;
  output chn_in_rsc_lz;
  input [31:0] cfg_offset_rsc_z;
  input [15:0] cfg_scale_rsc_z;
  input [5:0] cfg_truncate_rsc_z;
  input [1:0] cfg_proc_precision_rsc_z;
  input [1:0] cfg_out_precision_rsc_z;
  input cfg_mode_eql_rsc_z;
  output [271:0] chn_out_rsc_z;
  input chn_out_rsc_vz;
  output chn_out_rsc_lz;
  input chn_in_rsci_oswt;
  output chn_in_rsci_oswt_unreg;
  input chn_out_rsci_oswt;
  output chn_out_rsci_oswt_unreg;
// Interconnect Declarations
  wire core_wen;
  reg chn_in_rsci_iswt0;
  wire chn_in_rsci_bawt;
  wire chn_in_rsci_wen_comp;
  reg chn_in_rsci_ld_core_psct;
  wire [511:0] chn_in_rsci_d_mxwt;
  wire core_wten;
  wire [31:0] cfg_offset_rsci_d;
  wire [15:0] cfg_scale_rsci_d;
  wire [5:0] cfg_truncate_rsci_d;
  wire [1:0] cfg_proc_precision_rsci_d;
  wire [1:0] cfg_out_precision_rsci_d;
  wire cfg_mode_eql_rsci_d;
  reg chn_out_rsci_iswt0;
  wire chn_out_rsci_bawt;
  wire chn_out_rsci_wen_comp;
  reg chn_out_rsci_d_271;
  reg chn_out_rsci_d_270;
  reg chn_out_rsci_d_269;
  reg chn_out_rsci_d_268;
  reg chn_out_rsci_d_267;
  reg chn_out_rsci_d_266;
  reg chn_out_rsci_d_265;
  reg chn_out_rsci_d_264;
  reg chn_out_rsci_d_263;
  reg chn_out_rsci_d_262;
  reg chn_out_rsci_d_261;
  reg chn_out_rsci_d_260;
  reg chn_out_rsci_d_259;
  reg chn_out_rsci_d_258;
  reg chn_out_rsci_d_257;
  reg chn_out_rsci_d_256;
  reg chn_out_rsci_d_255;
  reg [8:0] chn_out_rsci_d_249_241;
  reg chn_out_rsci_d_240;
  reg chn_out_rsci_d_239;
  reg [8:0] chn_out_rsci_d_233_225;
  reg chn_out_rsci_d_224;
  reg chn_out_rsci_d_223;
  reg [8:0] chn_out_rsci_d_217_209;
  reg chn_out_rsci_d_208;
  reg chn_out_rsci_d_207;
  reg [8:0] chn_out_rsci_d_201_193;
  reg chn_out_rsci_d_192;
  reg chn_out_rsci_d_191;
  reg [8:0] chn_out_rsci_d_185_177;
  reg chn_out_rsci_d_176;
  reg chn_out_rsci_d_175;
  reg [8:0] chn_out_rsci_d_169_161;
  reg chn_out_rsci_d_160;
  reg chn_out_rsci_d_159;
  reg [8:0] chn_out_rsci_d_153_145;
  reg chn_out_rsci_d_144;
  reg chn_out_rsci_d_143;
  reg [8:0] chn_out_rsci_d_137_129;
  reg chn_out_rsci_d_128;
  reg chn_out_rsci_d_127;
  reg [8:0] chn_out_rsci_d_121_113;
  reg chn_out_rsci_d_112;
  reg chn_out_rsci_d_111;
  reg [8:0] chn_out_rsci_d_105_97;
  reg chn_out_rsci_d_96;
  reg chn_out_rsci_d_95;
  reg [8:0] chn_out_rsci_d_89_81;
  reg chn_out_rsci_d_80;
  reg chn_out_rsci_d_79;
  reg [8:0] chn_out_rsci_d_73_65;
  reg chn_out_rsci_d_64;
  reg chn_out_rsci_d_63;
  reg [8:0] chn_out_rsci_d_57_49;
  reg chn_out_rsci_d_48;
  reg chn_out_rsci_d_47;
  reg [8:0] chn_out_rsci_d_41_33;
  reg chn_out_rsci_d_32;
  reg chn_out_rsci_d_31;
  reg [8:0] chn_out_rsci_d_25_17;
  reg chn_out_rsci_d_16;
  reg chn_out_rsci_d_15;
  reg [8:0] chn_out_rsci_d_9_1;
  reg chn_out_rsci_d_0;
  reg chn_out_rsci_d_254;
  reg [3:0] chn_out_rsci_d_253_250;
  reg chn_out_rsci_d_238;
  reg [3:0] chn_out_rsci_d_237_234;
  reg chn_out_rsci_d_222;
  reg [3:0] chn_out_rsci_d_221_218;
  reg chn_out_rsci_d_206;
  reg [3:0] chn_out_rsci_d_205_202;
  reg chn_out_rsci_d_190;
  reg [3:0] chn_out_rsci_d_189_186;
  reg chn_out_rsci_d_174;
  reg [3:0] chn_out_rsci_d_173_170;
  reg chn_out_rsci_d_158;
  reg [3:0] chn_out_rsci_d_157_154;
  reg chn_out_rsci_d_142;
  reg [3:0] chn_out_rsci_d_141_138;
  reg chn_out_rsci_d_126;
  reg [3:0] chn_out_rsci_d_125_122;
  reg chn_out_rsci_d_110;
  reg [3:0] chn_out_rsci_d_109_106;
  reg chn_out_rsci_d_94;
  reg [3:0] chn_out_rsci_d_93_90;
  reg chn_out_rsci_d_78;
  reg [3:0] chn_out_rsci_d_77_74;
  reg chn_out_rsci_d_62;
  reg [3:0] chn_out_rsci_d_61_58;
  reg chn_out_rsci_d_46;
  reg [3:0] chn_out_rsci_d_45_42;
  reg chn_out_rsci_d_30;
  reg [3:0] chn_out_rsci_d_29_26;
  reg chn_out_rsci_d_14;
  reg [3:0] chn_out_rsci_d_13_10;
  wire [1:0] fsm_output;
  wire cvt_16_FpMantRNE_24U_11U_else_and_4_tmp;
  wire cvt_15_FpMantRNE_24U_11U_else_and_3_tmp;
  wire cvt_14_FpMantRNE_24U_11U_else_and_3_tmp;
  wire cvt_13_FpMantRNE_24U_11U_else_and_2_tmp;
  wire cvt_12_FpMantRNE_24U_11U_else_and_3_tmp;
  wire cvt_11_FpMantRNE_24U_11U_else_and_2_tmp;
  wire cvt_10_FpMantRNE_24U_11U_else_and_2_tmp;
  wire cvt_9_FpMantRNE_24U_11U_else_and_1_tmp;
  wire cvt_8_FpMantRNE_24U_11U_else_and_3_tmp;
  wire cvt_7_FpMantRNE_24U_11U_else_and_2_tmp;
  wire cvt_6_FpMantRNE_24U_11U_else_and_2_tmp;
  wire cvt_5_FpMantRNE_24U_11U_else_and_1_tmp;
  wire cvt_4_FpMantRNE_24U_11U_else_and_2_tmp;
  wire cvt_3_FpMantRNE_24U_11U_else_and_1_tmp;
  wire cvt_2_FpMantRNE_24U_11U_else_and_1_tmp;
  wire cvt_1_FpMantRNE_24U_11U_else_and_tmp;
  wire cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_tmp;
  wire cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_and_9_tmp;
  wire cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_nor_20_tmp;
  wire [49:0] cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_acc_4_tmp;
  wire [50:0] nl_cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_acc_4_tmp;
  wire cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp;
  wire cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp;
  wire cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp;
  wire [49:0] cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp;
  wire [50:0] nl_cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp;
  wire cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp;
  wire cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp;
  wire cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp;
  wire [49:0] cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp;
  wire [50:0] nl_cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp;
  wire cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  wire cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  wire cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  wire [49:0] cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  wire [50:0] nl_cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  wire cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp;
  wire cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp;
  wire cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp;
  wire [49:0] cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp;
  wire [50:0] nl_cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp;
  wire cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  wire cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  wire cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  wire [49:0] cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  wire [50:0] nl_cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  wire cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  wire cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  wire cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  wire [49:0] cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  wire [50:0] nl_cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  wire cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp;
  wire cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp;
  wire cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp;
  wire [49:0] cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp;
  wire [50:0] nl_cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp;
  wire cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp;
  wire cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp;
  wire cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp;
  wire [49:0] cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp;
  wire [50:0] nl_cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp;
  wire cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  wire cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  wire cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  wire [49:0] cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  wire [50:0] nl_cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  wire cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  wire cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  wire cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  wire [49:0] cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  wire [50:0] nl_cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  wire cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp;
  wire cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp;
  wire cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp;
  wire [49:0] cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp;
  wire [50:0] nl_cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp;
  wire cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
  wire cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  wire cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  wire [49:0] cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  wire [50:0] nl_cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp;
  wire cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp;
  wire cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp;
  wire cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp;
  wire [49:0] cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp;
  wire [50:0] nl_cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp;
  wire cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp;
  wire cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp;
  wire cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp;
  wire [49:0] cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp;
  wire [50:0] nl_cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp;
  wire cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_tmp;
  wire cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_and_1_tmp;
  wire cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_nor_tmp;
  wire [49:0] cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_acc_tmp;
  wire [50:0] nl_cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_acc_tmp;
  wire cvt_16_FpMantRNE_17U_11U_else_and_4_tmp;
  wire cvt_15_FpMantRNE_17U_11U_else_and_3_tmp;
  wire cvt_14_FpMantRNE_17U_11U_else_and_3_tmp;
  wire cvt_13_FpMantRNE_17U_11U_else_and_2_tmp;
  wire cvt_12_FpMantRNE_17U_11U_else_and_3_tmp;
  wire cvt_11_FpMantRNE_17U_11U_else_and_2_tmp;
  wire cvt_10_FpMantRNE_17U_11U_else_and_2_tmp;
  wire cvt_9_FpMantRNE_17U_11U_else_and_1_tmp;
  wire cvt_8_FpMantRNE_17U_11U_else_and_3_tmp;
  wire cvt_7_FpMantRNE_17U_11U_else_and_2_tmp;
  wire cvt_6_FpMantRNE_17U_11U_else_and_2_tmp;
  wire cvt_5_FpMantRNE_17U_11U_else_and_1_tmp;
  wire cvt_4_FpMantRNE_17U_11U_else_and_2_tmp;
  wire cvt_3_FpMantRNE_17U_11U_else_and_1_tmp;
  wire cvt_2_FpMantRNE_17U_11U_else_and_1_tmp;
  wire cvt_1_FpMantRNE_17U_11U_else_and_tmp;
  wire cvt_16_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_4_tmp;
  wire cvt_15_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp;
  wire cvt_14_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp;
  wire cvt_13_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp;
  wire cvt_12_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp;
  wire cvt_11_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp;
  wire cvt_10_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp;
  wire cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp;
  wire cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp;
  wire cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp;
  wire cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp;
  wire cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp;
  wire cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp;
  wire cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp;
  wire cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp;
  wire cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_tmp;
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_15_tmp;
  wire [4:0] cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_4_tmp;
  wire [5:0] nl_cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_4_tmp;
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_14_tmp;
  wire [4:0] cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp;
  wire [5:0] nl_cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp;
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_13_tmp;
  wire [4:0] cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp;
  wire [5:0] nl_cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp;
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_12_tmp;
  wire [4:0] cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  wire [5:0] nl_cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_11_tmp;
  wire [4:0] cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp;
  wire [5:0] nl_cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp;
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_10_tmp;
  wire [4:0] cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  wire [5:0] nl_cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_9_tmp;
  wire [4:0] cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  wire [5:0] nl_cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_8_tmp;
  wire [4:0] cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp;
  wire [5:0] nl_cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp;
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_7_tmp;
  wire [4:0] cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp;
  wire [5:0] nl_cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp;
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_6_tmp;
  wire [4:0] cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  wire [5:0] nl_cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_5_tmp;
  wire [4:0] cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  wire [5:0] nl_cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  wire IsNaN_8U_23U_IsNaN_8U_23U_nand_4_tmp;
  wire IsNaN_8U_23U_nor_4_tmp;
  wire [4:0] cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp;
  wire [5:0] nl_cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp;
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_3_tmp;
  wire [4:0] cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  wire [5:0] nl_cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_2_tmp;
  wire [4:0] cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp;
  wire [5:0] nl_cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp;
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_1_tmp;
  wire [4:0] cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp;
  wire [5:0] nl_cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp;
  wire IsNaN_8U_23U_IsNaN_8U_23U_nor_tmp;
  wire [4:0] cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_tmp;
  wire [5:0] nl_cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_tmp;
  wire and_dcpl_3;
  wire and_dcpl_4;
  wire and_dcpl_70;
  wire and_dcpl_71;
  wire and_dcpl_73;
  wire and_dcpl_75;
  wire and_dcpl_77;
  wire and_dcpl_80;
  wire and_dcpl_83;
  wire or_tmp_19;
  wire mux_tmp_6;
  wire or_tmp_24;
  wire mux_tmp_39;
  wire and_tmp_8;
  wire and_tmp_11;
  wire mux_tmp_114;
  wire and_tmp_12;
  wire mux_tmp_117;
  wire and_tmp_16;
  wire or_tmp_213;
  wire mux_tmp_120;
  wire not_tmp_119;
  wire or_tmp_218;
  wire and_tmp_18;
  wire mux_tmp_122;
  wire mux_tmp_123;
  wire and_tmp_19;
  wire mux_tmp_129;
  wire and_tmp_33;
  wire mux_tmp_151;
  wire mux_tmp_161;
  wire or_tmp_306;
  wire mux_tmp_189;
  wire or_tmp_378;
  wire mux_tmp_199;
  wire mux_tmp_200;
  wire or_tmp_389;
  wire mux_tmp_236;
  wire mux_tmp_239;
  wire mux_tmp_245;
  wire and_tmp_50;
  wire and_tmp_52;
  wire mux_tmp_249;
  wire mux_tmp_251;
  wire mux_tmp_253;
  wire mux_tmp_259;
  wire mux_tmp_263;
  wire not_tmp_249;
  wire not_tmp_269;
  wire not_tmp_270;
  wire and_tmp_67;
  wire mux_tmp_294;
  wire mux_tmp_298;
  wire mux_tmp_299;
  wire mux_tmp_305;
  wire or_tmp_533;
  wire mux_tmp_309;
  wire mux_tmp_311;
  wire mux_tmp_313;
  wire mux_tmp_317;
  wire not_tmp_312;
  wire mux_tmp_321;
  wire and_tmp_71;
  wire not_tmp_336;
  wire mux_tmp_345;
  wire mux_tmp_351;
  wire mux_tmp_356;
  wire mux_tmp_370;
  wire not_tmp_388;
  wire and_tmp_79;
  wire mux_tmp_386;
  wire mux_tmp_391;
  wire mux_tmp_405;
  wire not_tmp_436;
  wire mux_tmp_415;
  wire mux_tmp_416;
  wire mux_tmp_421;
  wire mux_tmp_422;
  wire mux_tmp_427;
  wire mux_tmp_428;
  wire mux_tmp_435;
  wire mux_tmp_440;
  wire mux_tmp_441;
  wire not_tmp_497;
  wire and_tmp_93;
  wire mux_tmp_455;
  wire and_tmp_94;
  wire not_tmp_520;
  wire mux_tmp_481;
  wire mux_tmp_487;
  wire mux_tmp_502;
  wire not_tmp_580;
  wire mux_tmp_519;
  wire mux_tmp_525;
  wire mux_tmp_541;
  wire not_tmp_638;
  wire mux_tmp_560;
  wire mux_tmp_565;
  wire mux_tmp_566;
  wire mux_tmp_577;
  wire mux_tmp_578;
  wire mux_tmp_579;
  wire mux_tmp_580;
  wire mux_tmp_585;
  wire mux_tmp_591;
  wire mux_tmp_592;
  wire mux_tmp_597;
  wire mux_tmp_600;
  wire mux_tmp_601;
  wire mux_tmp_602;
  wire mux_tmp_612;
  wire mux_tmp_613;
  wire mux_tmp_614;
  wire not_tmp_757;
  wire mux_tmp_634;
  wire mux_tmp_638;
  wire mux_tmp_639;
  wire mux_tmp_640;
  wire mux_tmp_641;
  wire not_tmp_811;
  wire mux_tmp_658;
  wire mux_tmp_678;
  wire mux_tmp_679;
  wire mux_tmp_680;
  wire mux_tmp_681;
  wire mux_tmp_692;
  wire mux_tmp_693;
  wire mux_tmp_694;
  wire mux_tmp_695;
  wire not_tmp_899;
  wire mux_tmp_719;
  wire mux_tmp_720;
  wire mux_tmp_723;
  wire mux_tmp_724;
  wire mux_tmp_725;
  wire mux_tmp_726;
  wire mux_tmp_727;
  wire mux_tmp_739;
  wire mux_tmp_740;
  wire mux_tmp_741;
  wire mux_tmp_742;
  wire mux_tmp_743;
  wire not_tmp_989;
  wire mux_tmp_765;
  wire mux_tmp_766;
  wire or_tmp_1375;
  wire or_tmp_1393;
  wire mux_tmp_944;
  wire mux_tmp_945;
  wire and_tmp_165;
  wire mux_tmp_946;
  wire mux_tmp_947;
  wire and_tmp_166;
  wire mux_tmp_960;
  wire mux_tmp_961;
  wire and_tmp_168;
  wire mux_tmp_962;
  wire mux_tmp_963;
  wire and_tmp_169;
  wire mux_tmp_986;
  wire mux_tmp_987;
  wire mux_tmp_992;
  wire mux_tmp_994;
  wire mux_tmp_1015;
  wire mux_tmp_1038;
  wire nand_tmp_30;
  wire mux_tmp_1039;
  wire and_tmp_171;
  wire or_tmp_1650;
  wire mux_tmp_1041;
  wire mux_tmp_1043;
  wire mux_tmp_1047;
  wire mux_tmp_1049;
  wire mux_tmp_1074;
  wire mux_tmp_1088;
  wire mux_tmp_1100;
  wire nand_tmp_36;
  wire mux_tmp_1101;
  wire and_tmp_175;
  wire or_tmp_1780;
  wire mux_tmp_1103;
  wire mux_tmp_1105;
  wire mux_tmp_1109;
  wire mux_tmp_1111;
  wire mux_tmp_1152;
  wire mux_tmp_1196;
  wire mux_tmp_1197;
  wire or_tmp_1981;
  wire or_tmp_1992;
  wire mux_tmp_1225;
  wire mux_tmp_1226;
  wire mux_tmp_1227;
  wire mux_tmp_1264;
  wire or_tmp_2136;
  wire or_tmp_2139;
  wire mux_tmp_1270;
  wire mux_tmp_1276;
  wire mux_tmp_1280;
  wire mux_tmp_1282;
  wire mux_tmp_1326;
  wire mux_tmp_1332;
  wire mux_tmp_1337;
  wire mux_tmp_1339;
  wire mux_tmp_1341;
  wire mux_tmp_1409;
  wire mux_tmp_1419;
  wire not_tmp_1709;
  wire nand_tmp_48;
  wire mux_tmp_1435;
  wire mux_tmp_1469;
  wire or_tmp_2432;
  wire or_tmp_2466;
  wire or_tmp_2469;
  wire mux_tmp_1566;
  wire or_tmp_2569;
  wire mux_tmp_1570;
  wire or_tmp_2571;
  wire mux_tmp_1574;
  wire or_tmp_2573;
  wire mux_tmp_1578;
  wire or_tmp_2575;
  wire mux_tmp_1582;
  wire or_tmp_2577;
  wire mux_tmp_1586;
  wire or_tmp_2579;
  wire mux_tmp_1592;
  wire or_tmp_2588;
  wire mux_tmp_1596;
  wire or_tmp_2590;
  wire mux_tmp_1600;
  wire or_tmp_2595;
  wire mux_tmp_1606;
  wire or_tmp_2604;
  wire mux_tmp_1610;
  wire or_tmp_2606;
  wire mux_tmp_1614;
  wire or_tmp_2608;
  wire mux_tmp_1618;
  wire or_tmp_2610;
  wire mux_tmp_1622;
  wire or_tmp_2612;
  wire and_dcpl_93;
  wire or_dcpl_4;
  wire and_dcpl_98;
  wire and_dcpl_102;
  wire and_dcpl_103;
  wire and_dcpl_105;
  wire and_dcpl_114;
  wire or_dcpl_15;
  wire or_dcpl_16;
  wire or_dcpl_30;
  wire or_dcpl_32;
  wire and_dcpl_204;
  wire and_dcpl_209;
  wire and_dcpl_217;
  wire and_dcpl_224;
  wire or_dcpl_108;
  wire and_dcpl_228;
  wire or_dcpl_109;
  wire nor_tmp_636;
  wire or_dcpl_110;
  wire or_dcpl_111;
  wire not_tmp_2254;
  wire or_tmp_2960;
  wire or_dcpl_113;
  wire or_dcpl_114;
  wire and_tmp_225;
  wire or_dcpl_115;
  wire or_dcpl_116;
  wire or_dcpl_119;
  wire or_dcpl_120;
  wire and_dcpl_301;
  wire or_dcpl_124;
  wire or_dcpl_125;
  wire or_dcpl_126;
  wire or_dcpl_127;
  wire or_dcpl_130;
  wire or_dcpl_131;
  wire or_dcpl_132;
  wire or_dcpl_133;
  wire or_tmp_3025;
  wire or_tmp_3032;
  wire or_dcpl_136;
  wire and_dcpl_363;
  wire or_dcpl_137;
  wire or_dcpl_139;
  wire or_dcpl_140;
  wire or_dcpl_143;
  wire or_dcpl_144;
  wire mux_tmp_1813;
  wire and_dcpl_401;
  wire and_dcpl_407;
  wire and_dcpl_408;
  wire or_dcpl_147;
  wire and_dcpl_409;
  wire and_dcpl_411;
  wire and_dcpl_417;
  wire and_dcpl_420;
  wire and_dcpl_424;
  wire and_dcpl_425;
  wire and_dcpl_433;
  wire or_dcpl_151;
  wire and_dcpl_444;
  wire and_dcpl_446;
  wire not_tmp_2422;
  wire and_dcpl_458;
  wire and_tmp_248;
  wire or_dcpl_160;
  wire and_dcpl_473;
  wire and_dcpl_479;
  wire or_dcpl_163;
  wire and_dcpl_481;
  wire mux_tmp_1899;
  wire and_dcpl_499;
  wire or_dcpl_178;
  wire and_dcpl_535;
  wire or_dcpl_181;
  wire or_dcpl_184;
  wire or_dcpl_188;
  wire or_dcpl_195;
  wire or_dcpl_197;
  wire or_dcpl_210;
  wire and_dcpl_617;
  wire and_dcpl_626;
  wire or_dcpl_243;
  wire and_dcpl_631;
  wire and_dcpl_648;
  wire or_tmp_3379;
  wire or_dcpl_277;
  wire or_dcpl_320;
  wire or_dcpl_322;
  wire or_dcpl_324;
  wire or_dcpl_326;
  wire or_dcpl_328;
  wire or_dcpl_330;
  wire or_dcpl_332;
  wire or_dcpl_334;
  wire or_dcpl_336;
  wire or_dcpl_338;
  wire or_dcpl_340;
  wire or_dcpl_342;
  wire or_dcpl_344;
  wire or_dcpl_346;
  wire or_dcpl_348;
  wire or_dcpl_350;
  wire or_dcpl_353;
  wire or_dcpl_386;
  wire or_dcpl_389;
  wire and_dcpl_942;
  wire or_dcpl_399;
  wire and_dcpl_946;
  wire and_dcpl_950;
  wire or_dcpl_420;
  wire and_dcpl_954;
  wire and_dcpl_958;
  wire or_dcpl_439;
  wire and_dcpl_962;
  wire or_dcpl_448;
  wire and_dcpl_966;
  wire and_dcpl_970;
  wire and_dcpl_974;
  wire or_dcpl_480;
  wire and_dcpl_978;
  wire or_dcpl_490;
  wire and_dcpl_982;
  wire and_dcpl_987;
  wire or_dcpl_511;
  wire and_dcpl_991;
  wire and_dcpl_995;
  wire and_dcpl_999;
  wire and_dcpl_1003;
  wire or_dcpl_612;
  wire or_tmp_3487;
  reg cvt_1_FpMantRNE_24U_11U_else_and_svs;
  reg cvt_2_FpMantRNE_24U_11U_else_and_1_svs;
  reg cvt_3_FpMantRNE_24U_11U_else_and_1_svs;
  reg cvt_4_FpMantRNE_24U_11U_else_and_2_svs;
  reg cvt_5_FpMantRNE_24U_11U_else_and_1_svs;
  reg cvt_6_FpMantRNE_24U_11U_else_and_2_svs;
  reg cvt_7_FpMantRNE_24U_11U_else_and_2_svs;
  reg cvt_8_FpMantRNE_24U_11U_else_and_3_svs;
  reg cvt_9_FpMantRNE_24U_11U_else_and_1_svs;
  reg cvt_10_FpMantRNE_24U_11U_else_and_2_svs;
  reg cvt_11_FpMantRNE_24U_11U_else_and_2_svs;
  reg cvt_12_FpMantRNE_24U_11U_else_and_3_svs;
  reg cvt_13_FpMantRNE_24U_11U_else_and_2_svs;
  reg cvt_14_FpMantRNE_24U_11U_else_and_3_svs;
  reg cvt_15_FpMantRNE_24U_11U_else_and_3_svs;
  reg cvt_16_FpMantRNE_24U_11U_else_and_4_svs;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_1_sva;
  reg IntShiftRightSat_49U_6U_17U_lor_2_lpi_1_dfm;
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp;
  reg cvt_1_FpMantRNE_17U_11U_else_and_svs;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_2_sva;
  reg IntShiftRightSat_49U_6U_17U_o_16_2_sva;
  reg IntShiftRightSat_49U_6U_17U_lor_3_lpi_1_dfm;
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_1;
  reg cvt_2_FpMantRNE_17U_11U_else_and_1_svs;
  reg cvt_else_equal_tmp_5;
  reg cvt_else_nor_dfs_2;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_3_sva;
  reg IntShiftRightSat_49U_6U_17U_lor_4_lpi_1_dfm;
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_2;
  reg cvt_3_FpMantRNE_17U_11U_else_and_1_svs;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_4_sva;
  reg IntShiftRightSat_49U_6U_17U_o_16_4_sva;
  reg IntShiftRightSat_49U_6U_17U_lor_5_lpi_1_dfm;
  reg cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs;
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_3;
  reg cvt_4_FpMantRNE_17U_11U_else_and_2_svs;
  reg FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_3;
  reg cvt_else_equal_tmp_9;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_5_sva;
  reg IntShiftRightSat_49U_6U_17U_lor_6_lpi_1_dfm;
  reg cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs;
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_4;
  reg cvt_5_FpMantRNE_17U_11U_else_and_1_svs;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_6_sva;
  reg IntShiftRightSat_49U_6U_17U_o_16_6_sva;
  reg IntShiftRightSat_49U_6U_17U_lor_7_lpi_1_dfm;
  reg cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs;
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_5;
  reg cvt_6_FpMantRNE_17U_11U_else_and_2_svs;
  reg FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_3;
  reg cvt_else_equal_tmp_16;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_7_sva;
  reg IntShiftRightSat_49U_6U_17U_o_16_7_sva;
  reg IntShiftRightSat_49U_6U_17U_lor_8_lpi_1_dfm;
  reg cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs;
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_6;
  reg cvt_7_FpMantRNE_17U_11U_else_and_2_svs;
  reg FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_3;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_8_sva;
  reg IntShiftRightSat_49U_6U_17U_o_16_8_sva;
  reg IntShiftRightSat_49U_6U_17U_lor_9_lpi_1_dfm;
  reg cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs;
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_7;
  reg cvt_8_FpMantRNE_17U_11U_else_and_3_svs;
  reg FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_3;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_9_sva;
  reg IntShiftRightSat_49U_6U_17U_lor_10_lpi_1_dfm;
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_8;
  reg cvt_9_FpMantRNE_17U_11U_else_and_1_svs;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_10_sva;
  reg IntShiftRightSat_49U_6U_17U_o_16_10_sva;
  reg IntShiftRightSat_49U_6U_17U_lor_11_lpi_1_dfm;
  reg cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs;
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_9;
  reg cvt_10_FpMantRNE_17U_11U_else_and_2_svs;
  reg FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_3;
  reg cvt_else_equal_tmp_28;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_11_sva;
  reg IntShiftRightSat_49U_6U_17U_o_16_11_sva;
  reg IntShiftRightSat_49U_6U_17U_lor_12_lpi_1_dfm;
  reg cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs;
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_10;
  reg cvt_11_FpMantRNE_17U_11U_else_and_2_svs;
  reg FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_3;
  reg cvt_else_nor_dfs_10;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_12_sva;
  reg IntShiftRightSat_49U_6U_17U_o_16_12_sva;
  reg IntShiftRightSat_49U_6U_17U_lor_13_lpi_1_dfm;
  reg cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs;
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_11;
  reg cvt_12_FpMantRNE_17U_11U_else_and_3_svs;
  reg FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_3;
  reg cvt_else_equal_tmp_33;
  reg cvt_else_equal_tmp_34;
  reg cvt_else_nor_dfs_11;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_13_sva;
  reg IntShiftRightSat_49U_6U_17U_o_16_13_sva;
  reg IntShiftRightSat_49U_6U_17U_lor_14_lpi_1_dfm;
  reg cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs;
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_12;
  reg cvt_13_FpMantRNE_17U_11U_else_and_2_svs;
  reg FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_3;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_14_sva;
  reg IntShiftRightSat_49U_6U_17U_o_16_14_sva;
  reg IntShiftRightSat_49U_6U_17U_lor_15_lpi_1_dfm;
  reg cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs;
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_13;
  reg cvt_14_FpMantRNE_17U_11U_else_and_3_svs;
  reg FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2;
  reg chn_odata_data_13_0_lpi_1_dfm_1;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_15_sva;
  reg IntShiftRightSat_49U_6U_17U_o_16_15_sva;
  reg IntShiftRightSat_49U_6U_17U_lor_16_lpi_1_dfm;
  reg cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs;
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_14;
  reg cvt_15_FpMantRNE_17U_11U_else_and_3_svs;
  reg FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_3;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_sva;
  reg IntShiftRightSat_49U_6U_17U_o_16_sva;
  reg IntShiftRightSat_49U_6U_17U_lor_lpi_1_dfm;
  reg cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_svs;
  reg FpIntToFloat_17U_5U_10U_else_unequal_tmp_15;
  reg cvt_16_FpMantRNE_17U_11U_else_and_4_svs;
  reg FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_3;
  reg cvt_else_equal_tmp_45;
  reg cvt_else_equal_tmp_46;
  reg cvt_else_nor_dfs_15;
  reg main_stage_v_1;
  reg main_stage_v_2;
  reg main_stage_v_3;
  reg IsNaN_5U_10U_land_1_lpi_1_dfm_3;
  reg cvt_1_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_svs_2;
  reg IntShiftRightSat_49U_6U_17U_o_0_1_sva_2;
  reg IsNaN_5U_10U_land_2_lpi_1_dfm_4;
  reg cvt_2_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2;
  reg IsNaN_5U_10U_land_4_lpi_1_dfm_4;
  reg IsNaN_5U_10U_land_4_lpi_1_dfm_5;
  reg cvt_4_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2;
  reg IsNaN_5U_10U_land_7_lpi_1_dfm_5;
  reg IsNaN_5U_10U_land_7_lpi_1_dfm_6;
  reg cvt_7_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2;
  reg IntShiftRightSat_49U_6U_17U_o_0_7_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_0_7_sva_3;
  reg IsNaN_5U_10U_land_8_lpi_1_dfm_4;
  reg IsNaN_5U_10U_land_8_lpi_1_dfm_5;
  reg cvt_8_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2;
  reg IsNaN_5U_10U_land_11_lpi_1_dfm_4;
  reg IsNaN_5U_10U_land_11_lpi_1_dfm_5;
  reg cvt_11_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2;
  reg IntShiftRightSat_49U_6U_17U_o_0_11_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_0_11_sva_3;
  reg IsNaN_5U_10U_land_13_lpi_1_dfm_4;
  reg IsNaN_5U_10U_land_13_lpi_1_dfm_5;
  reg cvt_13_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2;
  reg IntShiftRightSat_49U_6U_17U_o_0_13_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_0_13_sva_3;
  reg IsNaN_5U_10U_land_14_lpi_1_dfm_5;
  reg IsNaN_5U_10U_land_14_lpi_1_dfm_6;
  reg cvt_14_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2;
  reg IsNaN_5U_10U_land_lpi_1_dfm_4;
  reg IsNaN_5U_10U_land_lpi_1_dfm_5;
  reg cvt_16_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_4_svs_2;
  reg IsNaN_5U_10U_land_15_lpi_1_dfm_3;
  reg cvt_15_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2;
  reg IntShiftRightSat_49U_6U_17U_o_0_15_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_0_15_sva_3;
  reg IsNaN_5U_10U_land_12_lpi_1_dfm_4;
  reg IsNaN_5U_10U_land_12_lpi_1_dfm_5;
  reg cvt_12_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2;
  reg IsNaN_5U_10U_land_10_lpi_1_dfm_4;
  reg IsNaN_5U_10U_land_10_lpi_1_dfm_5;
  reg cvt_10_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2;
  reg IsNaN_5U_10U_land_9_lpi_1_dfm_4;
  reg IsNaN_5U_10U_land_9_lpi_1_dfm_5;
  reg cvt_9_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2;
  reg IntShiftRightSat_49U_6U_17U_o_0_9_sva_3;
  reg IntShiftRightSat_49U_6U_17U_o_0_9_sva_4;
  reg IsNaN_5U_10U_land_6_lpi_1_dfm_4;
  reg IsNaN_5U_10U_land_6_lpi_1_dfm_5;
  reg cvt_6_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2;
  reg IsNaN_5U_10U_land_5_lpi_1_dfm_4;
  reg IsNaN_5U_10U_land_5_lpi_1_dfm_5;
  reg cvt_5_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2;
  reg IntShiftRightSat_49U_6U_17U_o_0_5_sva_3;
  reg IntShiftRightSat_49U_6U_17U_o_0_5_sva_4;
  reg IsNaN_5U_10U_land_3_lpi_1_dfm_4;
  reg IsNaN_5U_10U_land_3_lpi_1_dfm_5;
  reg cvt_3_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2;
  reg IntShiftRightSat_49U_6U_17U_o_0_3_sva_3;
  reg IntShiftRightSat_49U_6U_17U_o_0_3_sva_4;
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_1_lpi_1_dfm_8;
  reg IntShiftRightSat_49U_6U_17U_o_16_1_sva_3;
  reg IntShiftRightSat_49U_6U_17U_o_16_1_sva_4;
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_2_lpi_1_dfm_8;
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_4_lpi_1_dfm_8;
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_7_lpi_1_dfm_8;
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_8_lpi_1_dfm_8;
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_11_lpi_1_dfm_8;
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_13_lpi_1_dfm_8;
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_14_lpi_1_dfm_8;
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_15_lpi_1_dfm_8;
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_12_lpi_1_dfm_8;
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_10_lpi_1_dfm_8;
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_9_lpi_1_dfm_8;
  reg IntShiftRightSat_49U_6U_17U_o_16_9_sva_3;
  reg IntShiftRightSat_49U_6U_17U_o_16_9_sva_4;
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_6_lpi_1_dfm_8;
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_5_lpi_1_dfm_8;
  reg IntShiftRightSat_49U_6U_17U_o_16_5_sva_3;
  reg IntShiftRightSat_49U_6U_17U_o_16_5_sva_4;
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_3_lpi_1_dfm_8;
  reg IntShiftRightSat_49U_6U_17U_o_16_3_sva_3;
  reg IntShiftRightSat_49U_6U_17U_o_16_3_sva_4;
  reg IntShiftRightSat_49U_6U_17U_o_0_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_0_sva_3;
  reg cvt_14_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_3_svs_1;
  reg IntShiftRightSat_49U_6U_17U_o_0_14_sva_3;
  reg IntShiftRightSat_49U_6U_17U_o_0_14_sva_4;
  reg IntShiftRightSat_49U_6U_17U_o_0_12_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_0_12_sva_3;
  reg IntShiftRightSat_49U_6U_17U_o_0_10_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_0_8_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_0_8_sva_3;
  reg IntShiftRightSat_49U_6U_17U_o_0_6_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_0_6_sva_3;
  reg IntShiftRightSat_49U_6U_17U_o_0_4_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_0_4_sva_3;
  reg IntShiftRightSat_49U_6U_17U_o_0_2_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_0_2_sva_3;
  reg FpFloatToInt_16U_5U_10U_internal_int_0_sva_3;
  reg FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_2;
  reg FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_2;
  reg FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_2;
  reg FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_2;
  reg FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_2;
  reg FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_2;
  reg FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_2;
  reg FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_2;
  reg FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_2;
  reg FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_2;
  reg FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_2;
  reg FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_2;
  reg FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_2;
  reg FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_2;
  reg FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_2;
  reg [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_lpi_1_dfm_9;
  reg [14:0] IntSaturation_17U_16U_o_15_1_lpi_1_dfm_9;
  reg [14:0] IntSaturation_17U_16U_o_15_1_15_lpi_1_dfm_8;
  reg [14:0] IntSaturation_17U_16U_o_15_1_14_lpi_1_dfm_8;
  reg [14:0] IntSaturation_17U_16U_o_15_1_13_lpi_1_dfm_7;
  reg [14:0] IntSaturation_17U_16U_o_15_1_12_lpi_1_dfm_8;
  reg [14:0] IntSaturation_17U_16U_o_15_1_11_lpi_1_dfm_7;
  reg [14:0] IntSaturation_17U_16U_o_15_1_10_lpi_1_dfm_7;
  reg [14:0] IntSaturation_17U_16U_o_15_1_9_lpi_1_dfm_6;
  reg [14:0] IntSaturation_17U_16U_o_15_1_8_lpi_1_dfm_8;
  reg [14:0] IntSaturation_17U_16U_o_15_1_7_lpi_1_dfm_7;
  reg [14:0] IntSaturation_17U_16U_o_15_1_6_lpi_1_dfm_7;
  reg [14:0] IntSaturation_17U_16U_o_15_1_5_lpi_1_dfm_6;
  reg [14:0] IntSaturation_17U_16U_o_15_1_4_lpi_1_dfm_7;
  reg [14:0] IntSaturation_17U_16U_o_15_1_3_lpi_1_dfm_6;
  reg [14:0] IntSaturation_17U_16U_o_15_1_2_lpi_1_dfm_6;
  reg [14:0] IntSaturation_17U_16U_o_15_1_1_lpi_1_dfm_5;
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_sva_9;
  reg cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_2;
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_sva_9;
  reg cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_2;
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_sva_9;
  reg cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_2;
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_sva_9;
  reg cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_2;
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_sva_9;
  reg cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_2;
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_sva_9;
  reg cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_2;
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_sva_9;
  reg cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_2;
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_sva_9;
  reg cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_2;
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_sva_9;
  reg cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_2;
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_sva_9;
  reg cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_2;
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_sva_9;
  reg cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_2;
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_sva_9;
  reg cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_2;
  reg [14:0] FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5;
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_sva_9;
  reg cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_2;
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_sva_9;
  reg cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_2;
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_sva_9;
  reg cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_2;
  reg [4:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_sva_9;
  reg cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_2;
  reg [5:0] cfg_truncate_1_sva_2;
  reg [1:0] cfg_out_precision_1_sva_6;
  reg cfg_mode_eql_1_sva_4;
  reg cfg_mode_eql_1_sva_5;
  reg cfg_mode_eql_1_sva_6;
  reg cvt_unequal_tmp_19;
  reg cvt_unequal_tmp_20;
  reg cvt_unequal_tmp_21;
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_2_sva_2;
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_1_sva_2;
  wire [5:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_1_sva_2;
  reg FpMantRNE_24U_11U_else_carry_1_sva_2;
  reg cvt_1_FpMantRNE_24U_11U_else_and_svs_2;
  reg IsNaN_8U_23U_land_1_lpi_1_dfm_3;
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_3_sva_2;
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_2_sva_2;
  wire [5:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_2_sva_2;
  reg FpMantRNE_24U_11U_else_carry_2_sva_2;
  reg cvt_2_FpMantRNE_24U_11U_else_and_1_svs_2;
  reg IsNaN_8U_23U_land_2_lpi_1_dfm_3;
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_4_sva_2;
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_3_sva_2;
  wire [5:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_3_sva_2;
  reg FpMantRNE_24U_11U_else_carry_3_sva_2;
  reg cvt_3_FpMantRNE_24U_11U_else_and_1_svs_2;
  reg IsNaN_8U_23U_land_3_lpi_1_dfm_3;
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_5_sva_2;
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_4_sva_2;
  wire [5:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_4_sva_2;
  reg FpMantRNE_24U_11U_else_carry_4_sva_2;
  reg cvt_4_FpMantRNE_24U_11U_else_and_2_svs_2;
  reg IsNaN_8U_23U_land_4_lpi_1_dfm_3;
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_6_sva_2;
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_5_sva_2;
  wire [5:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_5_sva_2;
  reg FpMantRNE_24U_11U_else_carry_5_sva_2;
  reg cvt_5_FpMantRNE_24U_11U_else_and_1_svs_2;
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_7_sva_2;
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_6_sva_2;
  wire [5:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_6_sva_2;
  reg FpMantRNE_24U_11U_else_carry_6_sva_2;
  reg cvt_6_FpMantRNE_24U_11U_else_and_2_svs_2;
  reg IsNaN_8U_23U_land_6_lpi_1_dfm_3;
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_8_sva_2;
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_7_sva_2;
  wire [5:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_7_sva_2;
  reg FpMantRNE_24U_11U_else_carry_7_sva_2;
  reg cvt_7_FpMantRNE_24U_11U_else_and_2_svs_2;
  reg IsNaN_8U_23U_land_7_lpi_1_dfm_3;
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_9_sva_2;
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_8_sva_2;
  wire [5:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_8_sva_2;
  reg FpMantRNE_24U_11U_else_carry_8_sva_2;
  reg cvt_8_FpMantRNE_24U_11U_else_and_3_svs_2;
  reg IsNaN_8U_23U_land_8_lpi_1_dfm_3;
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_10_sva_2;
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_9_sva_2;
  wire [5:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_9_sva_2;
  reg FpMantRNE_24U_11U_else_carry_9_sva_2;
  reg cvt_9_FpMantRNE_24U_11U_else_and_1_svs_2;
  reg IsNaN_8U_23U_land_9_lpi_1_dfm_3;
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_11_sva_2;
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_10_sva_2;
  wire [5:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_10_sva_2;
  reg FpMantRNE_24U_11U_else_carry_10_sva_2;
  reg cvt_10_FpMantRNE_24U_11U_else_and_2_svs_2;
  reg IsNaN_8U_23U_land_10_lpi_1_dfm_3;
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_12_sva_2;
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_11_sva_2;
  wire [5:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_11_sva_2;
  reg FpMantRNE_24U_11U_else_carry_11_sva_2;
  reg cvt_11_FpMantRNE_24U_11U_else_and_2_svs_2;
  reg IsNaN_8U_23U_land_11_lpi_1_dfm_3;
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_13_sva_2;
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_12_sva_2;
  wire [5:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_12_sva_2;
  reg FpMantRNE_24U_11U_else_carry_12_sva_2;
  reg cvt_12_FpMantRNE_24U_11U_else_and_3_svs_2;
  reg IsNaN_8U_23U_land_12_lpi_1_dfm_3;
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_14_sva_2;
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_13_sva_2;
  wire [5:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_13_sva_2;
  reg FpMantRNE_24U_11U_else_carry_13_sva_2;
  reg cvt_13_FpMantRNE_24U_11U_else_and_2_svs_2;
  reg IsNaN_8U_23U_land_13_lpi_1_dfm_3;
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_15_sva_2;
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_14_sva_2;
  wire [5:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_14_sva_2;
  reg FpMantRNE_24U_11U_else_carry_14_sva_2;
  reg cvt_14_FpMantRNE_24U_11U_else_and_3_svs_2;
  reg IsNaN_8U_23U_land_14_lpi_1_dfm_3;
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_16_sva_2;
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_15_sva_2;
  wire [5:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_15_sva_2;
  reg FpMantRNE_24U_11U_else_carry_15_sva_2;
  reg cvt_15_FpMantRNE_24U_11U_else_and_3_svs_2;
  reg IsNaN_8U_23U_land_15_lpi_1_dfm_3;
  reg [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_2;
  reg [4:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva_2;
  wire [5:0] nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva_2;
  reg FpMantRNE_24U_11U_else_carry_sva_2;
  reg cvt_16_FpMantRNE_24U_11U_else_and_4_svs_2;
  reg IsNaN_8U_23U_land_lpi_1_dfm_3;
  reg [48:0] IntMulExt_33U_16U_49U_return_1_sva_2;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_2;
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_1_sva_2;
  reg cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_svs_2;
  reg [14:0] FpIntToFloat_17U_5U_10U_else_i_abs_15_1_1_lpi_1_dfm_5;
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_1_lpi_1_dfm_5;
  reg FpIntToFloat_17U_5U_10U_is_inf_1_lpi_1_dfm_6;
  reg [48:0] IntMulExt_33U_16U_49U_return_2_sva_2;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_16_2_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_16_2_sva_3;
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_2_sva_2;
  reg cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  reg [14:0] FpIntToFloat_17U_5U_10U_else_i_abs_15_1_2_lpi_1_dfm_6;
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_2_lpi_1_dfm_6;
  reg FpIntToFloat_17U_5U_10U_is_inf_2_lpi_1_dfm_6;
  reg [48:0] IntMulExt_33U_16U_49U_return_3_sva_2;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_2;
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_3_sva_2;
  reg cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  reg [14:0] FpIntToFloat_17U_5U_10U_else_i_abs_15_1_3_lpi_1_dfm_6;
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_3_lpi_1_dfm_6;
  reg FpIntToFloat_17U_5U_10U_is_inf_3_lpi_1_dfm_7;
  reg [48:0] IntMulExt_33U_16U_49U_return_4_sva_1;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_16_4_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_16_4_sva_3;
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_4_sva_2;
  reg cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_4_lpi_1_dfm_7;
  reg FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_7;
  reg [48:0] IntMulExt_33U_16U_49U_return_5_sva_2;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_2;
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_5_sva_2;
  reg cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_5_lpi_1_dfm_6;
  reg FpIntToFloat_17U_5U_10U_is_inf_5_lpi_1_dfm_7;
  reg [48:0] IntMulExt_33U_16U_49U_return_6_sva_1;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_16_6_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_16_6_sva_3;
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_6_sva_2;
  reg cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_6_lpi_1_dfm_7;
  reg FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_7;
  reg [48:0] IntMulExt_33U_16U_49U_return_7_sva_1;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_16_7_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_16_7_sva_3;
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_7_sva_2;
  reg cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_7_lpi_1_dfm_7;
  reg FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_7;
  reg [48:0] IntMulExt_33U_16U_49U_return_8_sva_1;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_16_8_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_16_8_sva_3;
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_8_sva_2;
  reg cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_8_lpi_1_dfm_8;
  reg FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_8;
  reg [48:0] IntMulExt_33U_16U_49U_return_9_sva_2;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_2;
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_9_sva_2;
  reg cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_2;
  reg cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  reg [14:0] FpIntToFloat_17U_5U_10U_else_i_abs_15_1_9_lpi_1_dfm_6;
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_9_lpi_1_dfm_6;
  reg FpIntToFloat_17U_5U_10U_is_inf_9_lpi_1_dfm_7;
  reg [48:0] IntMulExt_33U_16U_49U_return_10_sva_1;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_16_10_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_16_10_sva_3;
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_10_sva_2;
  reg cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_10_lpi_1_dfm_7;
  reg FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_7;
  reg [48:0] IntMulExt_33U_16U_49U_return_11_sva_1;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_16_11_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_16_11_sva_3;
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_11_sva_2;
  reg cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_11_lpi_1_dfm_7;
  reg FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_7;
  reg [48:0] IntMulExt_33U_16U_49U_return_12_sva_1;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_16_12_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_16_12_sva_3;
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_12_sva_2;
  reg cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_12_lpi_1_dfm_8;
  reg FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_8;
  reg [48:0] IntMulExt_33U_16U_49U_return_13_sva_1;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_16_13_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_16_13_sva_3;
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_13_sva_2;
  reg cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_13_lpi_1_dfm_7;
  reg FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_7;
  reg [48:0] IntMulExt_33U_16U_49U_return_14_sva_1;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_16_14_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_16_14_sva_3;
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_14_sva_2;
  reg cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_14_lpi_1_dfm_8;
  reg FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_8;
  reg [48:0] IntMulExt_33U_16U_49U_return_15_sva_1;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_16_15_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_16_15_sva_3;
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_15_sva_2;
  reg cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_15_lpi_1_dfm_8;
  reg FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_8;
  reg [48:0] IntMulExt_33U_16U_49U_return_sva_1;
  reg [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_16_sva_2;
  reg IntShiftRightSat_49U_6U_17U_o_16_sva_3;
  reg [48:0] IntShiftRightSat_49U_6U_17U_i_sva_2;
  reg cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_svs_2;
  reg FpIntToFloat_17U_5U_10U_else_i_abs_0_lpi_1_dfm_9;
  reg FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_9;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_itm_2;
  reg [4:0] cvt_1_FpFloatToInt_16U_5U_10U_shift_acc_itm_2;
  wire [5:0] nl_cvt_1_FpFloatToInt_16U_5U_10U_shift_acc_itm_2;
  reg IsNaN_5U_10U_nor_itm_2;
  reg IsNaN_5U_10U_IsNaN_5U_10U_nand_itm_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_1_itm_2;
  reg [4:0] cvt_2_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2;
  wire [5:0] nl_cvt_2_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2;
  reg IsNaN_5U_10U_nor_1_itm_2;
  reg IsNaN_5U_10U_IsNaN_5U_10U_nand_1_itm_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_2_itm_2;
  reg [4:0] cvt_3_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2;
  wire [5:0] nl_cvt_3_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_3_itm_2;
  reg [4:0] cvt_4_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  wire [5:0] nl_cvt_4_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_4_itm_2;
  reg IsNaN_8U_23U_nor_4_itm_2;
  reg IsNaN_8U_23U_IsNaN_8U_23U_nand_4_itm_2;
  reg [4:0] cvt_5_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2;
  wire [5:0] nl_cvt_5_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_5_itm_2;
  reg [4:0] cvt_6_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  wire [5:0] nl_cvt_6_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_6_itm_2;
  reg [4:0] cvt_7_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  wire [5:0] nl_cvt_7_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_7_itm_2;
  reg [4:0] cvt_8_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2;
  wire [5:0] nl_cvt_8_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_8_itm_2;
  reg [4:0] cvt_9_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2;
  wire [5:0] nl_cvt_9_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_9_itm_2;
  reg [4:0] cvt_10_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  wire [5:0] nl_cvt_10_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_10_itm_2;
  reg [4:0] cvt_11_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  wire [5:0] nl_cvt_11_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_11_itm_2;
  reg [4:0] cvt_12_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2;
  wire [5:0] nl_cvt_12_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_12_itm_2;
  reg [4:0] cvt_13_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  wire [5:0] nl_cvt_13_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_13_itm_2;
  reg [4:0] cvt_14_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2;
  wire [5:0] nl_cvt_14_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_14_itm_2;
  reg [4:0] cvt_15_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2;
  wire [5:0] nl_cvt_15_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2;
  reg IsNaN_5U_10U_nor_14_itm_2;
  reg IsNaN_5U_10U_IsNaN_5U_10U_nand_14_itm_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_nand_15_itm_2;
  reg [4:0] cvt_16_FpFloatToInt_16U_5U_10U_shift_acc_4_itm_2;
  wire [5:0] nl_cvt_16_FpFloatToInt_16U_5U_10U_shift_acc_4_itm_2;
  reg cvt_1_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_itm_2;
  reg cvt_2_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2;
  reg cvt_3_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2;
  reg [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_7_itm_1;
  reg cvt_4_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2;
  reg cvt_5_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2;
  reg cvt_6_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2;
  reg cvt_7_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2;
  reg cvt_8_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2;
  reg cvt_9_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2;
  reg cvt_10_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2;
  reg cvt_11_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2;
  reg cvt_12_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2;
  reg cvt_13_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2;
  reg cvt_14_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2;
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm;
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm_3;
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm_4;
  reg cvt_15_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2;
  reg cvt_16_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_4_itm_2;
  reg cvt_16_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  reg cvt_15_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  reg cvt_14_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  reg cvt_13_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  reg cvt_12_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  reg cvt_11_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  reg cvt_10_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  reg cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  reg cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  reg cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  reg cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  reg cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  reg cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  reg cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  reg cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  reg cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2;
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_15_itm_2;
  reg cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1;
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_14_itm_2;
  reg cvt_15_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_2;
  reg cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1;
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_12_itm_2;
  reg cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1;
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_11_itm_2;
  reg cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1;
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_10_itm_2;
  reg cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1;
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_9_itm_2;
  reg cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1;
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_8_itm_2;
  reg cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1;
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_7_itm_2;
  reg cvt_8_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_2;
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_6_itm_2;
  reg cvt_7_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_2;
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_5_itm_2;
  reg cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1;
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_4_itm_2;
  reg cvt_5_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_2;
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_3_itm_2;
  reg cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1;
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_2_itm_2;
  reg cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1;
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_1_itm_2;
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_1_itm_3;
  reg cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1;
  reg IntSaturation_17U_16U_IntSaturation_17U_16U_or_itm_2;
  reg cvt_1_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_itm_2;
  reg [1:0] cfg_proc_precision_1_sva_st_64;
  reg cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_st_2;
  reg cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_2;
  reg [1:0] cfg_proc_precision_1_sva_st_65;
  reg [1:0] cfg_proc_precision_1_sva_st_66;
  reg cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_st_2;
  reg cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2;
  reg cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_st_2;
  reg cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2;
  reg cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_st_2;
  reg cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  reg cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_st_2;
  reg cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2;
  reg [1:0] cfg_out_precision_1_sva_st_113;
  reg cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_st_2;
  reg cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  reg cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_st_2;
  reg cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  reg cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_st_2;
  reg cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2;
  reg cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_st_2;
  reg cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2;
  reg cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_st_2;
  reg cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  reg cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_st_2;
  reg cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  reg cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_st_2;
  reg cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2;
  reg cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_st_2;
  reg cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2;
  reg cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_st_2;
  reg cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2;
  reg cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_st_2;
  reg cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2;
  reg cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_4_svs_st_2;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_2;
  reg cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_st_2;
  reg cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_svs_st_2;
  reg [1:0] cfg_out_precision_1_sva_st_136;
  reg cvt_1_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_svs_st_2;
  reg cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2;
  reg cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  reg cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2;
  reg cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  reg cvt_3_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2;
  reg cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2;
  reg cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2;
  reg cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  reg cvt_5_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2;
  reg cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2;
  reg cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2;
  reg cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_svs_st_2;
  reg [1:0] cfg_proc_precision_1_sva_st_89;
  reg [1:0] cfg_proc_precision_1_sva_st_90;
  reg cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  reg [1:0] cfg_out_precision_1_sva_st_144;
  reg cvt_9_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2;
  reg [1:0] cfg_proc_precision_1_sva_st_101;
  reg [1:0] cfg_proc_precision_1_sva_st_102;
  reg [1:0] cfg_out_precision_1_sva_st_149;
  reg [1:0] cfg_proc_precision_1_sva_st_108;
  reg [1:0] cfg_out_precision_1_sva_st_154;
  reg [1:0] cfg_out_precision_1_sva_st_156;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_9_4_1;
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_9_3_0_1;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_9_4_1;
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_9_3_0_1;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_9_4_1;
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_9_3_0_1;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_9_4_1;
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_9_3_0_1;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_9_4_1;
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_9_3_0_1;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_9_4_1;
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_9_3_0_1;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_9_4_1;
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_9_3_0_1;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_9_4_1;
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_9_3_0_1;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_9_4_1;
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_9_3_0_1;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_9_4_1;
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_9_3_0_1;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_9_4_1;
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_9_3_0_1;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_9_4_1;
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_9_3_0_1;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_9_4_1;
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_9_3_0_1;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_9_4_1;
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_9_3_0_1;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_9_4_1;
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_9_3_0_1;
  reg FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_9_4_1;
  reg [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_9_3_0_1;
  reg chn_idata_data_sva_1_511_1;
  reg [28:0] chn_idata_data_sva_1_507_479_1;
  reg [28:0] chn_idata_data_sva_1_475_447_1;
  reg [28:0] chn_idata_data_sva_1_443_415_1;
  reg [28:0] chn_idata_data_sva_1_411_383_1;
  reg [28:0] chn_idata_data_sva_1_379_351_1;
  reg [28:0] chn_idata_data_sva_1_347_319_1;
  reg [28:0] chn_idata_data_sva_1_315_287_1;
  reg [28:0] chn_idata_data_sva_1_283_255_1;
  reg [28:0] chn_idata_data_sva_1_251_223_1;
  reg [28:0] chn_idata_data_sva_1_219_191_1;
  reg [28:0] chn_idata_data_sva_1_187_159_1;
  reg [28:0] chn_idata_data_sva_1_155_127_1;
  reg [28:0] chn_idata_data_sva_1_123_95_1;
  reg [28:0] chn_idata_data_sva_1_91_63_1;
  reg [28:0] chn_idata_data_sva_1_59_31_1;
  reg [27:0] chn_idata_data_sva_1_27_0_1;
  reg chn_idata_data_sva_2_511_1;
  reg [16:0] chn_idata_data_sva_2_495_479_1;
  reg [16:0] chn_idata_data_sva_2_463_447_1;
  reg [16:0] chn_idata_data_sva_2_431_415_1;
  reg [16:0] chn_idata_data_sva_2_399_383_1;
  reg [16:0] chn_idata_data_sva_2_367_351_1;
  reg [16:0] chn_idata_data_sva_2_335_319_1;
  reg [16:0] chn_idata_data_sva_2_303_287_1;
  reg [16:0] chn_idata_data_sva_2_271_255_1;
  reg [16:0] chn_idata_data_sva_2_239_223_1;
  reg [16:0] chn_idata_data_sva_2_207_191_1;
  reg [16:0] chn_idata_data_sva_2_175_159_1;
  reg [16:0] chn_idata_data_sva_2_143_127_1;
  reg [16:0] chn_idata_data_sva_2_111_95_1;
  reg [16:0] chn_idata_data_sva_2_79_63_1;
  reg [16:0] chn_idata_data_sva_2_47_31_1;
  reg [15:0] chn_idata_data_sva_2_15_0_1;
  reg [16:0] chn_idata_data_sva_3_495_479_1;
  reg [16:0] chn_idata_data_sva_3_463_447_1;
  reg [16:0] chn_idata_data_sva_3_431_415_1;
  reg [16:0] chn_idata_data_sva_3_399_383_1;
  reg [16:0] chn_idata_data_sva_3_367_351_1;
  reg [16:0] chn_idata_data_sva_3_335_319_1;
  reg [16:0] chn_idata_data_sva_3_303_287_1;
  reg [16:0] chn_idata_data_sva_3_271_255_1;
  reg [16:0] chn_idata_data_sva_3_239_223_1;
  reg [16:0] chn_idata_data_sva_3_207_191_1;
  reg [16:0] chn_idata_data_sva_3_175_159_1;
  reg [16:0] chn_idata_data_sva_3_143_127_1;
  reg [16:0] chn_idata_data_sva_3_111_95_1;
  reg [16:0] chn_idata_data_sva_3_79_63_1;
  reg [16:0] chn_idata_data_sva_3_47_31_1;
  wire main_stage_en_1;
  wire cvt_else_equal_tmp_4_mx1;
  wire cvt_else_equal_tmp_3_mx0;
  wire cvt_else_nor_dfs_1_mx1;
  wire cvt_else_equal_tmp_10_mx0;
  wire cvt_else_equal_tmp_9_mx1;
  wire cvt_else_nor_dfs_3_mx1;
  wire cvt_else_equal_tmp_46_mx1;
  wire cvt_else_equal_tmp_45_mx1;
  wire cvt_else_nor_dfs_15_mx1;
  wire cvt_else_equal_tmp_43_mx0;
  wire cvt_else_equal_tmp_42_mx0;
  wire cvt_else_nor_dfs_14_mx1;
  wire cvt_else_equal_tmp_16_mx1;
  wire cvt_else_equal_tmp_15_mx0;
  wire cvt_else_nor_dfs_5_mx1;
  wire cvt_else_equal_tmp_40_mx1;
  wire cvt_else_equal_tmp_39_mx1;
  wire cvt_else_nor_dfs_13_mx1;
  wire cvt_else_equal_tmp_19_mx0;
  wire cvt_else_equal_tmp_18_mx0;
  wire cvt_else_nor_dfs_6_mx1;
  wire cvt_else_equal_tmp_37_mx0;
  wire cvt_else_equal_tmp_36_mx0;
  wire cvt_else_equal_tmp_22_mx1;
  wire cvt_and_147_m1c;
  wire cvt_else_equal_tmp_21_mx1;
  wire cvt_else_nor_dfs_7_mx1;
  wire cvt_else_equal_tmp_34_mx1;
  wire cvt_else_equal_tmp_33_mx1;
  wire cvt_else_nor_dfs_11_mx1;
  wire cvt_else_equal_tmp_1;
  wire cvt_else_equal_tmp;
  wire cvt_else_nor_dfs;
  wire cvt_else_equal_tmp_31_mx0;
  wire cvt_else_equal_tmp_30_mx0;
  wire cvt_else_nor_dfs_10_mx1;
  wire cvt_else_equal_tmp_28_mx1;
  wire cvt_else_equal_tmp_27_mx0;
  wire cvt_else_nor_dfs_9_mx1;
  wire cvt_if_unequal_tmp;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_15_tmp;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_14_tmp;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_13_tmp;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_12_tmp;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_11_tmp;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_10_tmp;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_9_tmp;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_8_tmp;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_7_tmp;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_6_tmp;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_5_tmp;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_4_tmp;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_3_tmp;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_2_tmp;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_1_tmp;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_tmp;
  wire IsNaN_5U_10U_land_15_lpi_1_dfm_mx0w0;
  wire IsNaN_5U_10U_land_2_lpi_1_dfm_mx0w0;
  wire IsNaN_5U_10U_land_1_lpi_1_dfm_mx0w0;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_7_4_mx0w0;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_15_ssc;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_lpi_1_dfm;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_31_m1c;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_7_4_mx0w0;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_14_ssc;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_15_lpi_1_dfm;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_29_m1c;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_7_4_mx0w0;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_13_ssc;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_14_lpi_1_dfm;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_27_m1c;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_7_4_mx0w0;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_12_ssc;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_13_lpi_1_dfm;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_25_m1c;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_7_4_mx0w0;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_11_ssc;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_12_lpi_1_dfm;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_23_m1c;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_7_4_mx0w0;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_10_ssc;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_11_lpi_1_dfm;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_21_m1c;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_7_4_mx0w0;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_9_ssc;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_10_lpi_1_dfm;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_19_m1c;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_7_4_mx0w0;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_8_ssc;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_9_lpi_1_dfm;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_17_m1c;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_7_4_mx0w0;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_7_ssc;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_8_lpi_1_dfm;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_15_m1c;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_7_4_mx0w0;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_6_ssc;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_7_lpi_1_dfm;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_13_m1c;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_7_4_mx0w0;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_5_ssc;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_6_lpi_1_dfm;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_11_m1c;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_7_4_mx0w0;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_4_ssc;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_5_lpi_1_dfm;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_9_m1c;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_7_4_mx0w0;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_3_ssc;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_4_lpi_1_dfm;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_7_m1c;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_7_4_mx0w0;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_2_ssc;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_3_lpi_1_dfm;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_5_m1c;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_7_4_mx0w0;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_1_ssc;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_2_lpi_1_dfm;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_3_m1c;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_7_4_mx0w0;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_ssc;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_1_lpi_1_dfm;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_and_1_m1c;
  wire IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0;
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva;
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva;
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva;
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva;
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva;
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva;
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva;
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva;
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva;
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva;
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva;
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva;
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva;
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva;
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva;
  wire [74:0] IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_lpi_1_dfm_5_mx0;
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_7_3_0_mx0w0;
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva;
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva;
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_7_3_0_mx0w0;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_15_lpi_1_dfm_5_mx0;
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_15_sva;
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_15_sva;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_14_lpi_1_dfm_5_mx0;
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_7_3_0_mx0w0;
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_14_sva;
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_14_sva;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_13_lpi_1_dfm_5_mx0;
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_7_3_0_mx0w0;
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_13_sva;
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_13_sva;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_12_lpi_1_dfm_5_mx0;
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_7_3_0_mx0w0;
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_12_sva;
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_12_sva;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_11_lpi_1_dfm_5_mx0;
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_7_3_0_mx0w0;
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_11_sva;
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_11_sva;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_10_lpi_1_dfm_5_mx0;
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_7_3_0_mx0w0;
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_10_sva;
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_10_sva;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_9_lpi_1_dfm_5_mx0;
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_7_3_0_mx0w0;
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_9_sva;
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_9_sva;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_8_lpi_1_dfm_5_mx0;
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_7_3_0_mx0w0;
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_8_sva;
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_8_sva;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_7_lpi_1_dfm_5_mx0;
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_7_3_0_mx0w0;
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_7_sva;
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_7_sva;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_6_lpi_1_dfm_5_mx0;
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_7_3_0_mx0w0;
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_6_sva;
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_6_sva;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_5_lpi_1_dfm_5_mx0;
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_7_3_0_mx0w0;
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_5_sva;
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_5_sva;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_4_lpi_1_dfm_5_mx0;
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_7_3_0_mx0w0;
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_4_sva;
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_4_sva;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_3_lpi_1_dfm_5_mx0;
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_7_3_0_mx0w0;
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_3_sva;
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_3_sva;
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_7_3_0_mx0w0;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_2_lpi_1_dfm_5_mx0;
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_2_sva;
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_2_sva;
  wire [3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_7_3_0_mx0w0;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_1_lpi_1_dfm_5_mx0;
  wire [10:0] FpMantDecShiftRight_23U_8U_10U_o_mant_sum_1_sva;
  wire [11:0] nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_1_sva;
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_sva_mx0w0;
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_mx0w0;
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_mx0w0;
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_mx0w0;
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_mx0w0;
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_mx0w0;
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_mx0w0;
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_mx0w0;
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_mx0w0;
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_mx0w0;
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_mx0w0;
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_mx0w0;
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_mx0w0;
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_mx0w0;
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_mx0w0;
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_mx0w0;
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_sva;
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_sva;
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_15_sva;
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_15_sva;
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_14_sva;
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_14_sva;
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_13_sva;
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_13_sva;
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_12_sva;
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_12_sva;
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_11_sva;
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_11_sva;
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_10_sva;
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_10_sva;
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_9_sva;
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_9_sva;
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_8_sva;
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_8_sva;
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_7_sva;
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_7_sva;
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_6_sva;
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_6_sva;
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_5_sva;
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_5_sva;
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_4_sva;
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_4_sva;
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_3_sva;
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_3_sva;
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_2_sva;
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_2_sva;
  wire [44:0] IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_1_sva;
  wire [45:0] nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_1_sva;
  wire and_1176_m1c;
  wire and_1172_m1c;
  wire and_1159_m1c;
  wire and_1155_m1c;
  wire and_1145_m1c;
  wire and_1141_m1c;
  wire and_1132_m1c;
  wire and_1123_m1c;
  wire and_1119_m1c;
  wire and_1115_m1c;
  wire and_1106_m1c;
  wire and_1097_m1c;
  wire and_1093_m1c;
  wire and_1084_m1c;
  wire and_1080_m1c;
  wire and_1069_m1c;
  wire cvt_or_cse;
  wire chn_out_and_cse;
  wire cvt_or_2_cse;
  wire cvt_or_6_cse;
  wire cvt_or_10_cse;
  wire cvt_or_12_cse;
  wire cvt_or_14_cse;
  wire cvt_or_18_cse;
  wire cvt_or_20_cse;
  wire cvt_or_22_cse;
  wire cvt_or_24_cse;
  wire cvt_or_26_cse;
  wire cvt_or_28_cse;
  wire cvt_or_30_cse;
  wire chn_out_and_32_cse;
  wire chn_out_and_77_cse;
  wire nor_2040_cse;
  wire nor_50_cse;
  wire or_419_cse;
  wire or_423_cse;
  wire or_451_cse;
  wire or_513_cse;
  wire or_4535_cse;
  wire nand_219_cse;
  wire nor_1056_cse;
  wire nor_1672_cse;
  wire FpFloatToInt_16U_5U_10U_internal_int_and_cse;
  wire nor_1664_cse;
  wire or_1176_cse;
  wire or_1157_cse;
  wire IsNaN_5U_10U_aelse_and_1_cse;
  wire nor_1666_cse;
  wire or_300_cse;
  wire nor_1669_cse;
  wire or_1159_cse;
  wire nor_1624_cse;
  wire nor_1630_cse;
  wire or_309_cse;
  wire IsNaN_5U_10U_aelse_and_cse;
  wire or_1196_cse;
  wire nor_151_cse;
  wire nor_1629_cse;
  wire IntShiftRightSat_49U_6U_17U_o_and_cse;
  wire cvt_else_and_cse;
  wire cvt_else_and_10_cse;
  wire cvt_else_and_19_cse;
  wire or_1202_cse;
  wire or_425_cse;
  wire nor_63_cse;
  wire or_1587_cse;
  wire nor_183_cse;
  wire and_2186_cse;
  wire FpIntToFloat_17U_5U_10U_is_inf_and_8_cse;
  wire nor_1589_cse;
  wire FpIntToFloat_17U_5U_10U_is_inf_and_10_cse;
  reg reg_chn_out_rsci_ld_core_psct_cse;
  wire nor_8_cse;
  wire or_4524_cse;
  wire or_2289_cse;
  wire nand_190_cse;
  wire nand_164_cse;
  wire nand_162_cse;
  wire nand_160_cse;
  wire nand_158_cse;
  wire nand_156_cse;
  wire nand_153_cse;
  wire nand_151_cse;
  wire nand_149_cse;
  wire nand_147_cse;
  wire nand_145_cse;
  wire nand_143_cse;
  wire nand_141_cse;
  wire nand_139_cse;
  wire nand_137_cse;
  wire nand_135_cse;
  wire nand_133_cse;
  wire and_2239_cse;
  wire nor_1185_cse;
  wire nor_1186_cse;
  wire or_1596_cse;
  wire or_1625_cse;
  wire or_1693_cse;
  wire or_1829_cse;
  wire nor_1099_cse;
  wire and_2237_cse;
  wire nor_57_cse;
  wire or_510_cse;
  wire and_2230_cse;
  wire or_600_cse;
  wire or_4536_cse;
  wire and_2206_cse;
  wire and_2199_cse;
  wire and_2194_cse;
  wire nor_1626_cse;
  wire or_3538_cse;
  wire or_3542_cse;
  wire nor_1556_cse;
  wire or_1919_cse;
  wire cvt_cvt_nand_cse;
  wire cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_nor_4_cse;
  wire cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse;
  wire cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse;
  wire cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse;
  wire cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse;
  wire cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse;
  wire cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse;
  wire cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse;
  wire cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse;
  wire cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse;
  wire cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse;
  wire cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse;
  wire cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse;
  wire cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse;
  wire cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse;
  wire cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_nor_24_cse;
  wire or_578_cse;
  wire nor_45_cse;
  wire or_tmp_3763;
  wire [14:0] FpIntToFloat_17U_5U_10U_else_if_mux1h_9_rgt;
  wire or_tmp_3768;
  wire [14:0] FpIntToFloat_17U_5U_10U_else_if_mux1h_12_rgt;
  wire [14:0] FpIntToFloat_17U_5U_10U_else_if_mux1h_15_rgt;
  wire [14:0] FpIntToFloat_17U_5U_10U_else_if_mux1h_18_rgt;
  wire [14:0] FpIntToFloat_17U_5U_10U_else_if_mux1h_21_rgt;
  wire [14:0] FpIntToFloat_17U_5U_10U_else_if_mux1h_27_rgt;
  wire [14:0] FpIntToFloat_17U_5U_10U_else_if_mux1h_30_rgt;
  wire [14:0] FpIntToFloat_17U_5U_10U_else_if_mux1h_33_rgt;
  wire [14:0] FpIntToFloat_17U_5U_10U_else_if_mux1h_36_rgt;
  wire or_tmp_3826;
  wire mux_tmp_2203;
  wire or_tmp_3832;
  wire mux_tmp_2206;
  wire [14:0] FpIntToFloat_17U_5U_10U_else_i_abs_mux1h_17_rgt;
  wire or_tmp_3840;
  wire [14:0] FpIntToFloat_17U_5U_10U_else_if_mux1h_41_rgt;
  wire or_tmp_3849;
  wire [14:0] FpIntToFloat_17U_5U_10U_else_if_mux1h_44_rgt;
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_1_rgt;
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_2_rgt;
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_4_rgt;
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_5_rgt;
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_6_rgt;
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_7_rgt;
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_8_rgt;
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_9_rgt;
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_10_rgt;
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_11_rgt;
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_12_rgt;
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_13_rgt;
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_14_rgt;
  wire [14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_15_rgt;
  wire [14:0] IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_mux_rgt;
  wire [15:0] chn_idata_data_mux1h_65_rgt;
  reg [4:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_4_lpi_1_dfm_6_reg;
  reg [9:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_4_lpi_1_dfm_6_1_reg;
  reg [4:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_5_lpi_1_dfm_5_reg;
  reg [9:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_5_lpi_1_dfm_5_1_reg;
  reg [4:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_6_lpi_1_dfm_6_reg;
  reg [9:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_6_lpi_1_dfm_6_1_reg;
  reg [4:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_7_lpi_1_dfm_6_reg;
  reg [9:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_7_lpi_1_dfm_6_1_reg;
  reg [4:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_8_lpi_1_dfm_7_reg;
  reg [9:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_8_lpi_1_dfm_7_1_reg;
  reg [4:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_10_lpi_1_dfm_6_reg;
  reg [9:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_10_lpi_1_dfm_6_1_reg;
  reg [4:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_11_lpi_1_dfm_6_reg;
  reg [9:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_11_lpi_1_dfm_6_1_reg;
  reg [4:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_12_lpi_1_dfm_7_reg;
  reg [9:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_12_lpi_1_dfm_7_1_reg;
  reg [4:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_13_lpi_1_dfm_6_reg;
  reg [9:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_13_lpi_1_dfm_6_1_reg;
  reg [4:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_14_lpi_1_dfm_7_reg;
  reg [9:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_14_lpi_1_dfm_7_1_reg;
  reg [4:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_15_lpi_1_dfm_7_reg;
  reg [9:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_15_lpi_1_dfm_7_1_reg;
  reg [4:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_lpi_1_dfm_8_reg;
  reg [9:0] reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_lpi_1_dfm_8_1_reg;
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_reg;
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_1_reg;
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_reg;
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_1_reg;
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_reg;
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_1_reg;
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_reg;
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_1_reg;
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_reg;
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_1_reg;
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_reg;
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_1_reg;
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_reg;
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_1_reg;
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_reg;
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_1_reg;
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_reg;
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_1_reg;
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_reg;
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_1_reg;
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_reg;
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_1_reg;
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_reg;
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_1_reg;
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_reg;
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_1_reg;
  reg [4:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_reg;
  reg [9:0] reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_1_reg;
  reg [4:0] reg_IntShiftRightSat_49U_6U_17U_o_15_1_14_1_reg;
  reg [9:0] reg_IntShiftRightSat_49U_6U_17U_o_15_1_14_3_reg;
  reg reg_chn_idata_data_sva_3_15_0_reg;
  reg [4:0] reg_chn_idata_data_sva_3_15_0_1_reg;
  reg [9:0] reg_chn_idata_data_sva_3_15_0_2_reg;
  wire mux_813_cse;
  wire nand_207_cse;
  wire mux_827_cse;
  wire nor_2099_cse;
  wire mux_1436_cse;
  wire mux_1126_cse;
  wire mux_1464_cse;
  wire nor_1320_cse;
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_10_itm_mx0w0;
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_13_itm_mx0w0;
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_16_itm_mx0w0;
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_19_itm_mx0w0;
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_22_itm_mx0w0;
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_28_itm_mx0w0;
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_31_itm_mx0w0;
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_34_itm_mx0w0;
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_37_itm_mx0w0;
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_40_itm_mx0w0;
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_43_itm_mx0w0;
  wire [9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_46_itm_mx0w0;
  wire [16:0] FpIntToFloat_17U_5U_10U_else_int_mant_2_sva;
  wire FpMantRNE_17U_11U_else_carry_2_sva;
  wire [16:0] FpIntToFloat_17U_5U_10U_else_int_mant_9_sva;
  wire FpMantRNE_17U_11U_else_carry_9_sva;
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_1_sva;
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_1_sva;
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_1_sva;
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_1_lpi_1_dfm_mx0;
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_m1c;
  wire [16:0] FpIntToFloat_17U_5U_10U_else_int_mant_1_sva;
  wire FpMantRNE_17U_11U_else_carry_1_sva;
  wire or_4550_cse;
  wire and_2360_cse;
  wire or_4709_cse;
  wire nor_2285_cse;
  wire mux_2230_cse;
  wire or_4714_cse;
  wire nor_2219_cse;
  wire mux_344_cse;
  wire mux_474_cse;
  wire and_1386_cse;
  wire and_1078_cse;
  wire mux_1494_cse;
  wire mux_660_cse;
  wire mux_201_cse;
  wire mux_1142_cse;
  wire and_550_cse;
  wire and_2365_cse;
  wire and_2369_cse;
  wire nand_202_cse;
  wire mux_767_cse;
  wire or_4749_cse;
  wire or_4788_cse;
  wire and_2388_cse;
  wire and_2422_cse;
  wire and_637_rgt;
  wire and_639_rgt;
  wire and_641_rgt;
  wire and_643_rgt;
  wire and_646_rgt;
  wire and_648_rgt;
  wire and_650_rgt;
  wire and_652_rgt;
  wire and_654_rgt;
  wire and_656_rgt;
  wire and_658_rgt;
  wire and_660_rgt;
  wire and_662_rgt;
  wire and_664_rgt;
  wire and_666_rgt;
  wire and_668_rgt;
  wire and_685_rgt;
  wire and_704_rgt;
  wire and_719_rgt;
  wire and_734_rgt;
  wire and_749_rgt;
  wire and_766_rgt;
  wire and_787_rgt;
  wire and_801_rgt;
  wire and_816_rgt;
  wire and_830_rgt;
  wire and_849_rgt;
  wire and_866_rgt;
  wire and_881_rgt;
  wire and_896_rgt;
  wire and_900_rgt;
  wire and_954_rgt;
  wire and_956_rgt;
  wire and_957_rgt;
  wire and_984_rgt;
  wire and_986_rgt;
  wire and_987_rgt;
  wire and_989_rgt;
  wire and_1009_rgt;
  wire and_1011_rgt;
  wire and_1077_rgt;
  wire [16:0] cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp;
  wire and_1091_rgt;
  wire [16:0] cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp;
  wire and_dcpl_1319;
  wire [16:0] cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp;
  wire and_1104_rgt;
  wire [16:0] cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp;
  wire [16:0] cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp;
  wire [16:0] cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp;
  wire [16:0] cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp;
  wire [16:0] cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp;
  wire [16:0] cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp;
  wire [16:0] cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp;
  wire [16:0] cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp;
  wire [16:0] cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp;
  wire [16:0] cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_tmp;
  wire and_1213_rgt;
  wire and_1247_rgt;
  wire and_1250_rgt;
  wire and_1321_rgt;
  wire and_1325_rgt;
  wire and_1329_rgt;
  wire and_1333_rgt;
  wire and_1337_rgt;
  wire and_1341_rgt;
  wire and_1345_rgt;
  wire and_1349_rgt;
  wire and_1353_rgt;
  wire and_1357_rgt;
  wire and_1361_rgt;
  wire and_1365_rgt;
  wire and_1369_rgt;
  wire and_1373_rgt;
  wire and_1377_rgt;
  wire and_1381_rgt;
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_rgt;
  wire IntSaturation_17U_16U_and_31_rgt;
  wire IntSaturation_17U_16U_o_and_31_rgt;
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_1_rgt;
  wire IntSaturation_17U_16U_and_29_rgt;
  wire IntSaturation_17U_16U_o_and_29_rgt;
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_2_rgt;
  wire IntSaturation_17U_16U_and_27_rgt;
  wire IntSaturation_17U_16U_o_and_27_rgt;
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_3_rgt;
  wire IntSaturation_17U_16U_and_25_rgt;
  wire IntSaturation_17U_16U_o_and_25_rgt;
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_4_rgt;
  wire IntSaturation_17U_16U_and_23_rgt;
  wire IntSaturation_17U_16U_o_and_23_rgt;
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_5_rgt;
  wire IntSaturation_17U_16U_and_21_rgt;
  wire IntSaturation_17U_16U_o_and_21_rgt;
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_6_rgt;
  wire IntSaturation_17U_16U_and_19_rgt;
  wire IntSaturation_17U_16U_o_and_19_rgt;
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_7_rgt;
  wire IntSaturation_17U_16U_and_17_rgt;
  wire IntSaturation_17U_16U_o_and_17_rgt;
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_8_rgt;
  wire IntSaturation_17U_16U_and_15_rgt;
  wire IntSaturation_17U_16U_o_and_15_rgt;
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_9_rgt;
  wire IntSaturation_17U_16U_and_13_rgt;
  wire IntSaturation_17U_16U_o_and_13_rgt;
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_10_rgt;
  wire IntSaturation_17U_16U_and_11_rgt;
  wire IntSaturation_17U_16U_o_and_11_rgt;
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_11_rgt;
  wire IntSaturation_17U_16U_and_9_rgt;
  wire IntSaturation_17U_16U_o_and_9_rgt;
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_12_rgt;
  wire IntSaturation_17U_16U_and_7_rgt;
  wire IntSaturation_17U_16U_o_and_7_rgt;
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_13_rgt;
  wire IntSaturation_17U_16U_and_5_rgt;
  wire IntSaturation_17U_16U_o_and_5_rgt;
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_14_rgt;
  wire IntSaturation_17U_16U_and_3_rgt;
  wire IntSaturation_17U_16U_o_and_3_rgt;
  wire IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_15_rgt;
  wire IntSaturation_17U_16U_and_1_rgt;
  wire IntSaturation_17U_16U_o_and_1_rgt;
  wire and_1385_rgt;
  wire and_1467_rgt;
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_1_itm;
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_1_lpi_1_dfm_7_itm;
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_1_lpi_1_dfm_7_1_itm;
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_3_itm;
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_2_lpi_1_dfm_8_itm;
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_2_lpi_1_dfm_8_1_itm;
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_5_itm;
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_3_lpi_1_dfm_8_itm;
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_3_lpi_1_dfm_8_1_itm;
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_7_itm;
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_4_lpi_1_dfm_9_itm;
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_4_lpi_1_dfm_9_1_itm;
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_9_itm;
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_5_lpi_1_dfm_8_itm;
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_5_lpi_1_dfm_8_1_itm;
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_11_itm;
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_6_lpi_1_dfm_9_itm;
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_6_lpi_1_dfm_9_1_itm;
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_13_itm;
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_7_lpi_1_dfm_9_itm;
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_7_lpi_1_dfm_9_1_itm;
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_15_itm;
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_8_lpi_1_dfm_10_itm;
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_8_lpi_1_dfm_10_1_itm;
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_17_itm;
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_9_lpi_1_dfm_8_itm;
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_9_lpi_1_dfm_8_1_itm;
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_19_itm;
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_10_lpi_1_dfm_9_itm;
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_10_lpi_1_dfm_9_1_itm;
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_21_itm;
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_11_lpi_1_dfm_9_itm;
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_11_lpi_1_dfm_9_1_itm;
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_23_itm;
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_12_lpi_1_dfm_10_itm;
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_12_lpi_1_dfm_10_1_itm;
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_25_itm;
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_13_lpi_1_dfm_9_itm;
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_13_lpi_1_dfm_9_1_itm;
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_27_itm;
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_14_lpi_1_dfm_10_itm;
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_14_lpi_1_dfm_10_1_itm;
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_29_itm;
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_15_lpi_1_dfm_10_itm;
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_15_lpi_1_dfm_10_1_itm;
  wire [4:0] FpIntToFloat_17U_5U_10U_o_expo_mux1h_31_itm;
  reg reg_FpIntToFloat_17U_5U_10U_o_expo_lpi_1_dfm_11_itm;
  reg [3:0] reg_FpIntToFloat_17U_5U_10U_o_expo_lpi_1_dfm_11_1_itm;
  wire [23:0] cvt_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_itm;
  wire [23:0] cvt_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_itm;
  wire [23:0] cvt_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_itm;
  wire [23:0] cvt_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm;
  wire [23:0] cvt_5_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_itm;
  wire [23:0] cvt_6_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm;
  wire [23:0] cvt_7_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm;
  wire [23:0] cvt_8_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_itm;
  wire [23:0] cvt_9_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_itm;
  wire [23:0] cvt_10_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm;
  wire [23:0] cvt_11_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm;
  wire [23:0] cvt_12_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_itm;
  wire [23:0] cvt_13_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm;
  wire [23:0] cvt_14_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_itm;
  wire [23:0] cvt_15_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_itm;
  wire [23:0] cvt_16_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_4_itm;
  wire mux_1966_itm;
  wire cvt_and_tmp_1;
  wire chn_in_rsci_ld_core_psct_mx0c0;
  wire cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
  wire cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
  wire cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_sig_mx0w1;
  wire cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1_sig_mx0w1;
  wire main_stage_v_1_mx0c1;
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_2_sva_mx0w0;
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_2_sva_mx0w0;
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_3_sva_mx0w0;
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_3_sva_mx0w0;
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_4_sva_mx0w0;
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_4_sva_mx0w0;
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_5_sva_mx0w0;
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_5_sva_mx0w0;
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_6_sva_mx0w0;
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_6_sva_mx0w0;
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_7_sva_mx0w0;
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_7_sva_mx0w0;
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_8_sva_mx0w0;
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_8_sva_mx0w0;
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_9_sva_mx0w0;
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_9_sva_mx0w0;
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_10_sva_mx0w0;
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_10_sva_mx0w0;
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_11_sva_mx0w0;
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_11_sva_mx0w0;
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_12_sva_mx0w0;
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_12_sva_mx0w0;
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_13_sva_mx0w0;
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_13_sva_mx0w0;
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_14_sva_mx0w0;
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_14_sva_mx0w0;
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_15_sva_mx0w0;
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_15_sva_mx0w0;
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_16_sva_mx0w0;
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_16_sva_mx0w0;
  wire [2:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_mx0w0;
  wire [3:0] nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_mx0w0;
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_4_sva_mx0w1;
  wire IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1;
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_6_sva_mx0w1;
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_8_sva_mx0w1;
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_7_sva_mx0w1;
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_10_sva_mx0w1;
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_12_sva_mx0w1;
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_11_sva_mx0w1;
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_14_sva_mx0w1;
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_sva_mx0w1;
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_15_sva_mx0w1;
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_13_sva_mx0w1;
  wire main_stage_v_2_mx0c1;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_mx0w1;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_1_mx0w1;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_2_mx0w1;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_3_mx0w1;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_4_mx0w1;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_5_mx0w1;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_6_mx0w1;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_7_mx0w1;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_8_mx0w1;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_9_mx0w1;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_10_mx0w1;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_11_mx0w1;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_12_mx0w1;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_13_mx0w1;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_14_mx0w1;
  wire [9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_15_mx0w1;
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_1_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_0_1_sva_mx0w0;
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_2_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_0_2_sva_mx0w0;
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_3_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_0_3_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_0_4_sva_mx0w0;
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_5_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_0_5_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_0_6_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_0_7_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_0_8_sva_mx0w0;
  wire [48:0] IntShiftRightSat_49U_6U_17U_i_9_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_0_9_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_0_10_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_0_11_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_0_12_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_0_13_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_0_14_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_0_15_sva_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_o_0_sva_mx0w0;
  wire main_stage_v_3_mx0c1;
  wire FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_mx0w0;
  wire FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_mx0w0;
  wire cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c0;
  wire cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c1;
  wire FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_mx0w0;
  wire cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c0;
  wire cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c1;
  wire FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_mx0w0;
  wire cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0;
  wire cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1;
  wire FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c1;
  wire FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c2;
  wire FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_mx0w0;
  wire FpFloatToInt_16U_5U_10U_internal_int_0_sva_mx0w0;
  wire cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1_mx0c0;
  wire cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1_mx0c1;
  wire FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_mx0w0;
  wire cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0;
  wire cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1;
  wire FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_mx0w0;
  wire FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_mx0w0;
  wire FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_mx0w0;
  wire cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c0;
  wire cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c1;
  wire FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_mx0w0;
  wire FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_mx0w0;
  wire cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0;
  wire cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1;
  wire FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_mx0w0;
  wire cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c0;
  wire cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c1;
  wire FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_mx0w0;
  wire cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c0;
  wire cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c1;
  wire FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_mx0w0;
  wire cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0;
  wire cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1;
  wire FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_mx0w0;
  wire cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0;
  wire cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1;
  wire chn_odata_data_13_0_lpi_1_dfm_1_mx0w0;
  wire FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_2_mx1w0;
  wire FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_2_mx1w0;
  wire FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_2_mx1w0;
  wire FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_2_mx1w0;
  wire FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_2_mx0w0;
  wire FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_2_mx1w0;
  wire FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_2_mx1w0;
  wire FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_2_mx0w0;
  wire FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2_mx0w0;
  wire FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_2_mx0w0;
  wire FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_2_mx0w0;
  wire FpMantRNE_24U_11U_else_carry_1_sva_mx0w0;
  wire FpMantRNE_24U_11U_else_carry_2_sva_mx0w0;
  wire FpMantRNE_24U_11U_else_carry_3_sva_mx0w0;
  wire FpMantRNE_24U_11U_else_carry_4_sva_mx0w0;
  wire FpMantRNE_24U_11U_else_carry_5_sva_mx0w0;
  wire FpMantRNE_24U_11U_else_carry_6_sva_mx0w0;
  wire FpMantRNE_24U_11U_else_carry_7_sva_mx0w0;
  wire FpMantRNE_24U_11U_else_carry_8_sva_mx0w0;
  wire FpMantRNE_24U_11U_else_carry_9_sva_mx0w0;
  wire FpMantRNE_24U_11U_else_carry_10_sva_mx0w0;
  wire FpMantRNE_24U_11U_else_carry_11_sva_mx0w0;
  wire FpMantRNE_24U_11U_else_carry_12_sva_mx0w0;
  wire FpMantRNE_24U_11U_else_carry_13_sva_mx0w0;
  wire FpMantRNE_24U_11U_else_carry_14_sva_mx0w0;
  wire FpMantRNE_24U_11U_else_carry_15_sva_mx0w0;
  wire FpMantRNE_24U_11U_else_carry_sva_mx0w0;
  wire IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm_mx0w0;
  wire IntShiftRightSat_49U_6U_17U_lor_3_lpi_1_dfm_mx1w0;
  wire IntShiftRightSat_49U_6U_17U_lor_5_lpi_1_dfm_mx1w0;
  wire IntShiftRightSat_49U_6U_17U_lor_4_lpi_1_dfm_mx1w0;
  wire IntShiftRightSat_49U_6U_17U_lor_7_lpi_1_dfm_mx1w0;
  wire IntShiftRightSat_49U_6U_17U_lor_9_lpi_1_dfm_mx1w0;
  wire IntShiftRightSat_49U_6U_17U_lor_8_lpi_1_dfm_mx1w0;
  wire IntShiftRightSat_49U_6U_17U_lor_6_lpi_1_dfm_mx1w0;
  wire IntShiftRightSat_49U_6U_17U_lor_11_lpi_1_dfm_mx1w0;
  wire IntShiftRightSat_49U_6U_17U_lor_13_lpi_1_dfm_mx1w0;
  wire IntShiftRightSat_49U_6U_17U_lor_12_lpi_1_dfm_mx1w0;
  wire IntShiftRightSat_49U_6U_17U_lor_15_lpi_1_dfm_mx1w0;
  wire IntShiftRightSat_49U_6U_17U_lor_lpi_1_dfm_mx1w0;
  wire IntShiftRightSat_49U_6U_17U_lor_16_lpi_1_dfm_mx1w0;
  wire IntShiftRightSat_49U_6U_17U_lor_14_lpi_1_dfm_mx1w0;
  wire IntShiftRightSat_49U_6U_17U_lor_10_lpi_1_dfm_mx1w0;
  wire IntShiftRightSat_49U_6U_17U_lor_2_lpi_1_dfm_mx1w0;
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva;
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva;
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva;
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva;
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva;
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva;
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva;
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva;
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva;
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva;
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva;
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva;
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva;
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva;
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva;
  wire [111:0] IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_1_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_1_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_2_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_2_sva;
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_2_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_3_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_3_sva;
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_3_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_4_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_4_sva;
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_4_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_5_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_5_sva;
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_5_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_6_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_6_sva;
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_6_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_7_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_7_sva;
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_7_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_8_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_8_sva;
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_8_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_9_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_9_sva;
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_9_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_10_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_10_sva;
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_10_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_11_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_11_sva;
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_11_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_12_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_12_sva;
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_12_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_13_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_13_sva;
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_13_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_14_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_14_sva;
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_14_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_15_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_15_sva;
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_15_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_sva;
  wire IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_sva;
  wire [23:0] FpFloatToInt_16U_5U_10U_internal_int_24_1_sva;
  wire FpMantRNE_17U_11U_else_carry_3_sva;
  wire FpMantRNE_17U_11U_else_carry_4_sva;
  wire FpMantRNE_17U_11U_else_carry_5_sva;
  wire FpMantRNE_17U_11U_else_carry_6_sva;
  wire FpMantRNE_17U_11U_else_carry_7_sva;
  wire FpMantRNE_17U_11U_else_carry_8_sva;
  wire FpMantRNE_17U_11U_else_carry_10_sva;
  wire FpMantRNE_17U_11U_else_carry_11_sva;
  wire FpMantRNE_17U_11U_else_carry_12_sva;
  wire FpMantRNE_17U_11U_else_carry_13_sva;
  wire FpMantRNE_17U_11U_else_carry_14_sva;
  wire FpMantRNE_17U_11U_else_carry_15_sva;
  wire FpMantRNE_17U_11U_else_carry_sva;
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_1_lpi_1_dfm_1;
  wire [6:0] IntSaturation_17U_8U_o_7_1_1_lpi_1_dfm_1;
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_2_lpi_1_dfm_1;
  wire [6:0] IntSaturation_17U_8U_o_7_1_2_lpi_1_dfm_1;
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_3_lpi_1_dfm_1;
  wire [6:0] IntSaturation_17U_8U_o_7_1_3_lpi_1_dfm_1;
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_4_lpi_1_dfm_1;
  wire [6:0] IntSaturation_17U_8U_o_7_1_4_lpi_1_dfm_1;
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_5_lpi_1_dfm_1;
  wire [6:0] IntSaturation_17U_8U_o_7_1_5_lpi_1_dfm_1;
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_6_lpi_1_dfm_1;
  wire [6:0] IntSaturation_17U_8U_o_7_1_6_lpi_1_dfm_1;
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_7_lpi_1_dfm_1;
  wire [6:0] IntSaturation_17U_8U_o_7_1_7_lpi_1_dfm_1;
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_8_lpi_1_dfm_1;
  wire [6:0] IntSaturation_17U_8U_o_7_1_8_lpi_1_dfm_1;
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_9_lpi_1_dfm_1;
  wire [6:0] IntSaturation_17U_8U_o_7_1_9_lpi_1_dfm_1;
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_10_lpi_1_dfm_1;
  wire [6:0] IntSaturation_17U_8U_o_7_1_10_lpi_1_dfm_1;
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_11_lpi_1_dfm_1;
  wire [6:0] IntSaturation_17U_8U_o_7_1_11_lpi_1_dfm_1;
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_12_lpi_1_dfm_1;
  wire [6:0] IntSaturation_17U_8U_o_7_1_12_lpi_1_dfm_1;
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_13_lpi_1_dfm_1;
  wire [6:0] IntSaturation_17U_8U_o_7_1_13_lpi_1_dfm_1;
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_14_lpi_1_dfm_1;
  wire [6:0] IntSaturation_17U_8U_o_7_1_14_lpi_1_dfm_1;
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_15_lpi_1_dfm_1;
  wire [6:0] IntSaturation_17U_8U_o_7_1_15_lpi_1_dfm_1;
  wire [9:0] FpIntToFloat_17U_5U_10U_o_mant_lpi_1_dfm_1;
  wire [6:0] IntSaturation_17U_8U_o_7_1_lpi_1_dfm_1;
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_2_lpi_1_dfm_mx0;
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_2_sva;
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_2_sva;
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_3_lpi_1_dfm_mx0;
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_3_sva;
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_3_sva;
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_4_lpi_1_dfm_mx0;
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_4_sva;
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_4_sva;
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_5_lpi_1_dfm_mx0;
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_5_sva;
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_5_sva;
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_6_lpi_1_dfm_mx0;
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_6_sva;
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_6_sva;
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_7_lpi_1_dfm_mx0;
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_7_sva;
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_7_sva;
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_8_lpi_1_dfm_mx0;
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_8_sva;
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_8_sva;
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_9_lpi_1_dfm_mx0;
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_9_sva;
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_9_sva;
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_10_lpi_1_dfm_mx0;
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_10_sva;
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_10_sva;
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_11_lpi_1_dfm_mx0;
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_11_sva;
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_11_sva;
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_12_lpi_1_dfm_mx0;
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_12_sva;
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_12_sva;
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_13_lpi_1_dfm_mx0;
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_13_sva;
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_13_sva;
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_14_lpi_1_dfm_mx0;
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_14_sva;
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_14_sva;
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_15_lpi_1_dfm_mx0;
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_15_sva;
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_15_sva;
  wire [15:0] FpFloatToInt_16U_5U_10U_if_qr_lpi_1_dfm_mx0;
  wire [15:0] FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_sva;
  wire [16:0] nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_1_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_1_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_1_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_1_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_1_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_2_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_2_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_2_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_2_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_2_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_3_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_3_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_3_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_3_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_3_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_4_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_4_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_4_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_4_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_4_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_5_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_5_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_5_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_5_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_5_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_6_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_6_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_6_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_6_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_6_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_7_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_7_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_7_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_7_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_7_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_8_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_8_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_8_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_8_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_8_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_9_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_9_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_9_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_9_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_9_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_10_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_10_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_10_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_10_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_10_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_11_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_11_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_11_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_11_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_11_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_12_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_12_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_12_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_12_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_12_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_13_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_13_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_13_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_13_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_13_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_14_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_14_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_14_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_14_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_14_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_15_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_15_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_15_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_15_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_15_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_guard_mask_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_sva;
  wire [22:0] FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_sva;
  wire [23:0] FpMantDecShiftRight_23U_8U_10U_least_mask_sva;
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_1_sva;
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_1_sva;
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_2_sva;
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_2_sva;
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_3_sva;
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_3_sva;
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_4_sva;
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_4_sva;
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_5_sva;
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_5_sva;
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_6_sva;
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_6_sva;
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_7_sva;
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_7_sva;
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_8_sva;
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_8_sva;
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_9_sva;
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_9_sva;
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_10_sva;
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_10_sva;
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_11_sva;
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_11_sva;
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_12_sva;
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_12_sva;
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_13_sva;
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_13_sva;
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_14_sva;
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_14_sva;
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_15_sva;
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_15_sva;
  wire [16:0] FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_sva;
  wire [17:0] nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_sva;
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_1_m1c;
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_2_m1c;
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_3_m1c;
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_4_m1c;
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_5_m1c;
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_6_m1c;
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_7_m1c;
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_8_m1c;
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_9_m1c;
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_10_m1c;
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_11_m1c;
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_12_m1c;
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_13_m1c;
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_14_m1c;
  wire FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_15_m1c;
  wire cvt_asn_319;
  wire cvt_asn_321;
  wire cvt_asn_323;
  wire cvt_asn_327;
  wire cvt_asn_329;
  wire cvt_asn_333;
  wire cvt_asn_335;
  wire cvt_asn_339;
  wire cvt_asn_341;
  wire cvt_asn_345;
  wire cvt_asn_347;
  wire cvt_asn_351;
  wire cvt_asn_353;
  wire cvt_asn_357;
  wire cvt_asn_359;
  wire cvt_asn_363;
  wire cvt_asn_365;
  wire cvt_asn_369;
  wire cvt_asn_371;
  wire cvt_asn_375;
  wire cvt_asn_377;
  wire cvt_asn_381;
  wire cvt_asn_383;
  wire cvt_asn_387;
  wire cvt_asn_389;
  wire cvt_asn_393;
  wire cvt_asn_399;
  wire cvt_1_FpIntToFloat_17U_5U_10U_else_i_abs_conc_3_16;
  wire cvt_2_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16;
  wire cvt_3_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16;
  wire cvt_4_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16;
  wire cvt_5_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16;
  wire cvt_6_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16;
  wire cvt_7_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16;
  wire cvt_8_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16;
  wire cvt_9_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16;
  wire cvt_10_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16;
  wire cvt_11_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16;
  wire cvt_12_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16;
  wire cvt_13_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16;
  wire cvt_14_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16;
  wire cvt_15_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16;
  wire cvt_16_FpIntToFloat_17U_5U_10U_else_i_abs_conc_7_16;
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_16;
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_17;
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_18;
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_19;
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_20;
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_21;
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_22;
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_23;
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_24;
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_25;
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_26;
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_27;
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_28;
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_29;
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_30;
  wire [4:0] libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_31;
  wire chn_idata_data_and_1_cse;
  wire FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse;
  reg [1:0] reg_cfg_proc_precision_1_sva_st_40_cse;
  wire cfg_proc_precision_and_11_cse;
  wire chn_idata_data_and_16_cse;
  wire FpIntToFloat_17U_5U_10U_else_i_abs_and_cse;
  wire IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse;
  wire FpIntToFloat_17U_5U_10U_else_i_abs_and_13_cse;
  wire FpIntToFloat_17U_5U_10U_else_i_abs_and_15_cse;
  wire FpIntToFloat_17U_5U_10U_else_i_abs_and_22_cse;
  wire cfg_proc_precision_and_24_cse;
  wire cfg_proc_precision_and_27_cse;
  wire FpFloatToInt_16U_5U_10U_if_and_cse;
  wire IsNaN_5U_10U_aelse_or_cse;
  wire IsNaN_5U_10U_aelse_or_1_cse;
  wire cvt_else_and_24_cse;
  wire cvt_else_and_34_cse;
  wire IntShiftRightSat_49U_6U_17U_o_and_103_cse;
  wire or_4862_cse;
  wire or_1659_cse_1;
  wire or_1720_cse_1;
  wire or_1752_cse_1;
  wire or_1789_cse_1;
  wire or_1851_cse_1;
  wire or_1892_cse_1;
  wire or_1925_cse_1;
  wire cfg_proc_precision_and_40_cse;
  wire cfg_proc_precision_and_43_cse;
  wire cfg_out_precision_and_32_cse;
  wire FpIntToFloat_17U_5U_10U_if_and_16_cse;
  wire IntShiftRightSat_49U_6U_17U_o_and_115_cse;
  wire IntSaturation_17U_16U_and_33_cse;
  wire IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_27_cse;
  wire IntShiftRightSat_49U_6U_17U_o_and_107_cse;
  wire IntShiftRightSat_49U_6U_17U_o_and_108_cse;
  wire IntShiftRightSat_49U_6U_17U_o_and_109_cse;
  wire IntShiftRightSat_49U_6U_17U_o_and_111_cse;
  wire IntShiftRightSat_49U_6U_17U_o_and_112_cse;
  wire IntShiftRightSat_49U_6U_17U_o_and_114_cse;
  wire or_5038_cse;
  wire or_5053_cse;
  wire or_5069_cse;
  wire or_5086_cse;
  wire nor_1309_cse;
  wire nor_213_cse;
  wire and_976_cse;
  wire and_2396_cse;
  wire and_2402_cse;
  wire and_1038_cse;
  wire and_1039_cse;
  wire or_1198_cse;
  wire or_3817_cse;
  wire nor_1310_cse;
  wire FpIntToFloat_17U_5U_10U_if_and_33_cse;
  wire and_676_cse;
  wire nor_2011_cse;
  wire nor_2004_cse;
  wire nor_2005_cse;
  wire and_978_cse;
  wire mux_1882_cse;
  wire reg_cvt_else_cvt_else_nor_4_cse;
  wire IntShiftRightSat_49U_6U_17U_oelse_and_cse;
  wire IntShiftRightSat_49U_6U_17U_oelse_and_18_cse;
  wire IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_19_cse;
  wire mux_382_cse;
  wire and_283_cse;
  wire IntMulExt_33U_16U_49U_and_11_cse;
  wire or_461_cse;
  wire IntShiftRightSat_49U_6U_17U_if_and_cse;
  wire mux_1762_cse;
  wire and_2275_cse;
  wire IntShiftRightSat_49U_6U_17U_if_and_3_cse;
  wire FpIntToFloat_17U_5U_10U_is_inf_FpIntToFloat_17U_5U_10U_is_inf_or_15_cse;
  wire mux_1071_cse;
  wire FpIntToFloat_17U_5U_10U_is_inf_or_cse;
  wire FpFloatToInt_16U_5U_10U_shift_and_5_cse;
  reg reg_cvt_else_nor_dfs_9_cse;
  wire nor_2150_cse;
  wire mux_110_cse;
  wire mux_1460_cse;
  wire mux_320_cse;
  wire or_3063_cse;
  wire and_2257_cse;
  wire or_4559_cse;
  wire FpIntToFloat_17U_5U_10U_if_and_31_cse;
  wire FpIntToFloat_17U_5U_10U_if_FpIntToFloat_17U_5U_10U_if_or_11_cse;
  wire and_dcpl_1742;
  wire or_tmp;
  wire mux_tmp_2294;
  wire or_tmp_4080;
  wire mux_tmp_2298;
  wire mux_tmp_2300;
  wire or_tmp_4081;
  wire mux_tmp_2304;
  wire mux_tmp_2306;
  wire or_tmp_4082;
  wire mux_tmp_2310;
  wire mux_tmp_2312;
  wire or_tmp_4084;
  wire mux_tmp_2315;
  wire mux_tmp_2317;
  wire mux_tmp_2319;
  wire or_tmp_4086;
  wire mux_tmp_2322;
  wire mux_tmp_2324;
  wire or_tmp_4087;
  wire mux_tmp_2328;
  wire mux_tmp_2330;
  wire mux_tmp_2334;
  wire mux_tmp_2336;
  wire or_tmp_4092;
  wire mux_tmp_2339;
  wire mux_tmp_2341;
  wire or_tmp_4095;
  wire mux_tmp_2345;
  wire mux_tmp_2347;
  wire or_tmp_4097;
  wire mux_tmp_2351;
  wire mux_tmp_2353;
  wire or_5188_tmp;
  wire or_5187_tmp;
  wire or_5186_tmp;
  wire or_5185_tmp;
  wire or_5184_tmp;
  wire or_5183_tmp;
  wire or_5182_tmp;
  wire or_5181_tmp;
  wire or_5180_tmp;
  wire or_5179_tmp;
  wire or_5178_tmp;
  wire or_5177_tmp;
  wire or_5176_tmp;
  wire or_5175_tmp;
  wire or_5174_tmp;
  wire or_tmp_4102;
  wire or_5189_cse;
  wire or_5254_cse;
  wire and_2136_cse;
  wire and_3024_cse;
  wire and_178_itm;
  wire cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_itm_8_1;
  wire cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1;
  wire cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1;
  wire cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1;
  wire cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1;
  wire cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1;
  wire cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1;
  wire cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1;
  wire cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1;
  wire cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1;
  wire cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1;
  wire cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1;
  wire cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1;
  wire cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1;
  wire cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1;
  wire cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1;
  wire cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1;
  wire cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1;
  wire cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1;
  wire cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1;
  wire cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1;
  wire cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1;
  wire cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1;
  wire cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1;
  wire cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1;
  wire cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1;
  wire cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1;
  wire cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1;
  wire cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1;
  wire cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1;
  wire cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_itm_8_1;
  wire cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_itm_7_1;
  wire cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_itm_8_1;
  wire cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1;
  wire cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1;
  wire cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1;
  wire cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1;
  wire cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1;
  wire cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1;
  wire cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1;
  wire cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1;
  wire cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1;
  wire cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1;
  wire cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1;
  wire cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1;
  wire cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1;
  wire cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1;
  wire cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_itm_8_1;
  wire cvt_1_FpFloatToInt_16U_5U_10U_if_acc_itm_11_1;
  wire cvt_2_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1;
  wire cvt_3_IntSaturation_17U_8U_if_acc_1_itm_10_1;
  wire cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1;
  wire cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1;
  wire cvt_5_IntSaturation_17U_8U_if_acc_1_itm_10_1;
  wire cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1;
  wire cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_itm_11_1;
  wire cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1;
  wire cvt_1_IntSaturation_17U_8U_if_acc_itm_10_1;
  wire cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1;
  wire cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1;
  wire cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1;
  wire cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1;
  wire cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1;
  wire cvt_9_IntSaturation_17U_8U_if_acc_1_itm_10_1;
  wire cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1;
  wire cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1;
  wire cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1;
  wire cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1;
  wire cvt_1_IntSaturation_17U_16U_if_acc_itm_2_1;
  wire cvt_2_IntSaturation_17U_16U_if_acc_1_itm_2_1;
  wire cvt_3_IntSaturation_17U_16U_if_acc_1_itm_2_1;
  wire cvt_4_IntSaturation_17U_16U_if_acc_2_itm_2_1;
  wire cvt_5_IntSaturation_17U_16U_if_acc_1_itm_2_1;
  wire cvt_6_IntSaturation_17U_16U_if_acc_2_itm_2_1;
  wire cvt_7_IntSaturation_17U_16U_if_acc_2_itm_2_1;
  wire cvt_8_IntSaturation_17U_16U_if_acc_3_itm_2_1;
  wire cvt_9_IntSaturation_17U_16U_if_acc_1_itm_2_1;
  wire cvt_10_IntSaturation_17U_16U_if_acc_2_itm_2_1;
  wire cvt_11_IntSaturation_17U_16U_if_acc_2_itm_2_1;
  wire cvt_12_IntSaturation_17U_16U_if_acc_3_itm_2_1;
  wire cvt_13_IntSaturation_17U_16U_if_acc_2_itm_2_1;
  wire cvt_14_IntSaturation_17U_16U_if_acc_3_itm_2_1;
  wire cvt_15_IntSaturation_17U_16U_if_acc_3_itm_2_1;
  wire cvt_16_IntSaturation_17U_16U_if_acc_4_itm_2_1;
  wire cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_1_itm_4;
  wire cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4;
  wire cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4;
  wire cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4;
  wire cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4;
  wire cvt_1_IntSaturation_17U_8U_else_if_acc_itm_10;
  wire cvt_2_IntSaturation_17U_8U_else_if_acc_1_itm_10;
  wire cvt_3_IntSaturation_17U_8U_else_if_acc_1_itm_10;
  wire cvt_4_IntSaturation_17U_8U_else_if_acc_2_itm_10;
  wire cvt_5_IntSaturation_17U_8U_else_if_acc_1_itm_10;
  wire cvt_6_IntSaturation_17U_8U_else_if_acc_2_itm_10;
  wire cvt_7_IntSaturation_17U_8U_else_if_acc_2_itm_10;
  wire cvt_8_IntSaturation_17U_8U_else_if_acc_3_itm_10;
  wire cvt_9_IntSaturation_17U_8U_else_if_acc_1_itm_10;
  wire cvt_10_IntSaturation_17U_8U_else_if_acc_2_itm_10;
  wire cvt_11_IntSaturation_17U_8U_else_if_acc_2_itm_10;
  wire cvt_12_IntSaturation_17U_8U_else_if_acc_3_itm_10;
  wire cvt_13_IntSaturation_17U_8U_else_if_acc_2_itm_10;
  wire cvt_15_IntSaturation_17U_8U_else_if_acc_3_itm_10;
  wire cvt_16_IntSaturation_17U_8U_else_if_acc_4_itm_10;
  wire cvt_14_IntSaturation_17U_8U_else_if_acc_3_itm_10;
  wire cvt_1_IntSaturation_17U_16U_else_if_acc_itm_2_1;
  wire cvt_2_IntSaturation_17U_16U_else_if_acc_1_itm_2_1;
  wire cvt_3_IntSaturation_17U_16U_else_if_acc_1_itm_2_1;
  wire cvt_4_IntSaturation_17U_16U_else_if_acc_2_itm_2_1;
  wire cvt_5_IntSaturation_17U_16U_else_if_acc_1_itm_2_1;
  wire cvt_6_IntSaturation_17U_16U_else_if_acc_2_itm_2_1;
  wire cvt_7_IntSaturation_17U_16U_else_if_acc_2_itm_2_1;
  wire cvt_8_IntSaturation_17U_16U_else_if_acc_3_itm_2_1;
  wire cvt_9_IntSaturation_17U_16U_else_if_acc_1_itm_2_1;
  wire cvt_10_IntSaturation_17U_16U_else_if_acc_2_itm_2_1;
  wire cvt_11_IntSaturation_17U_16U_else_if_acc_2_itm_2_1;
  wire cvt_12_IntSaturation_17U_16U_else_if_acc_3_itm_2_1;
  wire cvt_13_IntSaturation_17U_16U_else_if_acc_2_itm_2_1;
  wire cvt_15_IntSaturation_17U_16U_else_if_acc_3_itm_2_1;
  wire cvt_16_IntSaturation_17U_16U_else_if_acc_4_itm_2_1;
  wire cvt_14_IntSaturation_17U_16U_else_if_acc_3_itm_2_1;
  wire IntMulExt_33U_16U_49U_and_1_cse;
  wire or_183_cse_1;
  wire nor_2047_cse;
  wire or_303_cse;
  wire mux_166_cse;
  wire or_306_cse;
  wire nor_1980_cse;
  wire nor_1772_cse;
  wire or_400_cse_1;
  wire mux_1851_cse;
  wire and_2372_cse;
  wire FpIntToFloat_17U_5U_10U_is_inf_and_14_cse;
  wire nor_1500_cse;
  wire nor_1488_cse;
  wire nor_1489_cse;
  wire or_3623_cse;
  wire nand_171_cse;
  wire mux_272_cse;
  wire IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_8_cse;
  wire FpIntToFloat_17U_5U_10U_if_nor_10_cse;
  wire or_186_cse;
  wire mux_133_cse;
  wire or_5379_cse;
  wire mux_1466_cse;
  wire mux_989_cse;
  wire or_2140_cse;
  wire or_3696_cse;
  wire and_1021_cse;
  wire and_1059_cse;
  wire FpFloatToInt_16U_5U_10U_shift_and_1_cse;
  wire FpFloatToInt_16U_5U_10U_shift_and_8_cse;
  wire mux_1761_cse;
  wire mux_1779_cse;
  wire and_2317_cse;
  wire or_3151_cse;
  wire nor_1048_cse;
  wire mux_1881_cse;
  wire mux_1864_cse;
  wire and_2380_cse;
  wire mux_1463_cse;
  wire IntShiftRightSat_49U_6U_17U_o_and_90_cse;
  wire mux_1654_cse;
  wire IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_18_cse;
  wire IntShiftRightSat_49U_6U_17U_oelse_and_25_cse;
  wire FpIntToFloat_17U_5U_10U_if_nor_6_cse;
  wire nor_1486_cse;
  wire and_2246_cse;
  wire or_3774_cse;
  wire and_1249_cse;
  wire nor_2326_cse;
  wire mux_1849_cse;
  wire FpIntToFloat_17U_5U_10U_is_inf_FpIntToFloat_17U_5U_10U_is_inf_or_10_cse;
  wire mux_1437_cse;
  wire mux_786_cse_1;
  wire mux_1489_cse;
  wire mux_1521_cse;
  wire IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_15_cse;
  wire and_3063_cse;
  wire and_174_cse;
  wire and_2259_cse;
  wire nor_1898_cse;
  wire mux_417_cse;
  wire mux_1852_cse;
  wire and_2389_cse;
  wire and_2393_cse;
  wire FpIntToFloat_17U_5U_10U_is_inf_and_26_cse;
  wire FpIntToFloat_17U_5U_10U_if_and_18_cse;
  wire FpIntToFloat_17U_5U_10U_if_and_27_cse;
  wire mux_134_cse;
  wire FpIntToFloat_17U_5U_10U_if_and_22_cse;
  wire IntShiftRightSat_49U_6U_17U_oelse_and_22_cse;
  wire FpIntToFloat_17U_5U_10U_is_inf_and_28_cse;
  wire FpIntToFloat_17U_5U_10U_if_and_36_cse;
  wire mux_1053_cse;
  wire FpIntToFloat_17U_5U_10U_is_inf_and_23_cse;
  wire cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4;
  wire cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4;
  wire cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4;
  wire cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4;
  wire cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4;
  wire cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4;
  wire cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4;
  wire cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4;
  wire cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4;
  wire cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4;
  wire cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_8_tmp_4;
  wire[0:0] shift_0_prb;
  wire[0:0] and_15;
  wire[0:0] shift_0_prb_1;
  wire[0:0] and_19;
  wire[0:0] shift_0_prb_2;
  wire[0:0] and_23;
  wire[0:0] shift_0_prb_3;
  wire[0:0] and_27;
  wire[0:0] shift_0_prb_4;
  wire[0:0] and_32;
  wire[0:0] shift_0_prb_5;
  wire[0:0] and_37;
  wire[0:0] shift_0_prb_6;
  wire[0:0] and_41;
  wire[0:0] shift_0_prb_7;
  wire[0:0] and_45;
  wire[0:0] shift_0_prb_8;
  wire[0:0] and_49;
  wire[0:0] shift_0_prb_9;
  wire[0:0] and_54;
  wire[0:0] shift_0_prb_10;
  wire[0:0] and_58;
  wire[0:0] shift_0_prb_11;
  wire[0:0] and_62;
  wire[0:0] shift_0_prb_12;
  wire[0:0] and_67;
  wire[0:0] shift_0_prb_13;
  wire[0:0] and_71;
  wire[0:0] shift_0_prb_14;
  wire[0:0] and_75;
  wire[0:0] shift_0_prb_15;
  wire[0:0] and_79;
  wire[0:0] iMantWidth_oMantWidth_prb;
  wire[0:0] iExpoWidth_oExpoWidth_prb;
  wire[0:0] iMantWidth_oMantWidth_prb_1;
  wire[0:0] iExpoWidth_oExpoWidth_prb_1;
  wire[0:0] iMantWidth_oMantWidth_prb_2;
  wire[0:0] iExpoWidth_oExpoWidth_prb_2;
  wire[0:0] iMantWidth_oMantWidth_prb_3;
  wire[0:0] iExpoWidth_oExpoWidth_prb_3;
  wire[0:0] iMantWidth_oMantWidth_prb_4;
  wire[0:0] iExpoWidth_oExpoWidth_prb_4;
  wire[0:0] iMantWidth_oMantWidth_prb_5;
  wire[0:0] iExpoWidth_oExpoWidth_prb_5;
  wire[0:0] iMantWidth_oMantWidth_prb_6;
  wire[0:0] iExpoWidth_oExpoWidth_prb_6;
  wire[0:0] iMantWidth_oMantWidth_prb_7;
  wire[0:0] iExpoWidth_oExpoWidth_prb_7;
  wire[0:0] iMantWidth_oMantWidth_prb_8;
  wire[0:0] iExpoWidth_oExpoWidth_prb_8;
  wire[0:0] iMantWidth_oMantWidth_prb_9;
  wire[0:0] iExpoWidth_oExpoWidth_prb_9;
  wire[0:0] iMantWidth_oMantWidth_prb_10;
  wire[0:0] iExpoWidth_oExpoWidth_prb_10;
  wire[0:0] iMantWidth_oMantWidth_prb_11;
  wire[0:0] iExpoWidth_oExpoWidth_prb_11;
  wire[0:0] iMantWidth_oMantWidth_prb_12;
  wire[0:0] iExpoWidth_oExpoWidth_prb_12;
  wire[0:0] iMantWidth_oMantWidth_prb_13;
  wire[0:0] iExpoWidth_oExpoWidth_prb_13;
  wire[0:0] iMantWidth_oMantWidth_prb_14;
  wire[0:0] iExpoWidth_oExpoWidth_prb_14;
  wire[0:0] iMantWidth_oMantWidth_prb_15;
  wire[0:0] iExpoWidth_oExpoWidth_prb_15;
  wire[0:0] oWidth_mWidth_prb;
  wire[0:0] oWidth_aWidth_bWidth_prb;
  wire[0:0] oWidth_iWidth_prb;
  wire[0:0] oWidth_iWidth_prb_1;
  wire[0:0] oWidth_mWidth_prb_1;
  wire[0:0] oWidth_aWidth_bWidth_prb_1;
  wire[0:0] oWidth_iWidth_prb_2;
  wire[0:0] oWidth_iWidth_prb_3;
  wire[0:0] oWidth_mWidth_prb_2;
  wire[0:0] oWidth_aWidth_bWidth_prb_2;
  wire[0:0] oWidth_iWidth_prb_4;
  wire[0:0] oWidth_iWidth_prb_5;
  wire[0:0] oWidth_mWidth_prb_3;
  wire[0:0] oWidth_aWidth_bWidth_prb_3;
  wire[0:0] oWidth_iWidth_prb_6;
  wire[0:0] oWidth_iWidth_prb_7;
  wire[0:0] oWidth_mWidth_prb_4;
  wire[0:0] oWidth_aWidth_bWidth_prb_4;
  wire[0:0] oWidth_iWidth_prb_8;
  wire[0:0] oWidth_iWidth_prb_9;
  wire[0:0] oWidth_mWidth_prb_5;
  wire[0:0] oWidth_aWidth_bWidth_prb_5;
  wire[0:0] oWidth_iWidth_prb_10;
  wire[0:0] oWidth_iWidth_prb_11;
  wire[0:0] oWidth_mWidth_prb_6;
  wire[0:0] oWidth_aWidth_bWidth_prb_6;
  wire[0:0] oWidth_iWidth_prb_12;
  wire[0:0] oWidth_iWidth_prb_13;
  wire[0:0] oWidth_mWidth_prb_7;
  wire[0:0] oWidth_aWidth_bWidth_prb_7;
  wire[0:0] oWidth_iWidth_prb_14;
  wire[0:0] oWidth_iWidth_prb_15;
  wire[0:0] oWidth_mWidth_prb_8;
  wire[0:0] oWidth_aWidth_bWidth_prb_8;
  wire[0:0] oWidth_iWidth_prb_16;
  wire[0:0] oWidth_iWidth_prb_17;
  wire[0:0] oWidth_mWidth_prb_9;
  wire[0:0] oWidth_aWidth_bWidth_prb_9;
  wire[0:0] oWidth_iWidth_prb_18;
  wire[0:0] oWidth_iWidth_prb_19;
  wire[0:0] oWidth_mWidth_prb_10;
  wire[0:0] oWidth_aWidth_bWidth_prb_10;
  wire[0:0] oWidth_iWidth_prb_20;
  wire[0:0] oWidth_iWidth_prb_21;
  wire[0:0] oWidth_mWidth_prb_11;
  wire[0:0] oWidth_aWidth_bWidth_prb_11;
  wire[0:0] oWidth_iWidth_prb_22;
  wire[0:0] oWidth_iWidth_prb_23;
  wire[0:0] oWidth_mWidth_prb_12;
  wire[0:0] oWidth_aWidth_bWidth_prb_12;
  wire[0:0] oWidth_iWidth_prb_24;
  wire[0:0] oWidth_iWidth_prb_25;
  wire[0:0] oWidth_mWidth_prb_13;
  wire[0:0] oWidth_aWidth_bWidth_prb_13;
  wire[0:0] oWidth_iWidth_prb_26;
  wire[0:0] oWidth_iWidth_prb_27;
  wire[0:0] oWidth_mWidth_prb_14;
  wire[0:0] oWidth_aWidth_bWidth_prb_14;
  wire[0:0] oWidth_iWidth_prb_28;
  wire[0:0] oWidth_iWidth_prb_29;
  wire[0:0] oWidth_mWidth_prb_15;
  wire[0:0] oWidth_aWidth_bWidth_prb_15;
  wire[0:0] oWidth_iWidth_prb_30;
  wire[0:0] oWidth_iWidth_prb_31;
  wire[0:0] cvt_and_261_nl;
  wire[0:0] cvt_and_262_nl;
  wire[0:0] SetToInf_5U_10U_SetToInf_5U_10U_or_nl;
  wire[0:0] cvt_and_259_nl;
  wire[0:0] cvt_and_260_nl;
  wire[0:0] and_3148_nl;
  wire[0:0] mux_2302_nl;
  wire[0:0] mux_2301_nl;
  wire[0:0] SetToInf_5U_10U_SetToInf_5U_10U_or_1_nl;
  wire[0:0] cvt_and_257_nl;
  wire[0:0] cvt_and_258_nl;
  wire[0:0] SetToInf_5U_10U_SetToInf_5U_10U_or_2_nl;
  wire[0:0] and_3140_nl;
  wire[0:0] cvt_and_255_nl;
  wire[0:0] cvt_and_256_nl;
  wire[0:0] mux_2308_nl;
  wire[0:0] mux_2307_nl;
  wire[0:0] SetToInf_5U_10U_SetToInf_5U_10U_or_3_nl;
  wire[0:0] cvt_and_253_nl;
  wire[0:0] cvt_and_254_nl;
  wire[0:0] SetToInf_5U_10U_SetToInf_5U_10U_or_4_nl;
  wire[0:0] cvt_and_251_nl;
  wire[0:0] cvt_and_252_nl;
  wire[0:0] and_3136_nl;
  wire[0:0] mux_2314_nl;
  wire[0:0] mux_2313_nl;
  wire[0:0] SetToInf_5U_10U_SetToInf_5U_10U_or_5_nl;
  wire[0:0] cvt_and_249_nl;
  wire[0:0] cvt_and_250_nl;
  wire[0:0] and_3133_nl;
  wire[0:0] mux_2320_nl;
  wire[0:0] mux_2319_nl;
  wire[0:0] SetToInf_5U_10U_SetToInf_5U_10U_or_6_nl;
  wire[0:0] and_3128_nl;
  wire[0:0] cvt_and_247_nl;
  wire[0:0] cvt_and_248_nl;
  wire[0:0] and_3130_nl;
  wire[0:0] mux_2327_nl;
  wire[0:0] mux_2326_nl;
  wire[0:0] SetToInf_5U_10U_SetToInf_5U_10U_or_7_nl;
  wire[0:0] cvt_and_245_nl;
  wire[0:0] cvt_and_246_nl;
  wire[0:0] SetToInf_5U_10U_SetToInf_5U_10U_or_8_nl;
  wire[0:0] cvt_and_243_nl;
  wire[0:0] cvt_and_244_nl;
  wire[0:0] and_3124_nl;
  wire[0:0] mux_2332_nl;
  wire[0:0] mux_2331_nl;
  wire[0:0] SetToInf_5U_10U_SetToInf_5U_10U_or_9_nl;
  wire[0:0] cvt_and_241_nl;
  wire[0:0] cvt_and_242_nl;
  wire[0:0] and_3121_nl;
  wire[0:0] mux_2338_nl;
  wire[0:0] mux_2337_nl;
  wire[0:0] SetToInf_5U_10U_SetToInf_5U_10U_or_10_nl;
  wire[0:0] and_3116_nl;
  wire[0:0] cvt_and_239_nl;
  wire[0:0] cvt_and_240_nl;
  wire[0:0] and_3118_nl;
  wire[0:0] mux_2344_nl;
  wire[0:0] mux_2343_nl;
  wire[0:0] SetToInf_5U_10U_SetToInf_5U_10U_or_11_nl;
  wire[0:0] cvt_and_237_nl;
  wire[0:0] cvt_and_238_nl;
  wire[0:0] and_3115_nl;
  wire[0:0] mux_2349_nl;
  wire[0:0] mux_2348_nl;
  wire[0:0] SetToInf_5U_10U_SetToInf_5U_10U_or_12_nl;
  wire[0:0] mux_2355_nl;
  wire[0:0] mux_2354_nl;
  wire[0:0] and_3110_nl;
  wire[0:0] cvt_and_235_nl;
  wire[0:0] cvt_and_236_nl;
  wire[0:0] and_3112_nl;
  wire[0:0] SetToInf_5U_10U_SetToInf_5U_10U_or_13_nl;
  wire[0:0] cvt_and_233_nl;
  wire[0:0] cvt_and_234_nl;
  wire[0:0] and_3109_nl;
  wire[0:0] mux_2362_nl;
  wire[0:0] mux_2361_nl;
  wire[0:0] mux_2360_nl;
  wire[0:0] SetToInf_5U_10U_SetToInf_5U_10U_or_14_nl;
  wire[0:0] and_3104_nl;
  wire[0:0] cvt_and_231_nl;
  wire[0:0] cvt_and_232_nl;
  wire[0:0] and_3105_nl;
  wire[0:0] SetToInf_5U_10U_SetToInf_5U_10U_or_15_nl;
  wire[0:0] cvt_mux_2281_nl;
  wire[0:0] cvt_if_mux_10_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_mux_4_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_else_mux_2_nl;
  wire[0:0] cvt_mux_2280_nl;
  wire[0:0] cvt_else_mux1h_10_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_or_nl;
  wire[0:0] cvt_or_48_nl;
  wire[0:0] cvt_mux_2373_nl;
  wire[0:0] cvt_else_mux1h_8_nl;
  wire[0:0] cvt_if_mux_8_nl;
  wire[0:0] cvt_mux_2285_nl;
  wire[0:0] cvt_if_mux_25_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_1_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_mux_11_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_else_mux_5_nl;
  wire[0:0] cvt_mux_2284_nl;
  wire[0:0] cvt_else_mux1h_29_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_or_1_nl;
  wire[0:0] cvt_mux_2346_nl;
  wire[0:0] cvt_else_mux1h_27_nl;
  wire[0:0] cvt_if_mux_23_nl;
  wire[0:0] cvt_mux_2289_nl;
  wire[0:0] cvt_if_mux_40_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_2_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_mux_18_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_else_mux_8_nl;
  wire[0:0] cvt_mux_2288_nl;
  wire[0:0] cvt_else_mux1h_48_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_or_2_nl;
  wire[0:0] cvt_mux_2348_nl;
  wire[0:0] cvt_else_mux1h_46_nl;
  wire[0:0] cvt_if_mux_38_nl;
  wire[0:0] cvt_mux_2293_nl;
  wire[0:0] cvt_if_mux_55_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_3_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_mux_25_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_else_mux_11_nl;
  wire[0:0] cvt_mux_2292_nl;
  wire[0:0] cvt_else_mux1h_67_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_or_3_nl;
  wire[0:0] cvt_mux_2350_nl;
  wire[0:0] cvt_else_mux1h_65_nl;
  wire[0:0] cvt_if_mux_53_nl;
  wire[0:0] cvt_mux_2297_nl;
  wire[0:0] cvt_if_mux_70_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_4_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_mux_32_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_else_mux_14_nl;
  wire[0:0] cvt_mux_2296_nl;
  wire[0:0] cvt_else_mux1h_86_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_or_4_nl;
  wire[0:0] cvt_mux_2352_nl;
  wire[0:0] cvt_else_mux1h_84_nl;
  wire[0:0] cvt_if_mux_68_nl;
  wire[0:0] cvt_mux_2301_nl;
  wire[0:0] cvt_if_mux_85_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_5_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_mux_39_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_else_mux_17_nl;
  wire[0:0] cvt_mux_2300_nl;
  wire[0:0] cvt_else_mux1h_105_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_or_5_nl;
  wire[0:0] cvt_mux_2354_nl;
  wire[0:0] cvt_else_mux1h_103_nl;
  wire[0:0] cvt_if_mux_83_nl;
  wire[0:0] cvt_mux_2305_nl;
  wire[0:0] cvt_if_mux_100_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_6_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_mux_46_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_else_mux_20_nl;
  wire[0:0] cvt_mux_2304_nl;
  wire[0:0] cvt_else_mux1h_124_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_or_6_nl;
  wire[0:0] cvt_mux_2358_nl;
  wire[0:0] cvt_else_mux1h_122_nl;
  wire[0:0] cvt_if_mux_98_nl;
  wire[0:0] cvt_mux_2309_nl;
  wire[0:0] cvt_if_mux_115_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_7_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_mux_53_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_else_mux_23_nl;
  wire[0:0] cvt_mux_2308_nl;
  wire[0:0] cvt_else_mux1h_143_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_or_7_nl;
  wire[0:0] cvt_mux_2360_nl;
  wire[0:0] cvt_else_mux1h_141_nl;
  wire[0:0] cvt_if_mux_113_nl;
  wire[0:0] cvt_mux_2313_nl;
  wire[0:0] cvt_if_mux_130_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_8_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_mux_60_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_else_mux_26_nl;
  wire[0:0] cvt_mux_2312_nl;
  wire[0:0] cvt_else_mux1h_162_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_or_8_nl;
  wire[0:0] cvt_mux_2362_nl;
  wire[0:0] cvt_else_mux1h_160_nl;
  wire[0:0] cvt_if_mux_128_nl;
  wire[0:0] cvt_mux_2317_nl;
  wire[0:0] cvt_if_mux_145_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_9_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_mux_67_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_else_mux_29_nl;
  wire[0:0] cvt_mux_2316_nl;
  wire[0:0] cvt_else_mux1h_181_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_or_9_nl;
  wire[0:0] cvt_mux_2364_nl;
  wire[0:0] cvt_else_mux1h_179_nl;
  wire[0:0] cvt_if_mux_143_nl;
  wire[0:0] cvt_mux_2321_nl;
  wire[0:0] cvt_if_mux_160_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_10_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_mux_74_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_else_mux_32_nl;
  wire[0:0] cvt_mux_2320_nl;
  wire[0:0] cvt_else_mux1h_200_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_or_10_nl;
  wire[0:0] cvt_mux_2366_nl;
  wire[0:0] cvt_else_mux1h_198_nl;
  wire[0:0] cvt_if_mux_158_nl;
  wire[0:0] cvt_mux_2325_nl;
  wire[0:0] cvt_if_mux_175_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_11_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_mux_81_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_else_mux_35_nl;
  wire[0:0] cvt_mux_2324_nl;
  wire[0:0] cvt_else_mux1h_219_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_or_11_nl;
  wire[0:0] cvt_mux_2370_nl;
  wire[0:0] cvt_else_mux1h_217_nl;
  wire[0:0] cvt_if_mux_173_nl;
  wire[0:0] cvt_mux_2329_nl;
  wire[0:0] cvt_if_mux_190_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_12_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_mux_88_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_else_mux_38_nl;
  wire[0:0] cvt_mux_2328_nl;
  wire[0:0] cvt_else_mux1h_238_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_or_12_nl;
  wire[0:0] cvt_mux_2372_nl;
  wire[0:0] cvt_else_mux1h_236_nl;
  wire[0:0] cvt_if_mux_188_nl;
  wire[0:0] cvt_mux_2333_nl;
  wire[0:0] cvt_if_mux_205_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_13_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_mux_95_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_else_mux_41_nl;
  wire[0:0] cvt_mux_2332_nl;
  wire[0:0] chn_odata_data_mux_1_nl;
  wire[0:0] cvt_mux_2368_nl;
  wire[0:0] cvt_else_mux1h_255_nl;
  wire[0:0] cvt_if_mux_203_nl;
  wire[0:0] cvt_mux_2337_nl;
  wire[0:0] cvt_if_mux_220_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_14_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_mux_102_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_else_mux_44_nl;
  wire[0:0] cvt_mux_2336_nl;
  wire[0:0] cvt_else_mux1h_276_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_or_14_nl;
  wire[0:0] cvt_mux_2356_nl;
  wire[0:0] cvt_else_mux1h_274_nl;
  wire[0:0] cvt_if_mux_218_nl;
  wire[0:0] cvt_mux_2340_nl;
  wire[0:0] cvt_else_mux1h_295_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_or_15_nl;
  wire[0:0] cvt_if_mux_235_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_15_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_mux_109_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_else_mux_47_nl;
  wire[0:0] cvt_mux_2341_nl;
  wire[0:0] cvt_else_mux1h_292_nl;
  wire[0:0] cvt_if_mux_232_nl;
  wire[0:0] mux_nl;
  wire[0:0] nor_2081_nl;
  wire[0:0] nor_2082_nl;
  wire[0:0] mux_5_nl;
  wire[0:0] and_98_nl;
  wire[0:0] mux_2_nl;
  wire[0:0] or_9_nl;
  wire[0:0] mux_1_nl;
  wire[0:0] or_11_nl;
  wire[0:0] or_13_nl;
  wire[0:0] nor_2080_nl;
  wire[0:0] mux_4_nl;
  wire[0:0] mux_3_nl;
  wire[0:0] and_2240_nl;
  wire[0:0] or_14_nl;
  wire[0:0] and_2242_nl;
  wire[0:0] nor_2_nl;
  wire[0:0] mux_8_nl;
  wire[0:0] or_19_nl;
  wire[0:0] mux_7_nl;
  wire[0:0] nor_10_nl;
  wire[0:0] or_17_nl;
  wire[0:0] mux_10_nl;
  wire[0:0] mux_9_nl;
  wire[0:0] or_28_nl;
  wire[0:0] mux_11_nl;
  wire[0:0] nor_2075_nl;
  wire[0:0] nor_2076_nl;
  wire[0:0] mux_12_nl;
  wire[0:0] mux_14_nl;
  wire[0:0] mux_13_nl;
  wire[0:0] nor_12_nl;
  wire[0:0] or_35_nl;
  wire[0:0] nor_11_nl;
  wire[0:0] mux_16_nl;
  wire[0:0] mux_15_nl;
  wire[0:0] or_37_nl;
  wire[0:0] mux_17_nl;
  wire[0:0] nor_2073_nl;
  wire[0:0] nor_2074_nl;
  wire[0:0] mux_19_nl;
  wire[0:0] mux_18_nl;
  wire[0:0] nor_14_nl;
  wire[0:0] or_43_nl;
  wire[0:0] nor_13_nl;
  wire[0:0] mux_21_nl;
  wire[0:0] mux_20_nl;
  wire[0:0] or_45_nl;
  wire[0:0] mux_22_nl;
  wire[0:0] nor_2071_nl;
  wire[0:0] nor_2072_nl;
  wire[0:0] mux_24_nl;
  wire[0:0] mux_23_nl;
  wire[0:0] nor_16_nl;
  wire[0:0] or_51_nl;
  wire[0:0] nor_15_nl;
  wire[0:0] mux_26_nl;
  wire[0:0] mux_25_nl;
  wire[0:0] or_53_nl;
  wire[0:0] mux_28_nl;
  wire[0:0] mux_27_nl;
  wire[0:0] or_56_nl;
  wire[0:0] or_58_nl;
  wire[0:0] nor_17_nl;
  wire[0:0] mux_30_nl;
  wire[0:0] mux_29_nl;
  wire[0:0] or_61_nl;
  wire[0:0] or_63_nl;
  wire[0:0] nor_18_nl;
  wire[0:0] mux_32_nl;
  wire[0:0] mux_31_nl;
  wire[0:0] nand_235_nl;
  wire[0:0] or_68_nl;
  wire[0:0] mux_34_nl;
  wire[0:0] mux_33_nl;
  wire[0:0] or_71_nl;
  wire[0:0] or_73_nl;
  wire[0:0] nor_19_nl;
  wire[0:0] mux_36_nl;
  wire[0:0] mux_35_nl;
  wire[0:0] or_76_nl;
  wire[0:0] or_78_nl;
  wire[0:0] nor_20_nl;
  wire[0:0] mux_38_nl;
  wire[0:0] mux_37_nl;
  wire[0:0] nand_234_nl;
  wire[0:0] or_83_nl;
  wire[0:0] mux_41_nl;
  wire[0:0] mux_40_nl;
  wire[0:0] or_88_nl;
  wire[0:0] nor_21_nl;
  wire[0:0] mux_42_nl;
  wire[0:0] or_90_nl;
  wire[0:0] nor_22_nl;
  wire[0:0] mux_44_nl;
  wire[0:0] mux_43_nl;
  wire[0:0] nand_233_nl;
  wire[0:0] or_95_nl;
  wire[0:0] mux_45_nl;
  wire[0:0] nor_2069_nl;
  wire[0:0] nor_2070_nl;
  wire[0:0] mux_47_nl;
  wire[0:0] mux_46_nl;
  wire[0:0] nor_24_nl;
  wire[0:0] or_101_nl;
  wire[0:0] nor_23_nl;
  wire[0:0] mux_49_nl;
  wire[0:0] mux_48_nl;
  wire[0:0] or_103_nl;
  wire[0:0] mux_50_nl;
  wire[0:0] nor_2067_nl;
  wire[0:0] nor_2068_nl;
  wire[0:0] mux_52_nl;
  wire[0:0] mux_51_nl;
  wire[0:0] nor_26_nl;
  wire[0:0] or_109_nl;
  wire[0:0] nor_25_nl;
  wire[0:0] mux_54_nl;
  wire[0:0] mux_53_nl;
  wire[0:0] or_111_nl;
  wire[0:0] mux_56_nl;
  wire[0:0] mux_55_nl;
  wire[0:0] or_114_nl;
  wire[0:0] or_116_nl;
  wire[0:0] nor_27_nl;
  wire[0:0] mux_58_nl;
  wire[0:0] mux_57_nl;
  wire[0:0] or_119_nl;
  wire[0:0] or_121_nl;
  wire[0:0] nor_28_nl;
  wire[0:0] mux_60_nl;
  wire[0:0] mux_59_nl;
  wire[0:0] nand_232_nl;
  wire[0:0] or_126_nl;
  wire[0:0] mux_61_nl;
  wire[0:0] nor_2065_nl;
  wire[0:0] nor_2066_nl;
  wire[0:0] mux_63_nl;
  wire[0:0] mux_62_nl;
  wire[0:0] nor_30_nl;
  wire[0:0] or_132_nl;
  wire[0:0] nor_29_nl;
  wire[0:0] mux_65_nl;
  wire[0:0] mux_64_nl;
  wire[0:0] or_134_nl;
  wire[0:0] mux_66_nl;
  wire[0:0] nor_2063_nl;
  wire[0:0] nor_2064_nl;
  wire[0:0] mux_68_nl;
  wire[0:0] mux_67_nl;
  wire[0:0] nor_32_nl;
  wire[0:0] or_140_nl;
  wire[0:0] nor_31_nl;
  wire[0:0] mux_70_nl;
  wire[0:0] mux_69_nl;
  wire[0:0] or_142_nl;
  wire[0:0] mux_72_nl;
  wire[0:0] mux_71_nl;
  wire[0:0] or_145_nl;
  wire[0:0] or_147_nl;
  wire[0:0] nor_33_nl;
  wire[0:0] mux_74_nl;
  wire[0:0] mux_73_nl;
  wire[0:0] or_150_nl;
  wire[0:0] or_152_nl;
  wire[0:0] nor_34_nl;
  wire[0:0] mux_76_nl;
  wire[0:0] mux_75_nl;
  wire[0:0] nand_231_nl;
  wire[0:0] or_157_nl;
  wire[0:0] mux_77_nl;
  wire[0:0] nor_2061_nl;
  wire[0:0] nor_2062_nl;
  wire[0:0] mux_79_nl;
  wire[0:0] mux_78_nl;
  wire[0:0] nor_36_nl;
  wire[0:0] or_163_nl;
  wire[0:0] nor_35_nl;
  wire[0:0] mux_81_nl;
  wire[0:0] mux_80_nl;
  wire[0:0] or_165_nl;
  wire[0:0] mux_82_nl;
  wire[0:0] nor_2059_nl;
  wire[0:0] nor_2060_nl;
  wire[0:0] mux_84_nl;
  wire[0:0] mux_83_nl;
  wire[0:0] nor_38_nl;
  wire[0:0] or_171_nl;
  wire[0:0] nor_37_nl;
  wire[0:0] mux_86_nl;
  wire[0:0] mux_85_nl;
  wire[0:0] or_173_nl;
  wire[0:0] mux_87_nl;
  wire[0:0] nor_2057_nl;
  wire[0:0] nor_2058_nl;
  wire[0:0] mux_89_nl;
  wire[0:0] mux_88_nl;
  wire[0:0] nor_40_nl;
  wire[0:0] or_179_nl;
  wire[0:0] nor_39_nl;
  wire[0:0] mux_91_nl;
  wire[0:0] mux_90_nl;
  wire[0:0] or_181_nl;
  wire[32:0] cvt_2_IntSubExt_32U_32U_33U_o_acc_1_nl;
  wire[33:0] nl_cvt_2_IntSubExt_32U_32U_33U_o_acc_1_nl;
  wire[48:0] cvt_4_IntMulExt_33U_16U_49U_o_mul_2_nl;
  wire[32:0] cvt_4_IntSubExt_32U_32U_33U_o_acc_2_nl;
  wire[33:0] nl_cvt_4_IntSubExt_32U_32U_33U_o_acc_2_nl;
  wire[32:0] cvt_3_IntSubExt_32U_32U_33U_o_acc_1_nl;
  wire[33:0] nl_cvt_3_IntSubExt_32U_32U_33U_o_acc_1_nl;
  wire[48:0] cvt_6_IntMulExt_33U_16U_49U_o_mul_2_nl;
  wire[32:0] cvt_6_IntSubExt_32U_32U_33U_o_acc_2_nl;
  wire[33:0] nl_cvt_6_IntSubExt_32U_32U_33U_o_acc_2_nl;
  wire[48:0] cvt_8_IntMulExt_33U_16U_49U_o_mul_3_nl;
  wire[32:0] cvt_8_IntSubExt_32U_32U_33U_o_acc_3_nl;
  wire[33:0] nl_cvt_8_IntSubExt_32U_32U_33U_o_acc_3_nl;
  wire[48:0] cvt_7_IntMulExt_33U_16U_49U_o_mul_2_nl;
  wire[32:0] cvt_7_IntSubExt_32U_32U_33U_o_acc_2_nl;
  wire[33:0] nl_cvt_7_IntSubExt_32U_32U_33U_o_acc_2_nl;
  wire[32:0] cvt_5_IntSubExt_32U_32U_33U_o_acc_1_nl;
  wire[33:0] nl_cvt_5_IntSubExt_32U_32U_33U_o_acc_1_nl;
  wire[48:0] cvt_10_IntMulExt_33U_16U_49U_o_mul_2_nl;
  wire[32:0] cvt_10_IntSubExt_32U_32U_33U_o_acc_2_nl;
  wire[33:0] nl_cvt_10_IntSubExt_32U_32U_33U_o_acc_2_nl;
  wire[48:0] cvt_12_IntMulExt_33U_16U_49U_o_mul_3_nl;
  wire[32:0] cvt_12_IntSubExt_32U_32U_33U_o_acc_3_nl;
  wire[33:0] nl_cvt_12_IntSubExt_32U_32U_33U_o_acc_3_nl;
  wire[48:0] cvt_11_IntMulExt_33U_16U_49U_o_mul_2_nl;
  wire[32:0] cvt_11_IntSubExt_32U_32U_33U_o_acc_2_nl;
  wire[33:0] nl_cvt_11_IntSubExt_32U_32U_33U_o_acc_2_nl;
  wire[48:0] cvt_14_IntMulExt_33U_16U_49U_o_mul_3_nl;
  wire[32:0] cvt_14_IntSubExt_32U_32U_33U_o_acc_3_nl;
  wire[33:0] nl_cvt_14_IntSubExt_32U_32U_33U_o_acc_3_nl;
  wire[48:0] cvt_16_IntMulExt_33U_16U_49U_o_mul_4_nl;
  wire[32:0] cvt_16_IntSubExt_32U_32U_33U_o_acc_4_nl;
  wire[33:0] nl_cvt_16_IntSubExt_32U_32U_33U_o_acc_4_nl;
  wire[0:0] mux_159_nl;
  wire[0:0] and_132_nl;
  wire[0:0] mux_155_nl;
  wire[0:0] mux_154_nl;
  wire[48:0] cvt_15_IntMulExt_33U_16U_49U_o_mul_3_nl;
  wire[32:0] cvt_15_IntSubExt_32U_32U_33U_o_acc_3_nl;
  wire[33:0] nl_cvt_15_IntSubExt_32U_32U_33U_o_acc_3_nl;
  wire[48:0] cvt_13_IntMulExt_33U_16U_49U_o_mul_2_nl;
  wire[32:0] cvt_13_IntSubExt_32U_32U_33U_o_acc_2_nl;
  wire[33:0] nl_cvt_13_IntSubExt_32U_32U_33U_o_acc_2_nl;
  wire[32:0] cvt_9_IntSubExt_32U_32U_33U_o_acc_1_nl;
  wire[33:0] nl_cvt_9_IntSubExt_32U_32U_33U_o_acc_1_nl;
  wire[32:0] cvt_1_IntSubExt_32U_32U_33U_o_acc_nl;
  wire[33:0] nl_cvt_1_IntSubExt_32U_32U_33U_o_acc_nl;
  wire[0:0] mux_162_nl;
  wire[0:0] nor_2048_nl;
  wire[0:0] mux_163_nl;
  wire[0:0] nor_2046_nl;
  wire[0:0] mux_167_nl;
  wire[0:0] mux_169_nl;
  wire[0:0] mux_175_nl;
  wire[0:0] mux_191_nl;
  wire[0:0] mux_190_nl;
  wire[0:0] mux_192_nl;
  wire[0:0] nor_2026_nl;
  wire[0:0] mux_235_nl;
  wire[0:0] mux_232_nl;
  wire[0:0] and_143_nl;
  wire[0:0] and_145_nl;
  wire[0:0] mux_243_nl;
  wire[0:0] mux_238_nl;
  wire[0:0] mux_237_nl;
  wire[0:0] nor_2020_nl;
  wire[0:0] mux_242_nl;
  wire[0:0] mux_241_nl;
  wire[0:0] and_2857_nl;
  wire[0:0] mux_247_nl;
  wire[0:0] mux_246_nl;
  wire[0:0] nor_2016_nl;
  wire[0:0] nor_2017_nl;
  wire[0:0] mux_248_nl;
  wire[0:0] and_147_nl;
  wire[0:0] mux_257_nl;
  wire[0:0] mux_256_nl;
  wire[0:0] mux_255_nl;
  wire[0:0] mux_254_nl;
  wire[0:0] and_2234_nl;
  wire[0:0] mux_267_nl;
  wire[0:0] mux_261_nl;
  wire[0:0] mux_260_nl;
  wire[0:0] mux_266_nl;
  wire[0:0] mux_265_nl;
  wire[0:0] mux_264_nl;
  wire[0:0] and_2233_nl;
  wire[0:0] mux_271_nl;
  wire[0:0] mux_270_nl;
  wire[0:0] mux_273_nl;
  wire[0:0] mux_275_nl;
  wire[0:0] and_156_nl;
  wire[0:0] and_160_nl;
  wire[0:0] mux_285_nl;
  wire[0:0] mux_280_nl;
  wire[0:0] mux_279_nl;
  wire[0:0] mux_284_nl;
  wire[0:0] mux_283_nl;
  wire[0:0] and_161_nl;
  wire[0:0] mux_289_nl;
  wire[0:0] mux_288_nl;
  wire[0:0] nor_1992_nl;
  wire[0:0] nor_1993_nl;
  wire[0:0] mux_291_nl;
  wire[0:0] and_164_nl;
  wire[0:0] and_166_nl;
  wire[0:0] mux_290_nl;
  wire[0:0] nor_1991_nl;
  wire[0:0] mux_302_nl;
  wire[0:0] mux_296_nl;
  wire[0:0] mux_295_nl;
  wire[0:0] nor_1984_nl;
  wire[0:0] mux_301_nl;
  wire[0:0] mux_300_nl;
  wire[0:0] nor_1985_nl;
  wire[0:0] mux_316_nl;
  wire[0:0] mux_307_nl;
  wire[0:0] mux_306_nl;
  wire[0:0] mux_315_nl;
  wire[0:0] mux_314_nl;
  wire[0:0] and_696_nl;
  wire[0:0] and_699_nl;
  wire[0:0] mux_1752_nl;
  wire[0:0] mux_1751_nl;
  wire[0:0] mux_1750_nl;
  wire[0:0] mux_2174_nl;
  wire[0:0] mux_2173_nl;
  wire[0:0] mux_2172_nl;
  wire[0:0] mux_322_nl;
  wire[0:0] and_168_nl;
  wire[0:0] mux_329_nl;
  wire[0:0] mux_327_nl;
  wire[0:0] mux_328_nl;
  wire[0:0] and_171_nl;
  wire[0:0] mux_338_nl;
  wire[0:0] mux_333_nl;
  wire[0:0] mux_332_nl;
  wire[0:0] mux_337_nl;
  wire[0:0] mux_336_nl;
  wire[0:0] and_172_nl;
  wire[0:0] and_711_nl;
  wire[0:0] and_714_nl;
  wire[0:0] mux_1758_nl;
  wire[0:0] or_3070_nl;
  wire[0:0] mux_1757_nl;
  wire[0:0] mux_2170_nl;
  wire[0:0] mux_2176_nl;
  wire[0:0] mux_2175_nl;
  wire[0:0] and_2265_nl;
  wire[0:0] or_4569_nl;
  wire[0:0] mux_342_nl;
  wire[0:0] nor_1962_nl;
  wire[0:0] mux_341_nl;
  wire[0:0] nor_1958_nl;
  wire[0:0] mux_348_nl;
  wire[0:0] and_173_nl;
  wire[0:0] mux_347_nl;
  wire[0:0] and_2229_nl;
  wire[0:0] mux_359_nl;
  wire[0:0] mux_353_nl;
  wire[0:0] mux_352_nl;
  wire[0:0] nor_1951_nl;
  wire[0:0] mux_358_nl;
  wire[0:0] mux_357_nl;
  wire[0:0] nor_1952_nl;
  wire[0:0] mux_373_nl;
  wire[0:0] mux_364_nl;
  wire[0:0] mux_363_nl;
  wire[0:0] mux_372_nl;
  wire[0:0] mux_371_nl;
  wire[0:0] mux_1760_nl;
  wire[0:0] and_726_nl;
  wire[0:0] and_729_nl;
  wire[0:0] mux_2179_nl;
  wire[0:0] mux_2178_nl;
  wire[0:0] mux_2177_nl;
  wire[0:0] mux_378_nl;
  wire[0:0] nor_1939_nl;
  wire[0:0] mux_383_nl;
  wire[0:0] and_179_nl;
  wire[0:0] and_180_nl;
  wire[0:0] mux_394_nl;
  wire[0:0] mux_388_nl;
  wire[0:0] mux_387_nl;
  wire[0:0] nor_1931_nl;
  wire[0:0] mux_393_nl;
  wire[0:0] mux_392_nl;
  wire[0:0] nor_1932_nl;
  wire[0:0] mux_408_nl;
  wire[0:0] mux_399_nl;
  wire[0:0] mux_398_nl;
  wire[0:0] mux_407_nl;
  wire[0:0] mux_406_nl;
  wire[0:0] and_741_nl;
  wire[0:0] and_744_nl;
  wire[0:0] nor_1917_nl;
  wire[0:0] mux_418_nl;
  wire[0:0] and_182_nl;
  wire[0:0] and_183_nl;
  wire[0:0] mux_431_nl;
  wire[0:0] mux_424_nl;
  wire[0:0] mux_423_nl;
  wire[0:0] nor_1907_nl;
  wire[0:0] mux_430_nl;
  wire[0:0] mux_429_nl;
  wire[0:0] nor_1908_nl;
  wire[0:0] mux_444_nl;
  wire[0:0] mux_437_nl;
  wire[0:0] mux_436_nl;
  wire[0:0] mux_443_nl;
  wire[0:0] mux_442_nl;
  wire[0:0] and_185_nl;
  wire[0:0] and_756_nl;
  wire[0:0] and_759_nl;
  wire[0:0] mux_1772_nl;
  wire[0:0] mux_2186_nl;
  wire[0:0] mux_2185_nl;
  wire[0:0] mux_2183_nl;
  wire[0:0] mux_450_nl;
  wire[0:0] mux_453_nl;
  wire[0:0] mux_458_nl;
  wire[0:0] mux_456_nl;
  wire[0:0] and_2856_nl;
  wire[0:0] mux_467_nl;
  wire[0:0] mux_462_nl;
  wire[0:0] mux_461_nl;
  wire[0:0] mux_466_nl;
  wire[0:0] mux_465_nl;
  wire[0:0] and_194_nl;
  wire[0:0] mux_472_nl;
  wire[0:0] mux_471_nl;
  wire[0:0] nor_1875_nl;
  wire[0:0] mux_478_nl;
  wire[0:0] and_195_nl;
  wire[0:0] mux_477_nl;
  wire[0:0] and_2221_nl;
  wire[0:0] mux_490_nl;
  wire[0:0] mux_483_nl;
  wire[0:0] mux_482_nl;
  wire[0:0] nor_1868_nl;
  wire[0:0] mux_489_nl;
  wire[0:0] mux_488_nl;
  wire[0:0] nor_1869_nl;
  wire[0:0] mux_505_nl;
  wire[0:0] mux_495_nl;
  wire[0:0] mux_494_nl;
  wire[0:0] mux_504_nl;
  wire[0:0] mux_503_nl;
  wire[0:0] mux_2171_nl;
  wire[0:0] and_780_nl;
  wire[0:0] and_783_nl;
  wire[0:0] mux_1780_nl;
  wire[0:0] mux_516_nl;
  wire[0:0] and_199_nl;
  wire[0:0] mux_515_nl;
  wire[0:0] and_2217_nl;
  wire[0:0] mux_528_nl;
  wire[0:0] mux_521_nl;
  wire[0:0] mux_520_nl;
  wire[0:0] nor_1847_nl;
  wire[0:0] mux_527_nl;
  wire[0:0] mux_526_nl;
  wire[0:0] nor_1848_nl;
  wire[0:0] mux_544_nl;
  wire[0:0] mux_533_nl;
  wire[0:0] mux_532_nl;
  wire[0:0] mux_543_nl;
  wire[0:0] mux_542_nl;
  wire[0:0] and_794_nl;
  wire[0:0] and_797_nl;
  wire[0:0] mux_1785_nl;
  wire[0:0] mux_556_nl;
  wire[0:0] and_203_nl;
  wire[0:0] and_205_nl;
  wire[0:0] mux_555_nl;
  wire[0:0] and_2213_nl;
  wire[0:0] mux_569_nl;
  wire[0:0] mux_562_nl;
  wire[0:0] mux_561_nl;
  wire[0:0] nor_1822_nl;
  wire[0:0] mux_568_nl;
  wire[0:0] mux_567_nl;
  wire[0:0] nor_1823_nl;
  wire[0:0] mux_583_nl;
  wire[0:0] mux_575_nl;
  wire[0:0] mux_574_nl;
  wire[0:0] mux_582_nl;
  wire[0:0] mux_581_nl;
  wire[0:0] nor_1814_nl;
  wire[0:0] and_808_nl;
  wire[0:0] and_811_nl;
  wire[0:0] mux_1788_nl;
  wire[0:0] mux_2196_nl;
  wire[0:0] mux_2195_nl;
  wire[0:0] mux_2193_nl;
  wire[0:0] nor_2300_nl;
  wire[0:0] mux_594_nl;
  wire[0:0] and_210_nl;
  wire[0:0] and_212_nl;
  wire[0:0] mux_593_nl;
  wire[0:0] nor_1809_nl;
  wire[0:0] mux_605_nl;
  wire[0:0] mux_599_nl;
  wire[0:0] mux_598_nl;
  wire[0:0] nor_1800_nl;
  wire[0:0] mux_604_nl;
  wire[0:0] mux_603_nl;
  wire[0:0] nor_1801_nl;
  wire[0:0] mux_617_nl;
  wire[0:0] mux_610_nl;
  wire[0:0] mux_609_nl;
  wire[0:0] nor_1793_nl;
  wire[0:0] mux_616_nl;
  wire[0:0] mux_615_nl;
  wire[0:0] nor_1794_nl;
  wire[0:0] and_823_nl;
  wire[0:0] and_826_nl;
  wire[0:0] mux_1791_nl;
  wire[0:0] mux_1790_nl;
  wire[0:0] nand_51_nl;
  wire[0:0] mux_630_nl;
  wire[0:0] and_213_nl;
  wire[0:0] and_215_nl;
  wire[0:0] mux_629_nl;
  wire[0:0] and_2203_nl;
  wire[0:0] mux_644_nl;
  wire[0:0] mux_636_nl;
  wire[0:0] mux_635_nl;
  wire[0:0] or_961_nl;
  wire[0:0] mux_643_nl;
  wire[0:0] mux_642_nl;
  wire[0:0] nor_1773_nl;
  wire[9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_63_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_not_1_nl;
  wire[0:0] or_4348_nl;
  wire[0:0] mux_1799_nl;
  wire[0:0] mux_1794_nl;
  wire[0:0] or_3170_nl;
  wire[0:0] mux_1798_nl;
  wire[0:0] mux_1797_nl;
  wire[0:0] nand_225_nl;
  wire[0:0] mux_1796_nl;
  wire[0:0] and_840_nl;
  wire[0:0] and_843_nl;
  wire[0:0] mux_2214_nl;
  wire[0:0] mux_2213_nl;
  wire[0:0] mux_2212_nl;
  wire[0:0] mux_2211_nl;
  wire[0:0] mux_2210_nl;
  wire[0:0] and_2487_nl;
  wire[0:0] nor_1761_nl;
  wire[0:0] mux_671_nl;
  wire[0:0] and_216_nl;
  wire[0:0] and_218_nl;
  wire[0:0] mux_670_nl;
  wire[0:0] and_2201_nl;
  wire[0:0] mux_684_nl;
  wire[0:0] mux_677_nl;
  wire[0:0] mux_676_nl;
  wire[0:0] nor_1745_nl;
  wire[0:0] mux_683_nl;
  wire[0:0] mux_682_nl;
  wire[0:0] nor_1746_nl;
  wire[0:0] mux_698_nl;
  wire[0:0] mux_690_nl;
  wire[0:0] mux_689_nl;
  wire[0:0] mux_697_nl;
  wire[0:0] mux_696_nl;
  wire[0:0] nor_1737_nl;
  wire[0:0] and_856_nl;
  wire[0:0] and_859_nl;
  wire[0:0] mux_1808_nl;
  wire[0:0] mux_1807_nl;
  wire[0:0] or_3196_nl;
  wire[0:0] mux_2218_nl;
  wire[0:0] mux_2217_nl;
  wire[0:0] mux_2216_nl;
  wire[0:0] mux_2215_nl;
  wire[0:0] nor_2290_nl;
  wire[0:0] mux_715_nl;
  wire[0:0] and_219_nl;
  wire[0:0] and_221_nl;
  wire[0:0] mux_714_nl;
  wire[0:0] and_2196_nl;
  wire[0:0] mux_730_nl;
  wire[0:0] mux_722_nl;
  wire[0:0] mux_721_nl;
  wire[0:0] nor_1708_nl;
  wire[0:0] mux_729_nl;
  wire[0:0] mux_728_nl;
  wire[0:0] nor_1709_nl;
  wire[0:0] mux_746_nl;
  wire[0:0] mux_737_nl;
  wire[0:0] mux_736_nl;
  wire[0:0] nor_1697_nl;
  wire[0:0] mux_745_nl;
  wire[0:0] mux_744_nl;
  wire[0:0] nor_1698_nl;
  wire[0:0] and_873_nl;
  wire[0:0] and_876_nl;
  wire[0:0] mux_1817_nl;
  wire[0:0] mux_1816_nl;
  wire[0:0] mux_1815_nl;
  wire[0:0] or_3220_nl;
  wire[0:0] mux_1814_nl;
  wire[0:0] mux_2223_nl;
  wire[0:0] mux_2222_nl;
  wire[0:0] mux_2221_nl;
  wire[0:0] mux_2219_nl;
  wire[0:0] nor_2287_nl;
  wire[0:0] nor_1683_nl;
  wire[0:0] nor_1674_nl;
  wire[0:0] mux_794_nl;
  wire[0:0] mux_792_nl;
  wire[0:0] mux_793_nl;
  wire[0:0] and_136_nl;
  wire[0:0] mux_796_nl;
  wire[0:0] mux_800_nl;
  wire[10:0] cvt_10_IntSaturation_17U_8U_if_acc_2_nl;
  wire[11:0] nl_cvt_10_IntSaturation_17U_8U_if_acc_2_nl;
  wire[0:0] mux_811_nl;
  wire[0:0] mux_807_nl;
  wire[0:0] mux_805_nl;
  wire[0:0] nor_1667_nl;
  wire[0:0] mux_806_nl;
  wire[0:0] nor_1670_nl;
  wire[0:0] nor_1671_nl;
  wire[0:0] mux_810_nl;
  wire[0:0] mux_808_nl;
  wire[0:0] nand_208_nl;
  wire[0:0] mux_809_nl;
  wire[0:0] or_4532_nl;
  wire[0:0] mux_815_nl;
  wire[0:0] and_227_nl;
  wire[0:0] mux_812_nl;
  wire[0:0] nor_1665_nl;
  wire[0:0] and_228_nl;
  wire[0:0] mux_814_nl;
  wire[0:0] nand_2_nl;
  wire[0:0] mux_818_nl;
  wire[0:0] mux_816_nl;
  wire[0:0] nor_1659_nl;
  wire[0:0] mux_817_nl;
  wire[0:0] nor_1661_nl;
  wire[10:0] cvt_2_IntSaturation_17U_8U_if_acc_1_nl;
  wire[11:0] nl_cvt_2_IntSaturation_17U_8U_if_acc_1_nl;
  wire[0:0] mux_822_nl;
  wire[0:0] and_229_nl;
  wire[0:0] mux_819_nl;
  wire[0:0] nor_1658_nl;
  wire[0:0] and_230_nl;
  wire[0:0] mux_821_nl;
  wire[0:0] nand_3_nl;
  wire[0:0] mux_829_nl;
  wire[0:0] nor_1653_nl;
  wire[0:0] mux_826_nl;
  wire[0:0] mux_825_nl;
  wire[0:0] mux_823_nl;
  wire[0:0] or_1201_nl;
  wire[0:0] nand_4_nl;
  wire[0:0] and_2191_nl;
  wire[0:0] nor_1655_nl;
  wire[0:0] mux_828_nl;
  wire[0:0] or_1209_nl;
  wire[9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_1_nl;
  wire[9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_4_nl;
  wire[9:0] cvt_2_FpMantRNE_17U_11U_else_acc_1_nl;
  wire[10:0] nl_cvt_2_FpMantRNE_17U_11U_else_acc_1_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_if_not_179_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_33_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_34_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_3_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_o_int_and_nl;
  wire[0:0] and_916_nl;
  wire[0:0] and_921_nl;
  wire[0:0] mux_1831_nl;
  wire[0:0] mux_1828_nl;
  wire[0:0] nor_2100_nl;
  wire[0:0] mux_1830_nl;
  wire[0:0] nor_2101_nl;
  wire[0:0] mux_2224_nl;
  wire[0:0] and_2357_nl;
  wire[0:0] mux_833_nl;
  wire[0:0] and_233_nl;
  wire[0:0] mux_830_nl;
  wire[0:0] nor_1652_nl;
  wire[0:0] and_234_nl;
  wire[0:0] mux_832_nl;
  wire[0:0] nand_5_nl;
  wire[9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_2_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_35_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_36_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_5_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_o_int_and_29_nl;
  wire[0:0] mux_2226_nl;
  wire[0:0] mux_2225_nl;
  wire[0:0] nor_2284_nl;
  wire[0:0] or_4718_nl;
  wire[10:0] cvt_4_IntSaturation_17U_8U_if_acc_2_nl;
  wire[11:0] nl_cvt_4_IntSaturation_17U_8U_if_acc_2_nl;
  wire[0:0] mux_837_nl;
  wire[0:0] and_235_nl;
  wire[0:0] mux_834_nl;
  wire[0:0] nor_1649_nl;
  wire[0:0] and_236_nl;
  wire[0:0] mux_836_nl;
  wire[0:0] nand_6_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_37_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_38_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_7_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_o_int_and_28_nl;
  wire[0:0] nor_1049_nl;
  wire[9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_3_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_61_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_62_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_31_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_o_int_and_27_nl;
  wire[0:0] and_945_nl;
  wire[0:0] and_949_nl;
  wire[0:0] mux_2227_nl;
  wire[0:0] and_2371_nl;
  wire[0:0] mux_841_nl;
  wire[0:0] and_237_nl;
  wire[0:0] mux_838_nl;
  wire[0:0] nor_1646_nl;
  wire[0:0] and_238_nl;
  wire[0:0] mux_840_nl;
  wire[0:0] nand_7_nl;
  wire[0:0] mux_1859_nl;
  wire[0:0] and_2156_nl;
  wire[0:0] mux_849_nl;
  wire[0:0] mux_845_nl;
  wire[0:0] mux_843_nl;
  wire[0:0] mux_842_nl;
  wire[0:0] nor_1636_nl;
  wire[0:0] nor_1637_nl;
  wire[0:0] mux_844_nl;
  wire[0:0] nor_1640_nl;
  wire[0:0] nor_1641_nl;
  wire[0:0] mux_848_nl;
  wire[0:0] mux_846_nl;
  wire[0:0] nand_206_nl;
  wire[0:0] mux_847_nl;
  wire[0:0] or_4530_nl;
  wire[0:0] mux_853_nl;
  wire[0:0] and_240_nl;
  wire[0:0] mux_850_nl;
  wire[0:0] nor_1634_nl;
  wire[0:0] and_241_nl;
  wire[0:0] mux_852_nl;
  wire[0:0] nand_9_nl;
  wire[9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_4_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_39_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_40_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_9_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_o_int_and_26_nl;
  wire[0:0] mux_859_nl;
  wire[0:0] mux_856_nl;
  wire[0:0] mux_855_nl;
  wire[0:0] mux_854_nl;
  wire[0:0] nor_1625_nl;
  wire[0:0] mux_858_nl;
  wire[0:0] mux_857_nl;
  wire[0:0] nor_1628_nl;
  wire[0:0] or_1280_nl;
  wire[0:0] nor_1040_nl;
  wire[9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_5_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_59_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_60_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_29_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_o_int_and_25_nl;
  wire[0:0] and_961_nl;
  wire[0:0] and_966_nl;
  wire[0:0] mux_1867_nl;
  wire[0:0] or_4745_nl;
  wire[0:0] mux_2231_nl;
  wire[0:0] mux_2232_nl;
  wire[0:0] or_4755_nl;
  wire[0:0] mux_863_nl;
  wire[0:0] and_242_nl;
  wire[0:0] mux_860_nl;
  wire[0:0] nor_1623_nl;
  wire[0:0] and_243_nl;
  wire[0:0] mux_862_nl;
  wire[0:0] nand_10_nl;
  wire[10:0] cvt_6_IntSaturation_17U_8U_if_acc_2_nl;
  wire[11:0] nl_cvt_6_IntSaturation_17U_8U_if_acc_2_nl;
  wire[0:0] mux_867_nl;
  wire[0:0] and_244_nl;
  wire[0:0] mux_864_nl;
  wire[0:0] nor_1620_nl;
  wire[0:0] and_245_nl;
  wire[0:0] mux_866_nl;
  wire[0:0] nand_11_nl;
  wire[0:0] nor_1033_nl;
  wire[9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_6_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_41_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_42_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_11_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_o_int_and_24_nl;
  wire[0:0] mux_2233_nl;
  wire[0:0] and_2395_nl;
  wire[0:0] mux_1886_nl;
  wire[0:0] and_2154_nl;
  wire[0:0] mux_875_nl;
  wire[0:0] mux_871_nl;
  wire[0:0] mux_869_nl;
  wire[0:0] mux_868_nl;
  wire[0:0] nor_1610_nl;
  wire[0:0] nor_1611_nl;
  wire[0:0] mux_870_nl;
  wire[0:0] nor_1614_nl;
  wire[0:0] nor_1615_nl;
  wire[0:0] mux_874_nl;
  wire[0:0] mux_872_nl;
  wire[0:0] nand_205_nl;
  wire[0:0] mux_873_nl;
  wire[0:0] or_4528_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_57_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_58_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_27_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_o_int_and_23_nl;
  wire[0:0] mux_1889_nl;
  wire[0:0] nor_2142_nl;
  wire[0:0] mux_1888_nl;
  wire[0:0] nor_2143_nl;
  wire[0:0] mux_1832_nl;
  wire[0:0] mux_879_nl;
  wire[0:0] and_247_nl;
  wire[0:0] mux_876_nl;
  wire[0:0] nor_1608_nl;
  wire[0:0] and_248_nl;
  wire[0:0] mux_878_nl;
  wire[0:0] nand_13_nl;
  wire[10:0] cvt_7_IntSaturation_17U_8U_if_acc_2_nl;
  wire[11:0] nl_cvt_7_IntSaturation_17U_8U_if_acc_2_nl;
  wire[0:0] mux_1892_nl;
  wire[0:0] and_2153_nl;
  wire[0:0] mux_887_nl;
  wire[0:0] mux_883_nl;
  wire[0:0] mux_881_nl;
  wire[0:0] mux_880_nl;
  wire[0:0] nor_1598_nl;
  wire[0:0] nor_1599_nl;
  wire[0:0] mux_882_nl;
  wire[0:0] nor_1602_nl;
  wire[0:0] nor_1603_nl;
  wire[0:0] mux_886_nl;
  wire[0:0] mux_884_nl;
  wire[0:0] nand_204_nl;
  wire[0:0] mux_885_nl;
  wire[0:0] or_4526_nl;
  wire[0:0] mux_891_nl;
  wire[0:0] and_250_nl;
  wire[0:0] mux_888_nl;
  wire[0:0] nor_1596_nl;
  wire[0:0] and_251_nl;
  wire[0:0] mux_890_nl;
  wire[0:0] nand_15_nl;
  wire[0:0] mux_899_nl;
  wire[0:0] or_1375_nl;
  wire[0:0] mux_895_nl;
  wire[0:0] mux_894_nl;
  wire[0:0] nand_16_nl;
  wire[0:0] mux_892_nl;
  wire[0:0] nand_17_nl;
  wire[0:0] or_1374_nl;
  wire[0:0] and_2190_nl;
  wire[0:0] mux_898_nl;
  wire[0:0] or_1379_nl;
  wire[0:0] mux_897_nl;
  wire[0:0] or_1383_nl;
  wire[9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_7_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_43_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_44_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_13_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_o_int_and_22_nl;
  wire[10:0] cvt_16_IntSaturation_17U_8U_if_acc_4_nl;
  wire[11:0] nl_cvt_16_IntSaturation_17U_8U_if_acc_4_nl;
  wire[0:0] mux_909_nl;
  wire[0:0] and_2189_nl;
  wire[0:0] mux_906_nl;
  wire[0:0] nor_1584_nl;
  wire[0:0] nor_1585_nl;
  wire[0:0] mux_904_nl;
  wire[0:0] mux_902_nl;
  wire[0:0] or_1393_nl;
  wire[0:0] mux_903_nl;
  wire[0:0] or_1399_nl;
  wire[0:0] or_1396_nl;
  wire[0:0] nor_1588_nl;
  wire[0:0] mux_908_nl;
  wire[0:0] or_1402_nl;
  wire[0:0] or_1409_nl;
  wire[9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_8_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_55_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_56_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_25_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_o_int_and_21_nl;
  wire[0:0] and_999_nl;
  wire[0:0] and_1004_nl;
  wire[0:0] mux_1909_nl;
  wire[0:0] mux_2236_nl;
  wire[0:0] nor_2269_nl;
  wire[0:0] mux_2237_nl;
  wire[0:0] mux_2239_nl;
  wire[0:0] or_4793_nl;
  wire[0:0] mux_913_nl;
  wire[0:0] and_252_nl;
  wire[0:0] mux_910_nl;
  wire[0:0] nor_1583_nl;
  wire[0:0] and_253_nl;
  wire[0:0] mux_912_nl;
  wire[0:0] nand_21_nl;
  wire[10:0] cvt_8_IntSaturation_17U_8U_if_acc_3_nl;
  wire[11:0] nl_cvt_8_IntSaturation_17U_8U_if_acc_3_nl;
  wire[0:0] mux_1916_nl;
  wire[0:0] and_2151_nl;
  wire[0:0] mux_921_nl;
  wire[0:0] mux_917_nl;
  wire[0:0] mux_915_nl;
  wire[0:0] mux_914_nl;
  wire[0:0] nor_1574_nl;
  wire[0:0] nor_1575_nl;
  wire[0:0] mux_916_nl;
  wire[0:0] nor_1577_nl;
  wire[0:0] nor_1578_nl;
  wire[0:0] nor_1579_nl;
  wire[0:0] mux_920_nl;
  wire[0:0] mux_918_nl;
  wire[0:0] or_1431_nl;
  wire[0:0] nand_22_nl;
  wire[0:0] mux_919_nl;
  wire[0:0] mux_925_nl;
  wire[0:0] and_255_nl;
  wire[0:0] mux_922_nl;
  wire[0:0] nor_1572_nl;
  wire[0:0] and_256_nl;
  wire[0:0] mux_924_nl;
  wire[0:0] nand_23_nl;
  wire[9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_9_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_45_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_46_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_15_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_o_int_and_20_nl;
  wire[0:0] and_1013_nl;
  wire[10:0] cvt_15_IntSaturation_17U_8U_if_acc_3_nl;
  wire[11:0] nl_cvt_15_IntSaturation_17U_8U_if_acc_3_nl;
  wire[9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_10_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_53_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_54_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_23_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_o_int_and_19_nl;
  wire[0:0] and_1023_nl;
  wire[0:0] and_1027_nl;
  wire[0:0] mux_1933_nl;
  wire[0:0] mux_1930_nl;
  wire[0:0] and_2149_nl;
  wire[0:0] mux_929_nl;
  wire[0:0] and_257_nl;
  wire[0:0] mux_926_nl;
  wire[0:0] nor_1569_nl;
  wire[0:0] and_258_nl;
  wire[0:0] mux_928_nl;
  wire[0:0] nand_24_nl;
  wire[0:0] mux_933_nl;
  wire[0:0] and_259_nl;
  wire[0:0] mux_930_nl;
  wire[0:0] nor_1566_nl;
  wire[0:0] and_260_nl;
  wire[0:0] mux_932_nl;
  wire[0:0] nand_25_nl;
  wire[9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_11_nl;
  wire[9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_25_nl;
  wire[9:0] cvt_9_FpMantRNE_17U_11U_else_acc_1_nl;
  wire[10:0] nl_cvt_9_FpMantRNE_17U_11U_else_acc_1_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_if_not_200_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_47_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_48_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_17_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_o_int_and_18_nl;
  wire[10:0] cvt_13_IntSaturation_17U_8U_if_acc_2_nl;
  wire[11:0] nl_cvt_13_IntSaturation_17U_8U_if_acc_2_nl;
  wire[9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_12_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_51_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_52_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_21_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_o_int_and_17_nl;
  wire[0:0] mux_937_nl;
  wire[0:0] and_261_nl;
  wire[0:0] mux_934_nl;
  wire[0:0] nor_1563_nl;
  wire[0:0] and_262_nl;
  wire[0:0] mux_936_nl;
  wire[0:0] nand_26_nl;
  wire[10:0] cvt_11_IntSaturation_17U_8U_if_acc_2_nl;
  wire[11:0] nl_cvt_11_IntSaturation_17U_8U_if_acc_2_nl;
  wire[9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_13_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_49_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_50_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_19_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_o_int_and_16_nl;
  wire[10:0] cvt_12_IntSaturation_17U_8U_if_acc_3_nl;
  wire[11:0] nl_cvt_12_IntSaturation_17U_8U_if_acc_3_nl;
  wire[0:0] mux_938_nl;
  wire[0:0] mux_943_nl;
  wire[0:0] mux_940_nl;
  wire[0:0] nor_1557_nl;
  wire[0:0] mux_939_nl;
  wire[0:0] or_1483_nl;
  wire[0:0] or_1484_nl;
  wire[0:0] nor_1558_nl;
  wire[0:0] mux_948_nl;
  wire[0:0] mux_954_nl;
  wire[0:0] mux_950_nl;
  wire[0:0] mux_949_nl;
  wire[0:0] mux_953_nl;
  wire[0:0] mux_951_nl;
  wire[0:0] nor_1555_nl;
  wire[0:0] mux_952_nl;
  wire[0:0] mux_959_nl;
  wire[0:0] nor_1547_nl;
  wire[0:0] nor_1548_nl;
  wire[0:0] mux_964_nl;
  wire[0:0] mux_982_nl;
  wire[0:0] nor_1537_nl;
  wire[0:0] nor_1538_nl;
  wire[0:0] mux_991_nl;
  wire[0:0] mux_985_nl;
  wire[0:0] mux_984_nl;
  wire[0:0] mux_990_nl;
  wire[0:0] mux_988_nl;
  wire[0:0] nor_1536_nl;
  wire[0:0] mux_995_nl;
  wire[0:0] mux_1000_nl;
  wire[0:0] nor_1526_nl;
  wire[0:0] nor_1527_nl;
  wire[0:0] mux_1003_nl;
  wire[0:0] mux_1001_nl;
  wire[0:0] nor_1523_nl;
  wire[0:0] mux_1002_nl;
  wire[0:0] nor_1524_nl;
  wire[0:0] nor_1525_nl;
  wire[0:0] FpMantRNE_17U_11U_else_mux_1_nl;
  wire[0:0] or_3841_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_else_mux_1_nl;
  wire[0:0] mux_1004_nl;
  wire[0:0] nor_1519_nl;
  wire[0:0] nor_1521_nl;
  wire[4:0] cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_nl;
  wire[5:0] nl_cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_or_15_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_and_31_nl;
  wire[0:0] mux_2250_nl;
  wire[0:0] and_2811_nl;
  wire[0:0] mux_2251_nl;
  wire[0:0] nor_2461_nl;
  wire[0:0] mux_1011_nl;
  wire[0:0] nor_1510_nl;
  wire[0:0] mux_1010_nl;
  wire[0:0] nor_1511_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_nor_1_nl;
  wire[0:0] FpMantRNE_17U_11U_else_mux_3_nl;
  wire[0:0] or_3850_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_else_mux_4_nl;
  wire[0:0] mux_1018_nl;
  wire[0:0] mux_1016_nl;
  wire[0:0] mux_1012_nl;
  wire[0:0] nor_1508_nl;
  wire[0:0] mux_1017_nl;
  wire[4:0] cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl;
  wire[5:0] nl_cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_or_14_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_and_29_nl;
  wire[0:0] mux_2252_nl;
  wire[0:0] and_2809_nl;
  wire[0:0] mux_2253_nl;
  wire[0:0] nor_2457_nl;
  wire[9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_7_nl;
  wire[9:0] cvt_3_FpMantRNE_17U_11U_else_acc_1_nl;
  wire[10:0] nl_cvt_3_FpMantRNE_17U_11U_else_acc_1_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_if_not_182_nl;
  wire[0:0] mux_1027_nl;
  wire[0:0] nor_1498_nl;
  wire[0:0] FpMantRNE_17U_11U_else_mux_5_nl;
  wire[0:0] or_3860_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_else_mux_7_nl;
  wire[4:0] cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl;
  wire[5:0] nl_cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_or_13_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_and_27_nl;
  wire[0:0] mux_2254_nl;
  wire[0:0] and_2807_nl;
  wire[0:0] mux_2255_nl;
  wire[0:0] nor_2453_nl;
  wire[0:0] mux_1035_nl;
  wire[0:0] mux_1034_nl;
  wire[0:0] mux_1051_nl;
  wire[0:0] mux_1050_nl;
  wire[0:0] mux_1052_nl;
  wire[0:0] mux_1054_nl;
  wire[0:0] mux_1045_nl;
  wire[0:0] mux_1044_nl;
  wire[4:0] cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  wire[5:0] nl_cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_or_12_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_and_25_nl;
  wire[0:0] mux_2256_nl;
  wire[0:0] and_2805_nl;
  wire[0:0] mux_2257_nl;
  wire[0:0] nor_2449_nl;
  wire[0:0] FpMantRNE_17U_11U_else_mux_9_nl;
  wire[0:0] or_3879_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_else_mux_13_nl;
  wire[4:0] cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl;
  wire[5:0] nl_cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_or_11_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_and_23_nl;
  wire[0:0] mux_2258_nl;
  wire[0:0] and_2803_nl;
  wire[0:0] mux_2259_nl;
  wire[0:0] nor_2445_nl;
  wire[0:0] mux_1070_nl;
  wire[0:0] nor_1465_nl;
  wire[0:0] mux_1069_nl;
  wire[0:0] nor_1466_nl;
  wire[0:0] nor_1463_nl;
  wire[0:0] mux_1077_nl;
  wire[0:0] mux_1075_nl;
  wire[0:0] mux_1076_nl;
  wire[4:0] cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  wire[5:0] nl_cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_or_10_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_and_21_nl;
  wire[0:0] mux_2260_nl;
  wire[0:0] and_2801_nl;
  wire[0:0] mux_2261_nl;
  wire[0:0] nor_2441_nl;
  wire[0:0] mux_1091_nl;
  wire[0:0] mux_1089_nl;
  wire[0:0] mux_1090_nl;
  wire[4:0] cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  wire[5:0] nl_cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_or_9_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_and_19_nl;
  wire[0:0] mux_2262_nl;
  wire[0:0] and_2799_nl;
  wire[0:0] mux_2263_nl;
  wire[0:0] nor_2437_nl;
  wire[0:0] mux_1116_nl;
  wire[0:0] mux_1107_nl;
  wire[0:0] mux_1106_nl;
  wire[0:0] mux_1115_nl;
  wire[0:0] mux_1113_nl;
  wire[0:0] mux_1112_nl;
  wire[0:0] mux_1114_nl;
  wire[4:0] cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl;
  wire[5:0] nl_cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_or_8_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_and_17_nl;
  wire[0:0] mux_2264_nl;
  wire[0:0] and_2797_nl;
  wire[0:0] mux_2265_nl;
  wire[0:0] nor_2433_nl;
  wire[0:0] nor_1434_nl;
  wire[0:0] FpMantRNE_17U_11U_else_mux_17_nl;
  wire[0:0] or_3920_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_else_mux_25_nl;
  wire[0:0] mux_1127_nl;
  wire[0:0] nor_1433_nl;
  wire[4:0] cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl;
  wire[5:0] nl_cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_or_7_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_and_15_nl;
  wire[0:0] mux_2266_nl;
  wire[0:0] and_2795_nl;
  wire[0:0] mux_2267_nl;
  wire[0:0] nor_2429_nl;
  wire[0:0] mux_1134_nl;
  wire[0:0] mux_1133_nl;
  wire[4:0] cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  wire[5:0] nl_cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_or_6_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_and_13_nl;
  wire[0:0] mux_2268_nl;
  wire[0:0] and_2793_nl;
  wire[0:0] mux_2269_nl;
  wire[0:0] nor_2425_nl;
  wire[0:0] nor_1415_nl;
  wire[0:0] mux_1163_nl;
  wire[0:0] mux_1154_nl;
  wire[0:0] mux_1153_nl;
  wire[4:0] cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  wire[5:0] nl_cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_or_5_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_and_11_nl;
  wire[0:0] mux_2270_nl;
  wire[0:0] and_2791_nl;
  wire[0:0] mux_2271_nl;
  wire[0:0] and_2789_nl;
  wire[0:0] mux_1179_nl;
  wire[0:0] mux_1174_nl;
  wire[0:0] mux_1173_nl;
  wire[0:0] mux_1172_nl;
  wire[0:0] and_3372_nl;
  wire[0:0] mux_1178_nl;
  wire[0:0] mux_1177_nl;
  wire[0:0] mux_1176_nl;
  wire[0:0] mux_1175_nl;
  wire[0:0] nor_1403_nl;
  wire[0:0] or_1918_nl;
  wire[4:0] cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl;
  wire[5:0] nl_cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_or_4_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_and_9_nl;
  wire[0:0] mux_2272_nl;
  wire[0:0] and_2788_nl;
  wire[0:0] mux_2273_nl;
  wire[0:0] and_3373_nl;
  wire[4:0] cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  wire[5:0] nl_cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_or_3_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_and_7_nl;
  wire[0:0] mux_2274_nl;
  wire[0:0] and_2786_nl;
  wire[0:0] mux_2275_nl;
  wire[0:0] nor_2411_nl;
  wire[10:0] cvt_14_IntSaturation_17U_8U_if_acc_3_nl;
  wire[11:0] nl_cvt_14_IntSaturation_17U_8U_if_acc_3_nl;
  wire[0:0] mux_1204_nl;
  wire[0:0] nand_45_nl;
  wire[0:0] mux_1203_nl;
  wire[0:0] mux_1202_nl;
  wire[0:0] nand_201_nl;
  wire[0:0] mux_1213_nl;
  wire[0:0] nand_46_nl;
  wire[0:0] mux_1212_nl;
  wire[0:0] mux_1211_nl;
  wire[0:0] nand_199_nl;
  wire[4:0] cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl;
  wire[5:0] nl_cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_or_2_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_and_5_nl;
  wire[0:0] mux_2276_nl;
  wire[0:0] and_2784_nl;
  wire[0:0] mux_2277_nl;
  wire[0:0] nor_2406_nl;
  wire[0:0] mux_2000_nl;
  wire[4:0] cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl;
  wire[5:0] nl_cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_or_1_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_and_3_nl;
  wire[0:0] mux_2278_nl;
  wire[0:0] and_2782_nl;
  wire[0:0] mux_2279_nl;
  wire[0:0] nor_2401_nl;
  wire[4:0] cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_9_nl;
  wire[5:0] nl_cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_9_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_or_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_o_expo_and_1_nl;
  wire[0:0] mux_2280_nl;
  wire[0:0] and_2780_nl;
  wire[0:0] mux_2281_nl;
  wire[0:0] nor_2396_nl;
  wire[0:0] mux_1262_nl;
  wire[0:0] and_223_nl;
  wire[0:0] mux_1252_nl;
  wire[0:0] nor_1351_nl;
  wire[0:0] mux_1266_nl;
  wire[0:0] mux_1265_nl;
  wire[0:0] nor_1338_nl;
  wire[0:0] mux_1267_nl;
  wire[0:0] and_271_nl;
  wire[0:0] mux_1268_nl;
  wire[0:0] and_295_nl;
  wire[17:0] cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl;
  wire[18:0] nl_cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl;
  wire[0:0] IntShiftRightSat_49U_6U_17U_oelse_mux_24_nl;
  wire[14:0] FpFloatToInt_16U_5U_10U_o_int_mux1h_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_32_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_and_1_nl;
  wire[0:0] FpFloatToInt_16U_5U_10U_o_int_and_15_nl;
  wire[0:0] and_908_nl;
  wire[9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_14_nl;
  wire[9:0] FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_1_nl;
  wire[9:0] cvt_1_FpMantRNE_17U_11U_else_acc_nl;
  wire[10:0] nl_cvt_1_FpMantRNE_17U_11U_else_acc_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_if_not_176_nl;
  wire[0:0] and_1179_nl;
  wire[0:0] mux_2015_nl;
  wire[0:0] or_3597_nl;
  wire[0:0] mux_2011_nl;
  wire[0:0] mux_2010_nl;
  wire[0:0] mux_2014_nl;
  wire[0:0] mux_2012_nl;
  wire[0:0] mux_2013_nl;
  wire[0:0] or_3600_nl;
  wire[0:0] mux_2020_nl;
  wire[0:0] or_3606_nl;
  wire[0:0] mux_2017_nl;
  wire[0:0] mux_2019_nl;
  wire[0:0] or_3607_nl;
  wire[0:0] mux_2018_nl;
  wire[0:0] or_3609_nl;
  wire[0:0] mux_2249_nl;
  wire[0:0] mux_2248_nl;
  wire[0:0] nor_2251_nl;
  wire[0:0] or_4857_nl;
  wire[0:0] nor_2252_nl;
  wire[17:0] cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl;
  wire[18:0] nl_cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl;
  wire[0:0] IntShiftRightSat_49U_6U_17U_oelse_mux_26_nl;
  wire[17:0] cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl;
  wire[18:0] nl_cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl;
  wire[0:0] IntShiftRightSat_49U_6U_17U_oelse_mux_22_nl;
  wire[17:0] cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  wire[18:0] nl_cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  wire[0:0] IntShiftRightSat_49U_6U_17U_oelse_mux_28_nl;
  wire[17:0] cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl;
  wire[18:0] nl_cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl;
  wire[0:0] IntShiftRightSat_49U_6U_17U_oelse_mux_18_nl;
  wire[17:0] cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  wire[18:0] nl_cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  wire[0:0] IntShiftRightSat_49U_6U_17U_oelse_mux_20_nl;
  wire[17:0] cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  wire[18:0] nl_cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  wire[0:0] IntShiftRightSat_49U_6U_17U_oelse_mux_16_nl;
  wire[17:0] cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl;
  wire[18:0] nl_cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl;
  wire[0:0] IntShiftRightSat_49U_6U_17U_oelse_mux_30_nl;
  wire[17:0] cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl;
  wire[18:0] nl_cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl;
  wire[0:0] IntShiftRightSat_49U_6U_17U_oelse_mux_10_nl;
  wire[17:0] cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  wire[18:0] nl_cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  wire[0:0] IntShiftRightSat_49U_6U_17U_oelse_mux_12_nl;
  wire[17:0] cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  wire[18:0] nl_cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  wire[0:0] IntShiftRightSat_49U_6U_17U_oelse_mux_8_nl;
  wire[17:0] cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl;
  wire[18:0] nl_cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl;
  wire[0:0] IntShiftRightSat_49U_6U_17U_oelse_mux_14_nl;
  wire[17:0] cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  wire[18:0] nl_cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl;
  wire[0:0] IntShiftRightSat_49U_6U_17U_oelse_mux_4_nl;
  wire[17:0] cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl;
  wire[18:0] nl_cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl;
  wire[0:0] IntShiftRightSat_49U_6U_17U_oelse_mux_6_nl;
  wire[17:0] cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl;
  wire[18:0] nl_cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl;
  wire[0:0] IntShiftRightSat_49U_6U_17U_oelse_mux_2_nl;
  wire[17:0] cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl;
  wire[18:0] nl_cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl;
  wire[0:0] IntShiftRightSat_49U_6U_17U_oelse_mux_32_nl;
  wire[0:0] mux_1345_nl;
  wire[0:0] mux_1344_nl;
  wire[0:0] mux_1343_nl;
  wire[0:0] mux_1342_nl;
  wire[0:0] mux_1429_nl;
  wire[0:0] mux_1428_nl;
  wire[0:0] mux_1427_nl;
  wire[0:0] mux_1426_nl;
  wire[0:0] mux_1425_nl;
  wire[0:0] mux_1424_nl;
  wire[0:0] mux_1423_nl;
  wire[0:0] mux_1421_nl;
  wire[0:0] mux_1420_nl;
  wire[0:0] or_2251_nl;
  wire[0:0] or_2242_nl;
  wire[0:0] nor_1314_nl;
  wire[0:0] mux_1442_nl;
  wire[0:0] mux_1441_nl;
  wire[0:0] mux_1439_nl;
  wire[0:0] mux_1438_nl;
  wire[0:0] mux_1458_nl;
  wire[0:0] nor_1306_nl;
  wire[0:0] nor_2130_nl;
  wire[0:0] nor_1305_nl;
  wire[0:0] mux_1465_nl;
  wire[0:0] mux_1461_nl;
  wire[0:0] nor_2114_nl;
  wire[0:0] nor_1301_nl;
  wire[0:0] mux_1472_nl;
  wire[0:0] mux_1467_nl;
  wire[0:0] nor_2113_nl;
  wire[0:0] mux_1471_nl;
  wire[0:0] nor_1302_nl;
  wire[0:0] mux_1470_nl;
  wire[0:0] nor_1303_nl;
  wire[0:0] nor_2127_nl;
  wire[0:0] nor_1287_nl;
  wire[0:0] mux_1495_nl;
  wire[0:0] mux_1490_nl;
  wire[0:0] nor_2110_nl;
  wire[0:0] mux_1519_nl;
  wire[0:0] nor_1271_nl;
  wire[0:0] mux_124_nl;
  wire[0:0] mux_130_nl;
  wire[0:0] mux_118_nl;
  wire[0:0] mux_149_nl;
  wire[0:0] mux_152_nl;
  wire[0:0] mux_1533_nl;
  wire[0:0] mux_1532_nl;
  wire[0:0] mux_1531_nl;
  wire[0:0] or_2433_nl;
  wire[0:0] mux_1534_nl;
  wire[0:0] nor_1263_nl;
  wire[0:0] nor_1264_nl;
  wire[0:0] mux_1535_nl;
  wire[0:0] nor_1261_nl;
  wire[0:0] nor_1262_nl;
  wire[0:0] mux_1536_nl;
  wire[0:0] nor_1259_nl;
  wire[0:0] nor_1260_nl;
  wire[0:0] mux_1537_nl;
  wire[0:0] nor_1257_nl;
  wire[0:0] nor_1258_nl;
  wire[0:0] mux_1538_nl;
  wire[0:0] nor_1255_nl;
  wire[0:0] nor_1256_nl;
  wire[0:0] mux_1539_nl;
  wire[0:0] nor_1253_nl;
  wire[0:0] nor_1254_nl;
  wire[0:0] mux_1540_nl;
  wire[0:0] nor_1251_nl;
  wire[0:0] nor_1252_nl;
  wire[0:0] mux_1541_nl;
  wire[0:0] nor_1249_nl;
  wire[0:0] nor_1250_nl;
  wire[0:0] mux_1542_nl;
  wire[0:0] nor_1247_nl;
  wire[0:0] nor_1248_nl;
  wire[0:0] mux_1543_nl;
  wire[0:0] nor_1245_nl;
  wire[0:0] nor_1246_nl;
  wire[0:0] mux_1544_nl;
  wire[0:0] nor_1243_nl;
  wire[0:0] nor_1244_nl;
  wire[0:0] mux_1545_nl;
  wire[0:0] nor_1241_nl;
  wire[0:0] nor_1242_nl;
  wire[0:0] mux_1546_nl;
  wire[0:0] nor_1239_nl;
  wire[0:0] nor_1240_nl;
  wire[0:0] mux_1547_nl;
  wire[0:0] nor_1237_nl;
  wire[0:0] nor_1238_nl;
  wire[0:0] mux_1548_nl;
  wire[0:0] nor_1235_nl;
  wire[0:0] nor_1236_nl;
  wire[0:0] mux_1549_nl;
  wire[0:0] nor_1233_nl;
  wire[0:0] nor_1234_nl;
  wire[0:0] mux_1550_nl;
  wire[0:0] nor_1231_nl;
  wire[0:0] nor_1232_nl;
  wire[0:0] mux_1551_nl;
  wire[0:0] nor_1229_nl;
  wire[0:0] nor_1230_nl;
  wire[0:0] mux_1552_nl;
  wire[0:0] nor_1227_nl;
  wire[0:0] nor_1228_nl;
  wire[0:0] mux_1553_nl;
  wire[0:0] nor_1225_nl;
  wire[0:0] nor_1226_nl;
  wire[0:0] mux_1554_nl;
  wire[0:0] nor_1223_nl;
  wire[0:0] nor_1224_nl;
  wire[0:0] mux_1555_nl;
  wire[0:0] nor_1221_nl;
  wire[0:0] nor_1222_nl;
  wire[0:0] mux_1556_nl;
  wire[0:0] nor_1219_nl;
  wire[0:0] nor_1220_nl;
  wire[0:0] mux_1557_nl;
  wire[0:0] nor_1217_nl;
  wire[0:0] nor_1218_nl;
  wire[0:0] mux_1558_nl;
  wire[0:0] nor_1215_nl;
  wire[0:0] nor_1216_nl;
  wire[0:0] mux_1559_nl;
  wire[0:0] nor_1213_nl;
  wire[0:0] nor_1214_nl;
  wire[0:0] mux_1560_nl;
  wire[0:0] nor_1211_nl;
  wire[0:0] nor_1212_nl;
  wire[0:0] mux_1561_nl;
  wire[0:0] nor_1209_nl;
  wire[0:0] nor_1210_nl;
  wire[0:0] mux_1562_nl;
  wire[0:0] nor_1207_nl;
  wire[0:0] nor_1208_nl;
  wire[0:0] mux_1563_nl;
  wire[0:0] nor_1205_nl;
  wire[0:0] nor_1206_nl;
  wire[0:0] mux_1564_nl;
  wire[0:0] nor_1203_nl;
  wire[0:0] nor_1204_nl;
  wire[0:0] mux_1565_nl;
  wire[0:0] nor_1201_nl;
  wire[0:0] nor_1202_nl;
  wire[0:0] mux_1569_nl;
  wire[0:0] mux_1567_nl;
  wire[0:0] mux_1568_nl;
  wire[0:0] nor_597_nl;
  wire[0:0] FpMantRNE_24U_11U_else_mux_31_nl;
  wire[0:0] mux_1573_nl;
  wire[0:0] mux_1571_nl;
  wire[0:0] mux_1572_nl;
  wire[0:0] nor_598_nl;
  wire[0:0] FpMantRNE_24U_11U_else_mux_29_nl;
  wire[0:0] mux_1577_nl;
  wire[0:0] mux_1575_nl;
  wire[0:0] mux_1576_nl;
  wire[0:0] nor_599_nl;
  wire[0:0] FpMantRNE_24U_11U_else_mux_27_nl;
  wire[0:0] mux_1581_nl;
  wire[0:0] mux_1579_nl;
  wire[0:0] mux_1580_nl;
  wire[0:0] nor_600_nl;
  wire[0:0] FpMantRNE_24U_11U_else_mux_25_nl;
  wire[0:0] mux_1585_nl;
  wire[0:0] mux_1583_nl;
  wire[0:0] mux_1584_nl;
  wire[0:0] nor_601_nl;
  wire[0:0] FpMantRNE_24U_11U_else_mux_23_nl;
  wire[0:0] mux_1589_nl;
  wire[0:0] mux_1587_nl;
  wire[0:0] mux_1588_nl;
  wire[0:0] nor_602_nl;
  wire[0:0] FpMantRNE_24U_11U_else_mux_21_nl;
  wire[0:0] mux_1591_nl;
  wire[0:0] mux_1590_nl;
  wire[0:0] and_2243_nl;
  wire[0:0] and_2162_nl;
  wire[0:0] nor_603_nl;
  wire[0:0] nor_1200_nl;
  wire[0:0] FpMantRNE_24U_11U_else_mux_19_nl;
  wire[0:0] mux_1595_nl;
  wire[0:0] mux_1593_nl;
  wire[0:0] mux_1594_nl;
  wire[0:0] nor_605_nl;
  wire[0:0] FpMantRNE_24U_11U_else_mux_17_nl;
  wire[0:0] mux_1599_nl;
  wire[0:0] mux_1597_nl;
  wire[0:0] mux_1598_nl;
  wire[0:0] nor_606_nl;
  wire[0:0] FpMantRNE_24U_11U_else_mux_15_nl;
  wire[0:0] mux_1603_nl;
  wire[0:0] mux_1601_nl;
  wire[0:0] mux_1602_nl;
  wire[0:0] nor_607_nl;
  wire[0:0] FpMantRNE_24U_11U_else_mux_13_nl;
  wire[0:0] mux_1605_nl;
  wire[0:0] mux_1604_nl;
  wire[0:0] and_nl;
  wire[0:0] and_2161_nl;
  wire[0:0] nor_608_nl;
  wire[0:0] nor_1198_nl;
  wire[0:0] FpMantRNE_24U_11U_else_mux_11_nl;
  wire[0:0] mux_1609_nl;
  wire[0:0] mux_1607_nl;
  wire[0:0] mux_1608_nl;
  wire[0:0] nor_610_nl;
  wire[0:0] FpMantRNE_24U_11U_else_mux_9_nl;
  wire[0:0] mux_1613_nl;
  wire[0:0] mux_1611_nl;
  wire[0:0] mux_1612_nl;
  wire[0:0] nor_611_nl;
  wire[0:0] FpMantRNE_24U_11U_else_mux_7_nl;
  wire[0:0] mux_1617_nl;
  wire[0:0] mux_1615_nl;
  wire[0:0] mux_1616_nl;
  wire[0:0] nor_612_nl;
  wire[0:0] FpMantRNE_24U_11U_else_mux_5_nl;
  wire[0:0] mux_1621_nl;
  wire[0:0] mux_1619_nl;
  wire[0:0] mux_1620_nl;
  wire[0:0] nor_613_nl;
  wire[0:0] FpMantRNE_24U_11U_else_mux_3_nl;
  wire[0:0] mux_1625_nl;
  wire[0:0] mux_1623_nl;
  wire[0:0] mux_1624_nl;
  wire[0:0] nor_614_nl;
  wire[0:0] FpMantRNE_24U_11U_else_mux_1_nl;
  wire[0:0] mux_1626_nl;
  wire[0:0] nor_1195_nl;
  wire[0:0] mux_1627_nl;
  wire[0:0] and_2160_nl;
  wire[0:0] IsNaN_5U_10U_nor_nl;
  wire[0:0] mux_1640_nl;
  wire[0:0] mux_1633_nl;
  wire[0:0] mux_1632_nl;
  wire[0:0] mux_1639_nl;
  wire[0:0] mux_1638_nl;
  wire[0:0] IsNaN_5U_10U_IsNaN_5U_10U_nand_nl;
  wire[0:0] mux_1649_nl;
  wire[0:0] mux_1644_nl;
  wire[0:0] mux_1643_nl;
  wire[0:0] mux_1648_nl;
  wire[0:0] mux_1647_nl;
  wire[0:0] mux_1653_nl;
  wire[0:0] IsNaN_5U_10U_nor_1_nl;
  wire[0:0] mux_1660_nl;
  wire[0:0] mux_1659_nl;
  wire[0:0] mux_1658_nl;
  wire[0:0] IsNaN_5U_10U_IsNaN_5U_10U_nand_1_nl;
  wire[0:0] mux_1663_nl;
  wire[0:0] mux_1661_nl;
  wire[0:0] mux_1662_nl;
  wire[0:0] IsNaN_5U_10U_nor_14_nl;
  wire[0:0] mux_1674_nl;
  wire[0:0] mux_1673_nl;
  wire[0:0] mux_1672_nl;
  wire[0:0] IsNaN_5U_10U_IsNaN_5U_10U_nand_14_nl;
  wire[0:0] mux_1685_nl;
  wire[0:0] mux_1684_nl;
  wire[0:0] mux_1683_nl;
  wire[0:0] or_479_nl;
  wire[0:0] or_547_nl;
  wire[0:0] mux_377_nl;
  wire[0:0] or_626_nl;
  wire[0:0] mux_449_nl;
  wire[0:0] or_724_nl;
  wire[0:0] mux_454_nl;
  wire[0:0] or_733_nl;
  wire[0:0] mux_770_nl;
  wire[0:0] or_1118_nl;
  wire[0:0] mux_789_nl;
  wire[0:0] or_1134_nl;
  wire[0:0] mux_799_nl;
  wire[0:0] mux_798_nl;
  wire[0:0] or_1145_nl;
  wire[0:0] mux_803_nl;
  wire[0:0] mux_801_nl;
  wire[0:0] mux_92_nl;
  wire[0:0] mux_802_nl;
  wire[0:0] mux_208_nl;
  wire[0:0] mux_207_nl;
  wire[0:0] mux_1687_nl;
  wire[0:0] or_2688_nl;
  wire[0:0] or_2691_nl;
  wire[0:0] mux_1689_nl;
  wire[0:0] or_2696_nl;
  wire[0:0] or_2699_nl;
  wire[0:0] mux_1692_nl;
  wire[0:0] or_2705_nl;
  wire[0:0] or_2709_nl;
  wire[0:0] mux_1694_nl;
  wire[0:0] or_2714_nl;
  wire[0:0] or_2717_nl;
  wire[0:0] mux_1697_nl;
  wire[0:0] or_2723_nl;
  wire[0:0] or_2727_nl;
  wire[0:0] mux_1700_nl;
  wire[0:0] or_2733_nl;
  wire[0:0] or_2737_nl;
  wire[0:0] mux_1704_nl;
  wire[0:0] or_2744_nl;
  wire[0:0] or_2749_nl;
  wire[0:0] mux_1707_nl;
  wire[0:0] or_2754_nl;
  wire[0:0] or_2758_nl;
  wire[0:0] mux_1711_nl;
  wire[0:0] or_2764_nl;
  wire[0:0] or_2768_nl;
  wire[0:0] mux_1715_nl;
  wire[0:0] or_2774_nl;
  wire[0:0] or_2778_nl;
  wire[0:0] mux_1720_nl;
  wire[0:0] or_2784_nl;
  wire[0:0] or_2789_nl;
  wire[0:0] mux_1727_nl;
  wire[0:0] or_2796_nl;
  wire[0:0] or_2802_nl;
  wire[0:0] mux_1734_nl;
  wire[0:0] or_2809_nl;
  wire[0:0] or_2815_nl;
  wire[0:0] mux_1743_nl;
  wire[0:0] or_2823_nl;
  wire[0:0] or_2830_nl;
  wire[0:0] mux_1286_nl;
  wire[0:0] mux_1285_nl;
  wire[0:0] mux_1284_nl;
  wire[0:0] mux_1283_nl;
  wire[0:0] mux_1415_nl;
  wire[0:0] mux_1414_nl;
  wire[0:0] mux_1413_nl;
  wire[0:0] mux_1412_nl;
  wire[0:0] mux_119_nl;
  wire[0:0] or_217_nl;
  wire[0:0] mux_121_nl;
  wire[0:0] mux_125_nl;
  wire[0:0] or_226_nl;
  wire[0:0] mux_131_nl;
  wire[0:0] or_236_nl;
  wire[0:0] or_243_nl;
  wire[0:0] mux_143_nl;
  wire[0:0] or_263_nl;
  wire[0:0] mux_150_nl;
  wire[0:0] or_270_nl;
  wire[0:0] mux_153_nl;
  wire[0:0] or_275_nl;
  wire[0:0] or_2943_nl;
  wire[0:0] or_2944_nl;
  wire[0:0] or_2945_nl;
  wire[8:0] cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_nl;
  wire[9:0] nl_cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_nl;
  wire[7:0] cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_nl;
  wire[8:0] nl_cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_nl;
  wire[8:0] cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl;
  wire[9:0] nl_cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl;
  wire[7:0] cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl;
  wire[8:0] nl_cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl;
  wire[8:0] cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl;
  wire[9:0] nl_cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl;
  wire[7:0] cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl;
  wire[8:0] nl_cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl;
  wire[8:0] cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  wire[9:0] nl_cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  wire[7:0] cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  wire[8:0] nl_cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  wire[8:0] cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl;
  wire[9:0] nl_cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl;
  wire[7:0] cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl;
  wire[8:0] nl_cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl;
  wire[8:0] cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  wire[9:0] nl_cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  wire[7:0] cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  wire[8:0] nl_cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  wire[8:0] cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  wire[9:0] nl_cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  wire[7:0] cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  wire[8:0] nl_cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  wire[8:0] cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl;
  wire[9:0] nl_cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl;
  wire[7:0] cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl;
  wire[8:0] nl_cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl;
  wire[8:0] cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl;
  wire[9:0] nl_cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl;
  wire[7:0] cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl;
  wire[8:0] nl_cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl;
  wire[8:0] cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  wire[9:0] nl_cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  wire[7:0] cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  wire[8:0] nl_cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  wire[8:0] cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  wire[9:0] nl_cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  wire[7:0] cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  wire[8:0] nl_cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  wire[8:0] cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl;
  wire[9:0] nl_cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl;
  wire[7:0] cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl;
  wire[8:0] nl_cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl;
  wire[8:0] cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  wire[9:0] nl_cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl;
  wire[7:0] cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  wire[8:0] nl_cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl;
  wire[8:0] cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl;
  wire[9:0] nl_cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl;
  wire[7:0] cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl;
  wire[8:0] nl_cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl;
  wire[8:0] cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl;
  wire[9:0] nl_cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl;
  wire[7:0] cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl;
  wire[8:0] nl_cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl;
  wire[8:0] cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_nl;
  wire[9:0] nl_cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_nl;
  wire[7:0] cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_nl;
  wire[8:0] nl_cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_nl;
  wire[8:0] cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_nl;
  wire[9:0] nl_cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_nl;
  wire[8:0] cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl;
  wire[9:0] nl_cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl;
  wire[8:0] cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl;
  wire[9:0] nl_cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl;
  wire[8:0] cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  wire[9:0] nl_cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  wire[8:0] cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl;
  wire[9:0] nl_cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl;
  wire[8:0] cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  wire[9:0] nl_cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  wire[8:0] cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  wire[9:0] nl_cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  wire[8:0] cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl;
  wire[9:0] nl_cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl;
  wire[8:0] cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl;
  wire[9:0] nl_cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl;
  wire[8:0] cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  wire[9:0] nl_cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  wire[8:0] cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  wire[9:0] nl_cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  wire[8:0] cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl;
  wire[9:0] nl_cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl;
  wire[8:0] cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  wire[9:0] nl_cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl;
  wire[8:0] cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl;
  wire[9:0] nl_cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl;
  wire[8:0] cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl;
  wire[9:0] nl_cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl;
  wire[8:0] cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_nl;
  wire[9:0] nl_cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_1_nl;
  wire[9:0] cvt_1_FpMantRNE_24U_11U_else_acc_nl;
  wire[10:0] nl_cvt_1_FpMantRNE_24U_11U_else_acc_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_47_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_48_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_32_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_1_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_13_nl;
  wire[9:0] cvt_2_FpMantRNE_24U_11U_else_acc_1_nl;
  wire[10:0] nl_cvt_2_FpMantRNE_24U_11U_else_acc_1_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_2_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_1_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_49_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_50_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_33_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_2_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_25_nl;
  wire[9:0] cvt_3_FpMantRNE_24U_11U_else_acc_1_nl;
  wire[10:0] nl_cvt_3_FpMantRNE_24U_11U_else_acc_1_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_4_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_2_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_51_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_52_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_34_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_3_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_37_nl;
  wire[9:0] cvt_4_FpMantRNE_24U_11U_else_acc_2_nl;
  wire[10:0] nl_cvt_4_FpMantRNE_24U_11U_else_acc_2_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_6_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_3_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_53_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_54_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_35_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_4_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_49_nl;
  wire[9:0] cvt_5_FpMantRNE_24U_11U_else_acc_1_nl;
  wire[10:0] nl_cvt_5_FpMantRNE_24U_11U_else_acc_1_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_8_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_4_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_55_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_56_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_36_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_5_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_61_nl;
  wire[9:0] cvt_6_FpMantRNE_24U_11U_else_acc_2_nl;
  wire[10:0] nl_cvt_6_FpMantRNE_24U_11U_else_acc_2_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_10_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_5_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_57_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_58_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_37_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_6_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_73_nl;
  wire[9:0] cvt_7_FpMantRNE_24U_11U_else_acc_2_nl;
  wire[10:0] nl_cvt_7_FpMantRNE_24U_11U_else_acc_2_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_12_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_6_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_59_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_60_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_38_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_7_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_85_nl;
  wire[9:0] cvt_8_FpMantRNE_24U_11U_else_acc_3_nl;
  wire[10:0] nl_cvt_8_FpMantRNE_24U_11U_else_acc_3_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_14_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_7_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_61_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_62_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_39_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_8_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_97_nl;
  wire[9:0] cvt_9_FpMantRNE_24U_11U_else_acc_1_nl;
  wire[10:0] nl_cvt_9_FpMantRNE_24U_11U_else_acc_1_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_16_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_8_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_63_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_64_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_40_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_9_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_109_nl;
  wire[9:0] cvt_10_FpMantRNE_24U_11U_else_acc_2_nl;
  wire[10:0] nl_cvt_10_FpMantRNE_24U_11U_else_acc_2_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_18_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_9_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_65_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_66_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_41_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_10_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_121_nl;
  wire[9:0] cvt_11_FpMantRNE_24U_11U_else_acc_2_nl;
  wire[10:0] nl_cvt_11_FpMantRNE_24U_11U_else_acc_2_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_20_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_10_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_67_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_68_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_42_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_11_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_133_nl;
  wire[9:0] cvt_12_FpMantRNE_24U_11U_else_acc_3_nl;
  wire[10:0] nl_cvt_12_FpMantRNE_24U_11U_else_acc_3_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_22_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_11_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_69_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_70_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_43_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_12_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_145_nl;
  wire[9:0] cvt_13_FpMantRNE_24U_11U_else_acc_2_nl;
  wire[10:0] nl_cvt_13_FpMantRNE_24U_11U_else_acc_2_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_24_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_12_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_71_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_72_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_44_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_13_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_157_nl;
  wire[9:0] cvt_14_FpMantRNE_24U_11U_else_acc_3_nl;
  wire[10:0] nl_cvt_14_FpMantRNE_24U_11U_else_acc_3_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_26_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_13_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_73_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_74_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_45_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_14_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_169_nl;
  wire[9:0] cvt_15_FpMantRNE_24U_11U_else_acc_3_nl;
  wire[10:0] nl_cvt_15_FpMantRNE_24U_11U_else_acc_3_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_28_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_14_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_75_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_76_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_46_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_15_nl;
  wire[9:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_181_nl;
  wire[9:0] cvt_16_FpMantRNE_24U_11U_else_acc_4_nl;
  wire[10:0] nl_cvt_16_FpMantRNE_24U_11U_else_acc_4_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_30_nl;
  wire[3:0] FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_15_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_77_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_and_78_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_47_nl;
  wire[14:0] cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_nor_2_nl;
  wire[14:0] cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_nor_7_nl;
  wire[14:0] cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_nor_7_nl;
  wire[14:0] cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl;
  wire[14:0] cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_nor_7_nl;
  wire[14:0] cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl;
  wire[14:0] cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl;
  wire[14:0] cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_nor_17_nl;
  wire[14:0] cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_nor_7_nl;
  wire[14:0] cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl;
  wire[14:0] cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl;
  wire[14:0] cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_nor_17_nl;
  wire[14:0] cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl;
  wire[14:0] cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_nor_17_nl;
  wire[14:0] cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_nor_17_nl;
  wire[14:0] cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_nor_22_nl;
  wire[11:0] cvt_1_FpFloatToInt_16U_5U_10U_if_acc_nl;
  wire[12:0] nl_cvt_1_FpFloatToInt_16U_5U_10U_if_acc_nl;
  wire[0:0] cvt_1_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_nl;
  wire[11:0] cvt_2_FpFloatToInt_16U_5U_10U_if_acc_1_nl;
  wire[12:0] nl_cvt_2_FpFloatToInt_16U_5U_10U_if_acc_1_nl;
  wire[0:0] cvt_2_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_1_nl;
  wire[10:0] cvt_3_IntSaturation_17U_8U_if_acc_1_nl;
  wire[11:0] nl_cvt_3_IntSaturation_17U_8U_if_acc_1_nl;
  wire[11:0] cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_nl;
  wire[12:0] nl_cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_nl;
  wire[0:0] cvt_3_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_1_nl;
  wire[11:0] cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  wire[12:0] nl_cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  wire[0:0] cvt_4_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl;
  wire[10:0] cvt_5_IntSaturation_17U_8U_if_acc_1_nl;
  wire[11:0] nl_cvt_5_IntSaturation_17U_8U_if_acc_1_nl;
  wire[11:0] cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_nl;
  wire[12:0] nl_cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_nl;
  wire[0:0] cvt_5_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_1_nl;
  wire[11:0] cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_nl;
  wire[12:0] nl_cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_nl;
  wire[0:0] cvt_16_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_4_nl;
  wire[11:0] cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  wire[12:0] nl_cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  wire[0:0] cvt_6_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl;
  wire[10:0] cvt_1_IntSaturation_17U_8U_if_acc_nl;
  wire[11:0] nl_cvt_1_IntSaturation_17U_8U_if_acc_nl;
  wire[11:0] cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_nl;
  wire[12:0] nl_cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_nl;
  wire[0:0] cvt_15_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_3_nl;
  wire[11:0] cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  wire[12:0] nl_cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  wire[0:0] cvt_7_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl;
  wire[11:0] cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_nl;
  wire[12:0] nl_cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_nl;
  wire[0:0] cvt_14_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_3_nl;
  wire[11:0] cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_nl;
  wire[12:0] nl_cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_nl;
  wire[0:0] cvt_8_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_3_nl;
  wire[11:0] cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  wire[12:0] nl_cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  wire[0:0] cvt_13_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl;
  wire[10:0] cvt_9_IntSaturation_17U_8U_if_acc_1_nl;
  wire[11:0] nl_cvt_9_IntSaturation_17U_8U_if_acc_1_nl;
  wire[11:0] cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_nl;
  wire[12:0] nl_cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_nl;
  wire[0:0] cvt_9_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_1_nl;
  wire[11:0] cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_nl;
  wire[12:0] nl_cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_nl;
  wire[0:0] cvt_12_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_3_nl;
  wire[11:0] cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  wire[12:0] nl_cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  wire[0:0] cvt_10_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl;
  wire[11:0] cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  wire[12:0] nl_cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_nl;
  wire[0:0] cvt_11_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_or_13_nl;
  wire[0:0] cvt_else_mux_56_nl;
  wire[0:0] cvt_else_mux_62_nl;
  wire[0:0] cvt_else_mux_59_nl;
  wire[9:0] cvt_4_FpMantRNE_17U_11U_else_acc_2_nl;
  wire[10:0] nl_cvt_4_FpMantRNE_17U_11U_else_acc_2_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_if_not_185_nl;
  wire[0:0] FpMantRNE_17U_11U_else_mux_7_nl;
  wire[0:0] or_3872_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_else_mux_10_nl;
  wire[9:0] cvt_5_FpMantRNE_17U_11U_else_acc_1_nl;
  wire[10:0] nl_cvt_5_FpMantRNE_17U_11U_else_acc_1_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_if_not_188_nl;
  wire[9:0] cvt_6_FpMantRNE_17U_11U_else_acc_2_nl;
  wire[10:0] nl_cvt_6_FpMantRNE_17U_11U_else_acc_2_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_if_not_191_nl;
  wire[0:0] FpMantRNE_17U_11U_else_mux_11_nl;
  wire[0:0] or_3891_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_else_mux_16_nl;
  wire[9:0] cvt_7_FpMantRNE_17U_11U_else_acc_2_nl;
  wire[10:0] nl_cvt_7_FpMantRNE_17U_11U_else_acc_2_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_if_not_194_nl;
  wire[0:0] FpMantRNE_17U_11U_else_mux_13_nl;
  wire[0:0] or_3900_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_else_mux_19_nl;
  wire[9:0] cvt_8_FpMantRNE_17U_11U_else_acc_3_nl;
  wire[10:0] nl_cvt_8_FpMantRNE_17U_11U_else_acc_3_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_if_not_197_nl;
  wire[0:0] FpMantRNE_17U_11U_else_mux_15_nl;
  wire[0:0] or_3911_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_else_mux_22_nl;
  wire[9:0] cvt_10_FpMantRNE_17U_11U_else_acc_2_nl;
  wire[10:0] nl_cvt_10_FpMantRNE_17U_11U_else_acc_2_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_if_not_203_nl;
  wire[0:0] FpMantRNE_17U_11U_else_mux_19_nl;
  wire[0:0] or_3932_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_else_mux_28_nl;
  wire[9:0] cvt_11_FpMantRNE_17U_11U_else_acc_2_nl;
  wire[10:0] nl_cvt_11_FpMantRNE_17U_11U_else_acc_2_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_if_not_206_nl;
  wire[0:0] FpMantRNE_17U_11U_else_mux_21_nl;
  wire[0:0] or_3942_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_else_mux_31_nl;
  wire[9:0] cvt_12_FpMantRNE_17U_11U_else_acc_3_nl;
  wire[10:0] nl_cvt_12_FpMantRNE_17U_11U_else_acc_3_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_if_not_209_nl;
  wire[0:0] FpMantRNE_17U_11U_else_mux_23_nl;
  wire[0:0] or_3953_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_else_mux_34_nl;
  wire[9:0] cvt_13_FpMantRNE_17U_11U_else_acc_2_nl;
  wire[10:0] nl_cvt_13_FpMantRNE_17U_11U_else_acc_2_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_if_not_212_nl;
  wire[0:0] FpMantRNE_17U_11U_else_mux_25_nl;
  wire[0:0] or_3965_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_else_mux_37_nl;
  wire[9:0] cvt_14_FpMantRNE_17U_11U_else_acc_3_nl;
  wire[10:0] nl_cvt_14_FpMantRNE_17U_11U_else_acc_3_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_if_not_215_nl;
  wire[0:0] FpMantRNE_17U_11U_else_mux_27_nl;
  wire[0:0] or_3977_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_else_mux_40_nl;
  wire[9:0] cvt_15_FpMantRNE_17U_11U_else_acc_3_nl;
  wire[10:0] nl_cvt_15_FpMantRNE_17U_11U_else_acc_3_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_if_not_218_nl;
  wire[0:0] FpMantRNE_17U_11U_else_mux_29_nl;
  wire[0:0] or_3989_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_else_mux_43_nl;
  wire[9:0] cvt_16_FpMantRNE_17U_11U_else_acc_4_nl;
  wire[10:0] nl_cvt_16_FpMantRNE_17U_11U_else_acc_4_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_if_not_221_nl;
  wire[0:0] FpMantRNE_17U_11U_else_mux_31_nl;
  wire[0:0] or_3999_nl;
  wire[0:0] FpIntToFloat_17U_5U_10U_else_mux_46_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_32_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_33_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_34_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_35_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_36_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_37_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_38_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_39_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_40_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_41_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_42_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_43_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_44_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_45_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_46_nl;
  wire[0:0] FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_47_nl;
  wire[17:0] cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl;
  wire[18:0] nl_cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl;
  wire[17:0] cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  wire[18:0] nl_cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  wire[17:0] cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl;
  wire[18:0] nl_cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl;
  wire[17:0] cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  wire[18:0] nl_cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  wire[17:0] cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl;
  wire[18:0] nl_cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl;
  wire[17:0] cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  wire[18:0] nl_cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  wire[17:0] cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl;
  wire[18:0] nl_cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl;
  wire[17:0] cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  wire[18:0] nl_cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  wire[17:0] cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl;
  wire[18:0] nl_cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl;
  wire[17:0] cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  wire[18:0] nl_cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  wire[17:0] cvt_14_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl;
  wire[18:0] nl_cvt_14_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl;
  wire[17:0] cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl;
  wire[18:0] nl_cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl;
  wire[17:0] cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl;
  wire[18:0] nl_cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl;
  wire[17:0] cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  wire[18:0] nl_cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl;
  wire[17:0] cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl;
  wire[18:0] nl_cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl;
  wire[17:0] cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl;
  wire[18:0] nl_cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl;
  wire[2:0] cvt_1_IntSaturation_17U_16U_if_acc_nl;
  wire[3:0] nl_cvt_1_IntSaturation_17U_16U_if_acc_nl;
  wire[2:0] cvt_2_IntSaturation_17U_16U_if_acc_1_nl;
  wire[3:0] nl_cvt_2_IntSaturation_17U_16U_if_acc_1_nl;
  wire[0:0] cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_and_2_nl;
  wire[2:0] cvt_3_IntSaturation_17U_16U_if_acc_1_nl;
  wire[3:0] nl_cvt_3_IntSaturation_17U_16U_if_acc_1_nl;
  wire[2:0] cvt_4_IntSaturation_17U_16U_if_acc_2_nl;
  wire[3:0] nl_cvt_4_IntSaturation_17U_16U_if_acc_2_nl;
  wire[0:0] cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl;
  wire[0:0] cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_and_2_nl;
  wire[2:0] cvt_5_IntSaturation_17U_16U_if_acc_1_nl;
  wire[3:0] nl_cvt_5_IntSaturation_17U_16U_if_acc_1_nl;
  wire[2:0] cvt_6_IntSaturation_17U_16U_if_acc_2_nl;
  wire[3:0] nl_cvt_6_IntSaturation_17U_16U_if_acc_2_nl;
  wire[0:0] cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl;
  wire[2:0] cvt_7_IntSaturation_17U_16U_if_acc_2_nl;
  wire[3:0] nl_cvt_7_IntSaturation_17U_16U_if_acc_2_nl;
  wire[2:0] cvt_8_IntSaturation_17U_16U_if_acc_3_nl;
  wire[3:0] nl_cvt_8_IntSaturation_17U_16U_if_acc_3_nl;
  wire[0:0] cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_and_6_nl;
  wire[0:0] cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl;
  wire[0:0] cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_and_2_nl;
  wire[2:0] cvt_9_IntSaturation_17U_16U_if_acc_1_nl;
  wire[3:0] nl_cvt_9_IntSaturation_17U_16U_if_acc_1_nl;
  wire[2:0] cvt_10_IntSaturation_17U_16U_if_acc_2_nl;
  wire[3:0] nl_cvt_10_IntSaturation_17U_16U_if_acc_2_nl;
  wire[0:0] cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl;
  wire[2:0] cvt_11_IntSaturation_17U_16U_if_acc_2_nl;
  wire[3:0] nl_cvt_11_IntSaturation_17U_16U_if_acc_2_nl;
  wire[2:0] cvt_12_IntSaturation_17U_16U_if_acc_3_nl;
  wire[3:0] nl_cvt_12_IntSaturation_17U_16U_if_acc_3_nl;
  wire[0:0] cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_and_6_nl;
  wire[0:0] cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl;
  wire[2:0] cvt_13_IntSaturation_17U_16U_if_acc_2_nl;
  wire[3:0] nl_cvt_13_IntSaturation_17U_16U_if_acc_2_nl;
  wire[2:0] cvt_14_IntSaturation_17U_16U_if_acc_3_nl;
  wire[3:0] nl_cvt_14_IntSaturation_17U_16U_if_acc_3_nl;
  wire[0:0] cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_and_6_nl;
  wire[2:0] cvt_15_IntSaturation_17U_16U_if_acc_3_nl;
  wire[3:0] nl_cvt_15_IntSaturation_17U_16U_if_acc_3_nl;
  wire[2:0] cvt_16_IntSaturation_17U_16U_if_acc_4_nl;
  wire[3:0] nl_cvt_16_IntSaturation_17U_16U_if_acc_4_nl;
  wire[0:0] cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_and_8_nl;
  wire[0:0] cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_and_6_nl;
  wire[0:0] cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl;
  wire[0:0] cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_and_2_nl;
  wire[0:0] cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_and_nl;
  wire[0:0] cvt_1_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_nl;
  wire[23:0] cvt_1_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_2_nl;
  wire[0:0] cvt_2_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_2_nl;
  wire[23:0] cvt_2_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_7_nl;
  wire[0:0] cvt_3_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_2_nl;
  wire[23:0] cvt_3_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_7_nl;
  wire[0:0] cvt_4_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl;
  wire[23:0] cvt_4_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl;
  wire[0:0] cvt_5_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_2_nl;
  wire[23:0] cvt_5_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_7_nl;
  wire[0:0] cvt_6_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl;
  wire[23:0] cvt_6_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl;
  wire[0:0] cvt_7_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl;
  wire[23:0] cvt_7_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl;
  wire[0:0] cvt_8_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_6_nl;
  wire[23:0] cvt_8_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_17_nl;
  wire[0:0] cvt_9_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_2_nl;
  wire[23:0] cvt_9_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_7_nl;
  wire[0:0] cvt_10_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl;
  wire[23:0] cvt_10_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl;
  wire[0:0] cvt_11_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl;
  wire[23:0] cvt_11_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl;
  wire[0:0] cvt_12_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_6_nl;
  wire[23:0] cvt_12_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_17_nl;
  wire[0:0] cvt_13_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl;
  wire[23:0] cvt_13_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl;
  wire[0:0] cvt_14_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_6_nl;
  wire[23:0] cvt_14_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_17_nl;
  wire[0:0] cvt_15_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_6_nl;
  wire[23:0] cvt_15_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_17_nl;
  wire[0:0] cvt_16_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_8_nl;
  wire[23:0] cvt_16_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_22_nl;
  wire[4:0] cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_1_nl;
  wire[5:0] nl_cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_1_nl;
  wire[4:0] cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl;
  wire[5:0] nl_cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl;
  wire[4:0] cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl;
  wire[5:0] nl_cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl;
  wire[4:0] cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  wire[5:0] nl_cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  wire[4:0] cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl;
  wire[5:0] nl_cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl;
  wire[4:0] cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  wire[5:0] nl_cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  wire[4:0] cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  wire[5:0] nl_cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  wire[4:0] cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl;
  wire[5:0] nl_cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl;
  wire[4:0] cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl;
  wire[5:0] nl_cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl;
  wire[4:0] cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  wire[5:0] nl_cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  wire[4:0] cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  wire[5:0] nl_cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  wire[4:0] cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl;
  wire[5:0] nl_cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl;
  wire[4:0] cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  wire[5:0] nl_cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl;
  wire[4:0] cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl;
  wire[5:0] nl_cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl;
  wire[4:0] cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl;
  wire[5:0] nl_cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl;
  wire[4:0] cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_8_nl;
  wire[5:0] nl_cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_8_nl;
  wire[10:0] cvt_1_IntSaturation_17U_8U_else_if_acc_nl;
  wire[11:0] nl_cvt_1_IntSaturation_17U_8U_else_if_acc_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_nor_nl;
  wire[0:0] IntSaturation_17U_8U_and_1_nl;
  wire[10:0] cvt_2_IntSaturation_17U_8U_else_if_acc_1_nl;
  wire[11:0] nl_cvt_2_IntSaturation_17U_8U_else_if_acc_1_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_nor_1_nl;
  wire[0:0] IntSaturation_17U_8U_and_3_nl;
  wire[10:0] cvt_3_IntSaturation_17U_8U_else_if_acc_1_nl;
  wire[11:0] nl_cvt_3_IntSaturation_17U_8U_else_if_acc_1_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_nor_2_nl;
  wire[0:0] IntSaturation_17U_8U_and_5_nl;
  wire[10:0] cvt_4_IntSaturation_17U_8U_else_if_acc_2_nl;
  wire[11:0] nl_cvt_4_IntSaturation_17U_8U_else_if_acc_2_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_nor_3_nl;
  wire[0:0] IntSaturation_17U_8U_and_7_nl;
  wire[10:0] cvt_5_IntSaturation_17U_8U_else_if_acc_1_nl;
  wire[11:0] nl_cvt_5_IntSaturation_17U_8U_else_if_acc_1_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_nor_4_nl;
  wire[0:0] IntSaturation_17U_8U_and_9_nl;
  wire[10:0] cvt_6_IntSaturation_17U_8U_else_if_acc_2_nl;
  wire[11:0] nl_cvt_6_IntSaturation_17U_8U_else_if_acc_2_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_nor_5_nl;
  wire[0:0] IntSaturation_17U_8U_and_11_nl;
  wire[10:0] cvt_7_IntSaturation_17U_8U_else_if_acc_2_nl;
  wire[11:0] nl_cvt_7_IntSaturation_17U_8U_else_if_acc_2_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_nor_6_nl;
  wire[0:0] IntSaturation_17U_8U_and_13_nl;
  wire[10:0] cvt_8_IntSaturation_17U_8U_else_if_acc_3_nl;
  wire[11:0] nl_cvt_8_IntSaturation_17U_8U_else_if_acc_3_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_nor_7_nl;
  wire[0:0] IntSaturation_17U_8U_and_15_nl;
  wire[10:0] cvt_9_IntSaturation_17U_8U_else_if_acc_1_nl;
  wire[11:0] nl_cvt_9_IntSaturation_17U_8U_else_if_acc_1_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_nor_8_nl;
  wire[0:0] IntSaturation_17U_8U_and_17_nl;
  wire[10:0] cvt_10_IntSaturation_17U_8U_else_if_acc_2_nl;
  wire[11:0] nl_cvt_10_IntSaturation_17U_8U_else_if_acc_2_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_nor_9_nl;
  wire[0:0] IntSaturation_17U_8U_and_19_nl;
  wire[10:0] cvt_11_IntSaturation_17U_8U_else_if_acc_2_nl;
  wire[11:0] nl_cvt_11_IntSaturation_17U_8U_else_if_acc_2_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_nor_10_nl;
  wire[0:0] IntSaturation_17U_8U_and_21_nl;
  wire[10:0] cvt_12_IntSaturation_17U_8U_else_if_acc_3_nl;
  wire[11:0] nl_cvt_12_IntSaturation_17U_8U_else_if_acc_3_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_nor_11_nl;
  wire[0:0] IntSaturation_17U_8U_and_23_nl;
  wire[10:0] cvt_13_IntSaturation_17U_8U_else_if_acc_2_nl;
  wire[11:0] nl_cvt_13_IntSaturation_17U_8U_else_if_acc_2_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_nor_12_nl;
  wire[0:0] IntSaturation_17U_8U_and_25_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_nor_13_nl;
  wire[0:0] IntSaturation_17U_8U_and_27_nl;
  wire[10:0] cvt_15_IntSaturation_17U_8U_else_if_acc_3_nl;
  wire[11:0] nl_cvt_15_IntSaturation_17U_8U_else_if_acc_3_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_nor_14_nl;
  wire[0:0] IntSaturation_17U_8U_and_29_nl;
  wire[10:0] cvt_16_IntSaturation_17U_8U_else_if_acc_4_nl;
  wire[11:0] nl_cvt_16_IntSaturation_17U_8U_else_if_acc_4_nl;
  wire[0:0] IntSaturation_17U_8U_IntSaturation_17U_8U_nor_15_nl;
  wire[0:0] IntSaturation_17U_8U_and_31_nl;
  wire[10:0] cvt_14_IntSaturation_17U_8U_else_if_acc_3_nl;
  wire[11:0] nl_cvt_14_IntSaturation_17U_8U_else_if_acc_3_nl;
  wire[0:0] cvt_1_FpMantDecShiftRight_23U_8U_10U_carry_and_nl;
  wire[22:0] cvt_1_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl;
  wire[23:0] nl_cvt_1_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl;
  wire[0:0] cvt_2_FpMantDecShiftRight_23U_8U_10U_carry_and_1_nl;
  wire[22:0] cvt_2_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl;
  wire[23:0] nl_cvt_2_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl;
  wire[0:0] cvt_3_FpMantDecShiftRight_23U_8U_10U_carry_and_1_nl;
  wire[22:0] cvt_3_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl;
  wire[23:0] nl_cvt_3_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl;
  wire[0:0] cvt_4_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl;
  wire[22:0] cvt_4_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  wire[23:0] nl_cvt_4_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  wire[0:0] cvt_5_FpMantDecShiftRight_23U_8U_10U_carry_and_1_nl;
  wire[22:0] cvt_5_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl;
  wire[23:0] nl_cvt_5_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl;
  wire[0:0] cvt_6_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl;
  wire[22:0] cvt_6_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  wire[23:0] nl_cvt_6_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  wire[0:0] cvt_7_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl;
  wire[22:0] cvt_7_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  wire[23:0] nl_cvt_7_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  wire[0:0] cvt_8_FpMantDecShiftRight_23U_8U_10U_carry_and_3_nl;
  wire[22:0] cvt_8_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl;
  wire[23:0] nl_cvt_8_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl;
  wire[0:0] cvt_9_FpMantDecShiftRight_23U_8U_10U_carry_and_1_nl;
  wire[22:0] cvt_9_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl;
  wire[23:0] nl_cvt_9_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl;
  wire[0:0] cvt_10_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl;
  wire[22:0] cvt_10_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  wire[23:0] nl_cvt_10_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  wire[0:0] cvt_11_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl;
  wire[22:0] cvt_11_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  wire[23:0] nl_cvt_11_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  wire[0:0] cvt_12_FpMantDecShiftRight_23U_8U_10U_carry_and_3_nl;
  wire[22:0] cvt_12_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl;
  wire[23:0] nl_cvt_12_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl;
  wire[0:0] cvt_13_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl;
  wire[22:0] cvt_13_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  wire[23:0] nl_cvt_13_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl;
  wire[0:0] cvt_14_FpMantDecShiftRight_23U_8U_10U_carry_and_3_nl;
  wire[22:0] cvt_14_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl;
  wire[23:0] nl_cvt_14_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl;
  wire[0:0] cvt_15_FpMantDecShiftRight_23U_8U_10U_carry_and_3_nl;
  wire[22:0] cvt_15_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl;
  wire[23:0] nl_cvt_15_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl;
  wire[0:0] cvt_16_FpMantDecShiftRight_23U_8U_10U_carry_and_4_nl;
  wire[22:0] cvt_16_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_4_nl;
  wire[23:0] nl_cvt_16_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_4_nl;
  wire[2:0] cvt_1_IntSaturation_17U_16U_else_if_acc_nl;
  wire[3:0] nl_cvt_1_IntSaturation_17U_16U_else_if_acc_nl;
  wire[2:0] cvt_2_IntSaturation_17U_16U_else_if_acc_1_nl;
  wire[3:0] nl_cvt_2_IntSaturation_17U_16U_else_if_acc_1_nl;
  wire[2:0] cvt_3_IntSaturation_17U_16U_else_if_acc_1_nl;
  wire[3:0] nl_cvt_3_IntSaturation_17U_16U_else_if_acc_1_nl;
  wire[2:0] cvt_4_IntSaturation_17U_16U_else_if_acc_2_nl;
  wire[3:0] nl_cvt_4_IntSaturation_17U_16U_else_if_acc_2_nl;
  wire[2:0] cvt_5_IntSaturation_17U_16U_else_if_acc_1_nl;
  wire[3:0] nl_cvt_5_IntSaturation_17U_16U_else_if_acc_1_nl;
  wire[2:0] cvt_6_IntSaturation_17U_16U_else_if_acc_2_nl;
  wire[3:0] nl_cvt_6_IntSaturation_17U_16U_else_if_acc_2_nl;
  wire[2:0] cvt_7_IntSaturation_17U_16U_else_if_acc_2_nl;
  wire[3:0] nl_cvt_7_IntSaturation_17U_16U_else_if_acc_2_nl;
  wire[2:0] cvt_8_IntSaturation_17U_16U_else_if_acc_3_nl;
  wire[3:0] nl_cvt_8_IntSaturation_17U_16U_else_if_acc_3_nl;
  wire[2:0] cvt_9_IntSaturation_17U_16U_else_if_acc_1_nl;
  wire[3:0] nl_cvt_9_IntSaturation_17U_16U_else_if_acc_1_nl;
  wire[2:0] cvt_10_IntSaturation_17U_16U_else_if_acc_2_nl;
  wire[3:0] nl_cvt_10_IntSaturation_17U_16U_else_if_acc_2_nl;
  wire[2:0] cvt_11_IntSaturation_17U_16U_else_if_acc_2_nl;
  wire[3:0] nl_cvt_11_IntSaturation_17U_16U_else_if_acc_2_nl;
  wire[2:0] cvt_12_IntSaturation_17U_16U_else_if_acc_3_nl;
  wire[3:0] nl_cvt_12_IntSaturation_17U_16U_else_if_acc_3_nl;
  wire[2:0] cvt_13_IntSaturation_17U_16U_else_if_acc_2_nl;
  wire[3:0] nl_cvt_13_IntSaturation_17U_16U_else_if_acc_2_nl;
  wire[2:0] cvt_15_IntSaturation_17U_16U_else_if_acc_3_nl;
  wire[3:0] nl_cvt_15_IntSaturation_17U_16U_else_if_acc_3_nl;
  wire[2:0] cvt_16_IntSaturation_17U_16U_else_if_acc_4_nl;
  wire[3:0] nl_cvt_16_IntSaturation_17U_16U_else_if_acc_4_nl;
  wire[2:0] cvt_14_IntSaturation_17U_16U_else_if_acc_3_nl;
  wire[3:0] nl_cvt_14_IntSaturation_17U_16U_else_if_acc_3_nl;
  wire[0:0] or_23_nl;
  wire[0:0] or_86_nl;
  wire[0:0] mux_109_nl;
  wire[0:0] nor_2056_nl;
  wire[0:0] nor_2055_nl;
  wire[0:0] nor_2054_nl;
  wire[0:0] nor_2052_nl;
  wire[0:0] mux_148_nl;
  wire[0:0] nor_2050_nl;
  wire[0:0] nor_2049_nl;
  wire[0:0] nand_nl;
  wire[0:0] mux_188_nl;
  wire[0:0] nor_2029_nl;
  wire[0:0] or_378_nl;
  wire[0:0] nor_48_nl;
  wire[0:0] nor_2027_nl;
  wire[0:0] nor_2028_nl;
  wire[0:0] nor_2022_nl;
  wire[0:0] nor_2021_nl;
  wire[0:0] mux_244_nl;
  wire[0:0] or_429_nl;
  wire[0:0] or_431_nl;
  wire[0:0] or_434_nl;
  wire[0:0] or_448_nl;
  wire[0:0] and_152_nl;
  wire[0:0] mux_250_nl;
  wire[0:0] and_153_nl;
  wire[0:0] or_445_nl;
  wire[0:0] mux_252_nl;
  wire[0:0] nor_2015_nl;
  wire[0:0] nor_2013_nl;
  wire[0:0] nor_2007_nl;
  wire[0:0] nor_2009_nl;
  wire[0:0] nor_1995_nl;
  wire[0:0] nor_1997_nl;
  wire[0:0] nor_1988_nl;
  wire[0:0] nor_1987_nl;
  wire[0:0] and_167_nl;
  wire[0:0] or_520_nl;
  wire[0:0] nor_1983_nl;
  wire[0:0] mux_308_nl;
  wire[0:0] mux_310_nl;
  wire[0:0] mux_312_nl;
  wire[0:0] nor_1975_nl;
  wire[0:0] nor_1977_nl;
  wire[0:0] nor_1974_nl;
  wire[0:0] nor_1964_nl;
  wire[0:0] nor_1966_nl;
  wire[0:0] nor_1959_nl;
  wire[0:0] nor_1955_nl;
  wire[0:0] and_176_nl;
  wire[0:0] or_599_nl;
  wire[0:0] mux_369_nl;
  wire[0:0] nor_1942_nl;
  wire[0:0] nor_1944_nl;
  wire[0:0] nor_1935_nl;
  wire[0:0] and_181_nl;
  wire[0:0] or_645_nl;
  wire[0:0] mux_404_nl;
  wire[0:0] nor_1922_nl;
  wire[0:0] nor_1924_nl;
  wire[0:0] nor_1919_nl;
  wire[0:0] nor_1912_nl;
  wire[0:0] nor_1915_nl;
  wire[0:0] and_184_nl;
  wire[0:0] or_690_nl;
  wire[0:0] nor_1911_nl;
  wire[0:0] nor_1906_nl;
  wire[0:0] nor_1901_nl;
  wire[0:0] nor_1902_nl;
  wire[0:0] nor_1892_nl;
  wire[0:0] nor_1894_nl;
  wire[0:0] nor_1891_nl;
  wire[0:0] nor_1882_nl;
  wire[0:0] nor_1884_nl;
  wire[0:0] nor_1872_nl;
  wire[0:0] mux_486_nl;
  wire[0:0] and_2218_nl;
  wire[0:0] or_784_nl;
  wire[0:0] mux_500_nl;
  wire[0:0] or_795_nl;
  wire[0:0] nor_1858_nl;
  wire[0:0] nor_1860_nl;
  wire[0:0] nor_1851_nl;
  wire[0:0] mux_524_nl;
  wire[0:0] and_2214_nl;
  wire[0:0] or_828_nl;
  wire[0:0] mux_540_nl;
  wire[0:0] mux_538_nl;
  wire[0:0] nor_1838_nl;
  wire[0:0] nor_1840_nl;
  wire[0:0] nor_1828_nl;
  wire[0:0] and_2210_nl;
  wire[0:0] or_871_nl;
  wire[0:0] nor_1827_nl;
  wire[0:0] mux_576_nl;
  wire[0:0] and_2209_nl;
  wire[0:0] nor_1815_nl;
  wire[0:0] nor_1816_nl;
  wire[0:0] nor_1817_nl;
  wire[0:0] or_894_nl;
  wire[0:0] or_898_nl;
  wire[0:0] and_2208_nl;
  wire[0:0] nor_1810_nl;
  wire[0:0] nor_1807_nl;
  wire[0:0] or_921_nl;
  wire[0:0] nor_1803_nl;
  wire[0:0] nor_1804_nl;
  wire[0:0] mux_611_nl;
  wire[0:0] nor_1795_nl;
  wire[0:0] nor_1796_nl;
  wire[0:0] nor_1787_nl;
  wire[0:0] nor_1789_nl;
  wire[0:0] nor_1780_nl;
  wire[0:0] mux_637_nl;
  wire[0:0] and_2202_nl;
  wire[0:0] nor_1774_nl;
  wire[0:0] nor_1775_nl;
  wire[0:0] nor_1776_nl;
  wire[0:0] nor_1764_nl;
  wire[0:0] nor_1766_nl;
  wire[0:0] nor_1762_nl;
  wire[0:0] or_1015_nl;
  wire[0:0] nor_1748_nl;
  wire[0:0] nor_1749_nl;
  wire[0:0] nor_1750_nl;
  wire[0:0] mux_691_nl;
  wire[0:0] nor_1738_nl;
  wire[0:0] nor_1739_nl;
  wire[0:0] nor_1740_nl;
  wire[0:0] nor_1728_nl;
  wire[0:0] nor_1730_nl;
  wire[0:0] nor_1718_nl;
  wire[0:0] nor_1719_nl;
  wire[0:0] or_1072_nl;
  wire[0:0] nor_1711_nl;
  wire[0:0] nor_1712_nl;
  wire[0:0] nor_1713_nl;
  wire[0:0] nor_1714_nl;
  wire[0:0] mux_738_nl;
  wire[0:0] nor_1699_nl;
  wire[0:0] nor_1700_nl;
  wire[0:0] nor_1701_nl;
  wire[0:0] nor_1702_nl;
  wire[0:0] nor_1687_nl;
  wire[0:0] nor_1689_nl;
  wire[0:0] nor_1685_nl;
  wire[0:0] nor_1686_nl;
  wire[0:0] mux_969_nl;
  wire[0:0] nor_1545_nl;
  wire[0:0] nor_1534_nl;
  wire[0:0] nor_1535_nl;
  wire[0:0] mux_1014_nl;
  wire[0:0] mux_1013_nl;
  wire[0:0] and_2247_nl;
  wire[0:0] nor_208_nl;
  wire[0:0] or_1644_nl;
  wire[0:0] nor_1487_nl;
  wire[0:0] or_1643_nl;
  wire[0:0] mux_1040_nl;
  wire[0:0] mux_1042_nl;
  wire[0:0] mux_1046_nl;
  wire[0:0] mux_1048_nl;
  wire[0:0] mux_1073_nl;
  wire[0:0] mux_1072_nl;
  wire[0:0] nor_1464_nl;
  wire[0:0] nor_250_nl;
  wire[0:0] mux_1087_nl;
  wire[0:0] mux_1086_nl;
  wire[0:0] nor_1455_nl;
  wire[0:0] or_1745_nl;
  wire[0:0] mux_976_nl;
  wire[0:0] or_1774_nl;
  wire[0:0] nor_1446_nl;
  wire[0:0] or_1773_nl;
  wire[0:0] mux_1102_nl;
  wire[0:0] mux_1104_nl;
  wire[0:0] mux_1108_nl;
  wire[0:0] mux_1110_nl;
  wire[0:0] mux_1151_nl;
  wire[0:0] nor_1387_nl;
  wire[0:0] nor_1388_nl;
  wire[0:0] nor_1371_nl;
  wire[0:0] nor_1372_nl;
  wire[0:0] nor_1373_nl;
  wire[0:0] mux_1269_nl;
  wire[0:0] mux_1275_nl;
  wire[0:0] mux_1274_nl;
  wire[0:0] mux_1273_nl;
  wire[0:0] mux_1272_nl;
  wire[0:0] mux_1271_nl;
  wire[0:0] mux_1281_nl;
  wire[0:0] mux_1325_nl;
  wire[0:0] mux_1331_nl;
  wire[0:0] mux_1330_nl;
  wire[0:0] mux_1329_nl;
  wire[0:0] mux_1328_nl;
  wire[0:0] mux_1327_nl;
  wire[0:0] mux_1338_nl;
  wire[0:0] mux_1340_nl;
  wire[0:0] mux_1408_nl;
  wire[0:0] mux_1407_nl;
  wire[0:0] mux_1406_nl;
  wire[0:0] mux_1405_nl;
  wire[0:0] or_2232_nl;
  wire[0:0] mux_1418_nl;
  wire[0:0] mux_1417_nl;
  wire[0:0] mux_1416_nl;
  wire[0:0] or_2245_nl;
  wire[0:0] or_2246_nl;
  wire[0:0] mux_1434_nl;
  wire[0:0] mux_1433_nl;
  wire[0:0] mux_1432_nl;
  wire[0:0] mux_1431_nl;
  wire[0:0] mux_1430_nl;
  wire[0:0] and_306_nl;
  wire[0:0] or_2306_nl;
  wire[0:0] nand_230_nl;
  wire[0:0] nor_1063_nl;
  wire[0:0] mux_1839_nl;
  wire[0:0] mux_1841_nl;
  wire[0:0] nor_1053_nl;
  wire[0:0] nor_1025_nl;
  wire[0:0] mux_1836_nl;
  wire[0:0] and_2158_nl;
  wire[0:0] mux_1846_nl;
  wire[0:0] and_2157_nl;
  wire[0:0] mux_1876_nl;
  wire[0:0] and_2155_nl;
  wire[0:0] mux_1903_nl;
  wire[0:0] and_2152_nl;
  wire[0:0] mux_1927_nl;
  wire[0:0] and_2150_nl;
  wire[0:0] mux_1940_nl;
  wire[0:0] and_2148_nl;
  wire[0:0] mux_1943_nl;
  wire[0:0] and_2147_nl;
  wire[0:0] mux_1953_nl;
  wire[0:0] and_2146_nl;
  wire[0:0] mux_1964_nl;
  wire[0:0] and_2145_nl;
  wire[0:0] mux_2205_nl;
  wire[0:0] mux_2204_nl;
  wire[0:0] mux_2203_nl;
  wire[0:0] mux_2201_nl;
  wire[0:0] mux_2200_nl;
  wire[0:0] mux_2202_nl;
  wire[0:0] or_4667_nl;
  wire[0:0] mux_2208_nl;
  wire[0:0] mux_2207_nl;
  wire[0:0] or_4675_nl;
  wire[0:0] mux_2299_nl;
  wire[0:0] mux_2303_nl;
  wire[0:0] mux_2305_nl;
  wire[0:0] mux_2309_nl;
  wire[0:0] mux_2311_nl;
  wire[0:0] mux_2315_nl;
  wire[0:0] mux_2317_nl;
  wire[0:0] mux_2322_nl;
  wire[0:0] mux_2324_nl;
  wire[0:0] mux_2329_nl;
  wire[0:0] mux_2333_nl;
  wire[0:0] mux_2335_nl;
  wire[0:0] mux_2341_nl;
  wire[0:0] mux_2346_nl;
  wire[0:0] mux_2350_nl;
  wire[0:0] mux_2352_nl;
  wire[0:0] mux_2356_nl;
  wire[0:0] mux_2358_nl;
// Interconnect Declarations for Component Instantiations
  wire [111:0] nl_cvt_2_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg_a;
  assign nl_cvt_2_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg_a = {IntMulExt_33U_16U_49U_return_2_sva_2
      , 63'b0};
  wire [111:0] nl_cvt_4_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a;
  assign nl_cvt_4_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a = {IntMulExt_33U_16U_49U_return_4_sva_1
      , 63'b0};
  wire [111:0] nl_cvt_3_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg_a;
  assign nl_cvt_3_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg_a = {IntMulExt_33U_16U_49U_return_3_sva_2
      , 63'b0};
  wire [111:0] nl_cvt_6_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a;
  assign nl_cvt_6_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a = {IntMulExt_33U_16U_49U_return_6_sva_1
      , 63'b0};
  wire [111:0] nl_cvt_8_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg_a;
  assign nl_cvt_8_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg_a = {IntMulExt_33U_16U_49U_return_8_sva_1
      , 63'b0};
  wire [111:0] nl_cvt_7_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a;
  assign nl_cvt_7_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a = {IntMulExt_33U_16U_49U_return_7_sva_1
      , 63'b0};
  wire [111:0] nl_cvt_5_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg_a;
  assign nl_cvt_5_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg_a = {IntMulExt_33U_16U_49U_return_5_sva_2
      , 63'b0};
  wire [111:0] nl_cvt_10_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a;
  assign nl_cvt_10_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a = {IntMulExt_33U_16U_49U_return_10_sva_1
      , 63'b0};
  wire [111:0] nl_cvt_12_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg_a;
  assign nl_cvt_12_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg_a = {IntMulExt_33U_16U_49U_return_12_sva_1
      , 63'b0};
  wire [111:0] nl_cvt_11_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a;
  assign nl_cvt_11_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a = {IntMulExt_33U_16U_49U_return_11_sva_1
      , 63'b0};
  wire [111:0] nl_cvt_14_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg_a;
  assign nl_cvt_14_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg_a = {IntMulExt_33U_16U_49U_return_14_sva_1
      , 63'b0};
  wire [111:0] nl_cvt_16_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_4_rg_a;
  assign nl_cvt_16_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_4_rg_a = {IntMulExt_33U_16U_49U_return_sva_1
      , 63'b0};
  wire [111:0] nl_cvt_15_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg_a;
  assign nl_cvt_15_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg_a = {IntMulExt_33U_16U_49U_return_15_sva_1
      , 63'b0};
  wire [111:0] nl_cvt_13_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a;
  assign nl_cvt_13_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a = {IntMulExt_33U_16U_49U_return_13_sva_1
      , 63'b0};
  wire [111:0] nl_cvt_9_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg_a;
  assign nl_cvt_9_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg_a = {IntMulExt_33U_16U_49U_return_9_sva_2
      , 63'b0};
  wire [111:0] nl_cvt_1_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_rg_a;
  assign nl_cvt_1_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_rg_a = {IntMulExt_33U_16U_49U_return_1_sva_2
      , 63'b0};
  wire [41:0] nl_cvt_1_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_rg_a;
  assign nl_cvt_1_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_rg_a = {1'b1
      , FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_1_lpi_1_dfm_8 , 31'b0};
  wire [5:0] nl_cvt_1_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_rg_s;
  assign nl_cvt_1_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_rg_s = {cvt_1_FpFloatToInt_16U_5U_10U_shift_acc_itm_2
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_9_3_0_1[0]))};
  wire [41:0] nl_cvt_2_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_a;
  assign nl_cvt_2_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_a = {1'b1
      , FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_2_lpi_1_dfm_8 , 31'b0};
  wire [5:0] nl_cvt_2_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s;
  assign nl_cvt_2_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s = {cvt_2_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_9_3_0_1[0]))};
  wire [41:0] nl_cvt_3_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_a;
  assign nl_cvt_3_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_a = {1'b1
      , FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_3_lpi_1_dfm_8 , 31'b0};
  wire [5:0] nl_cvt_3_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s;
  assign nl_cvt_3_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s = {cvt_3_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_9_3_0_1[0]))};
  wire [41:0] nl_cvt_4_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a;
  assign nl_cvt_4_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a = {1'b1
      , FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_4_lpi_1_dfm_8 , 31'b0};
  wire [5:0] nl_cvt_4_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s;
  assign nl_cvt_4_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s = {cvt_4_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_9_3_0_1[0]))};
  wire [41:0] nl_cvt_5_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_a;
  assign nl_cvt_5_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_a = {1'b1
      , FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_5_lpi_1_dfm_8 , 31'b0};
  wire [5:0] nl_cvt_5_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s;
  assign nl_cvt_5_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s = {cvt_5_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_9_3_0_1[0]))};
  wire [41:0] nl_cvt_6_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a;
  assign nl_cvt_6_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a = {1'b1
      , FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_6_lpi_1_dfm_8 , 31'b0};
  wire [5:0] nl_cvt_6_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s;
  assign nl_cvt_6_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s = {cvt_6_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_9_3_0_1[0]))};
  wire [41:0] nl_cvt_7_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a;
  assign nl_cvt_7_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a = {1'b1
      , FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_7_lpi_1_dfm_8 , 31'b0};
  wire [5:0] nl_cvt_7_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s;
  assign nl_cvt_7_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s = {cvt_7_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_9_3_0_1[0]))};
  wire [41:0] nl_cvt_8_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_a;
  assign nl_cvt_8_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_a = {1'b1
      , FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_8_lpi_1_dfm_8 , 31'b0};
  wire [5:0] nl_cvt_8_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s;
  assign nl_cvt_8_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s = {cvt_8_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_9_3_0_1[0]))};
  wire [41:0] nl_cvt_9_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_a;
  assign nl_cvt_9_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_a = {1'b1
      , FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_9_lpi_1_dfm_8 , 31'b0};
  wire [5:0] nl_cvt_9_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s;
  assign nl_cvt_9_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s = {cvt_9_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_9_3_0_1[0]))};
  wire [41:0] nl_cvt_10_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a;
  assign nl_cvt_10_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a = {1'b1
      , FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_10_lpi_1_dfm_8 , 31'b0};
  wire [5:0] nl_cvt_10_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s;
  assign nl_cvt_10_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s = {cvt_10_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_9_3_0_1[0]))};
  wire [41:0] nl_cvt_11_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a;
  assign nl_cvt_11_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a = {1'b1
      , FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_11_lpi_1_dfm_8 , 31'b0};
  wire [5:0] nl_cvt_11_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s;
  assign nl_cvt_11_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s = {cvt_11_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_9_3_0_1[0]))};
  wire [41:0] nl_cvt_12_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_a;
  assign nl_cvt_12_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_a = {1'b1
      , FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_12_lpi_1_dfm_8 , 31'b0};
  wire [5:0] nl_cvt_12_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s;
  assign nl_cvt_12_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s = {cvt_12_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_9_3_0_1[0]))};
  wire [41:0] nl_cvt_13_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a;
  assign nl_cvt_13_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a = {1'b1
      , FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_13_lpi_1_dfm_8 , 31'b0};
  wire [5:0] nl_cvt_13_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s;
  assign nl_cvt_13_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s = {cvt_13_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_9_3_0_1[0]))};
  wire [41:0] nl_cvt_14_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_a;
  assign nl_cvt_14_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_a = {1'b1
      , FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_14_lpi_1_dfm_8 , 31'b0};
  wire [5:0] nl_cvt_14_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s;
  assign nl_cvt_14_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s = {cvt_14_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_9_3_0_1[0]))};
  wire [41:0] nl_cvt_15_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_a;
  assign nl_cvt_15_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_a = {1'b1
      , FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_15_lpi_1_dfm_8 , 31'b0};
  wire [5:0] nl_cvt_15_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s;
  assign nl_cvt_15_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s = {cvt_15_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_9_3_0_1[0]))};
  wire [41:0] nl_cvt_16_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_4_rg_a;
  assign nl_cvt_16_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_4_rg_a = {1'b1
      , FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_lpi_1_dfm_9 , 31'b0};
  wire [5:0] nl_cvt_16_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_4_rg_s;
  assign nl_cvt_16_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_4_rg_s = {cvt_16_FpFloatToInt_16U_5U_10U_shift_acc_4_itm_2
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_9_3_0_1[0]))};
  wire [16:0] nl_cvt_1_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_rg_a;
  assign nl_cvt_1_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_rg_a = {cvt_1_FpIntToFloat_17U_5U_10U_else_i_abs_conc_3_16
      , FpIntToFloat_17U_5U_10U_else_i_abs_15_1_1_lpi_1_dfm_5 , FpIntToFloat_17U_5U_10U_else_i_abs_0_1_lpi_1_dfm_5};
  wire [16:0] nl_cvt_1_leading_sign_17_0_rg_mantissa;
  assign nl_cvt_1_leading_sign_17_0_rg_mantissa = {cvt_1_FpIntToFloat_17U_5U_10U_else_i_abs_conc_3_16
      , FpIntToFloat_17U_5U_10U_else_i_abs_15_1_1_lpi_1_dfm_5 , FpIntToFloat_17U_5U_10U_else_i_abs_0_1_lpi_1_dfm_5};
  wire [16:0] nl_cvt_2_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg_a;
  assign nl_cvt_2_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg_a = {cvt_2_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16
      , FpIntToFloat_17U_5U_10U_else_i_abs_15_1_2_lpi_1_dfm_6 , FpIntToFloat_17U_5U_10U_else_i_abs_0_2_lpi_1_dfm_6};
  wire [16:0] nl_cvt_2_leading_sign_17_0_1_rg_mantissa;
  assign nl_cvt_2_leading_sign_17_0_1_rg_mantissa = {cvt_2_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16
      , FpIntToFloat_17U_5U_10U_else_i_abs_15_1_2_lpi_1_dfm_6 , FpIntToFloat_17U_5U_10U_else_i_abs_0_2_lpi_1_dfm_6};
  wire [16:0] nl_cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg_a;
  assign nl_cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg_a = {cvt_3_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16
      , FpIntToFloat_17U_5U_10U_else_i_abs_15_1_3_lpi_1_dfm_6 , FpIntToFloat_17U_5U_10U_else_i_abs_0_3_lpi_1_dfm_6};
  wire [16:0] nl_cvt_3_leading_sign_17_0_1_rg_mantissa;
  assign nl_cvt_3_leading_sign_17_0_1_rg_mantissa = {cvt_3_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16
      , FpIntToFloat_17U_5U_10U_else_i_abs_15_1_3_lpi_1_dfm_6 , FpIntToFloat_17U_5U_10U_else_i_abs_0_3_lpi_1_dfm_6};
  wire [16:0] nl_cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a;
  assign nl_cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a = {cvt_4_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16
      , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_4_lpi_1_dfm_6_reg , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_4_lpi_1_dfm_6_1_reg
      , FpIntToFloat_17U_5U_10U_else_i_abs_0_4_lpi_1_dfm_7};
  wire [16:0] nl_cvt_4_leading_sign_17_0_2_rg_mantissa;
  assign nl_cvt_4_leading_sign_17_0_2_rg_mantissa = {cvt_4_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16
      , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_4_lpi_1_dfm_6_reg , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_4_lpi_1_dfm_6_1_reg
      , FpIntToFloat_17U_5U_10U_else_i_abs_0_4_lpi_1_dfm_7};
  wire [16:0] nl_cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg_a;
  assign nl_cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg_a = {cvt_5_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16
      , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_5_lpi_1_dfm_5_reg , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_5_lpi_1_dfm_5_1_reg
      , FpIntToFloat_17U_5U_10U_else_i_abs_0_5_lpi_1_dfm_6};
  wire [16:0] nl_cvt_5_leading_sign_17_0_1_rg_mantissa;
  assign nl_cvt_5_leading_sign_17_0_1_rg_mantissa = {cvt_5_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16
      , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_5_lpi_1_dfm_5_reg , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_5_lpi_1_dfm_5_1_reg
      , FpIntToFloat_17U_5U_10U_else_i_abs_0_5_lpi_1_dfm_6};
  wire [16:0] nl_cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a;
  assign nl_cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a = {cvt_6_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16
      , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_6_lpi_1_dfm_6_reg , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_6_lpi_1_dfm_6_1_reg
      , FpIntToFloat_17U_5U_10U_else_i_abs_0_6_lpi_1_dfm_7};
  wire [16:0] nl_cvt_6_leading_sign_17_0_2_rg_mantissa;
  assign nl_cvt_6_leading_sign_17_0_2_rg_mantissa = {cvt_6_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16
      , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_6_lpi_1_dfm_6_reg , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_6_lpi_1_dfm_6_1_reg
      , FpIntToFloat_17U_5U_10U_else_i_abs_0_6_lpi_1_dfm_7};
  wire [16:0] nl_cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a;
  assign nl_cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a = {cvt_7_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16
      , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_7_lpi_1_dfm_6_reg , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_7_lpi_1_dfm_6_1_reg
      , FpIntToFloat_17U_5U_10U_else_i_abs_0_7_lpi_1_dfm_7};
  wire [16:0] nl_cvt_7_leading_sign_17_0_2_rg_mantissa;
  assign nl_cvt_7_leading_sign_17_0_2_rg_mantissa = {cvt_7_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16
      , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_7_lpi_1_dfm_6_reg , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_7_lpi_1_dfm_6_1_reg
      , FpIntToFloat_17U_5U_10U_else_i_abs_0_7_lpi_1_dfm_7};
  wire [16:0] nl_cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg_a;
  assign nl_cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg_a = {cvt_8_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16
      , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_8_lpi_1_dfm_7_reg , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_8_lpi_1_dfm_7_1_reg
      , FpIntToFloat_17U_5U_10U_else_i_abs_0_8_lpi_1_dfm_8};
  wire [16:0] nl_cvt_8_leading_sign_17_0_3_rg_mantissa;
  assign nl_cvt_8_leading_sign_17_0_3_rg_mantissa = {cvt_8_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16
      , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_8_lpi_1_dfm_7_reg , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_8_lpi_1_dfm_7_1_reg
      , FpIntToFloat_17U_5U_10U_else_i_abs_0_8_lpi_1_dfm_8};
  wire [16:0] nl_cvt_9_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg_a;
  assign nl_cvt_9_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg_a = {cvt_9_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16
      , FpIntToFloat_17U_5U_10U_else_i_abs_15_1_9_lpi_1_dfm_6 , FpIntToFloat_17U_5U_10U_else_i_abs_0_9_lpi_1_dfm_6};
  wire [16:0] nl_cvt_9_leading_sign_17_0_1_rg_mantissa;
  assign nl_cvt_9_leading_sign_17_0_1_rg_mantissa = {cvt_9_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16
      , FpIntToFloat_17U_5U_10U_else_i_abs_15_1_9_lpi_1_dfm_6 , FpIntToFloat_17U_5U_10U_else_i_abs_0_9_lpi_1_dfm_6};
  wire [16:0] nl_cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a;
  assign nl_cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a = {cvt_10_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16
      , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_10_lpi_1_dfm_6_reg , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_10_lpi_1_dfm_6_1_reg
      , FpIntToFloat_17U_5U_10U_else_i_abs_0_10_lpi_1_dfm_7};
  wire [16:0] nl_cvt_10_leading_sign_17_0_2_rg_mantissa;
  assign nl_cvt_10_leading_sign_17_0_2_rg_mantissa = {cvt_10_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16
      , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_10_lpi_1_dfm_6_reg , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_10_lpi_1_dfm_6_1_reg
      , FpIntToFloat_17U_5U_10U_else_i_abs_0_10_lpi_1_dfm_7};
  wire [16:0] nl_cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a;
  assign nl_cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a = {cvt_11_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16
      , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_11_lpi_1_dfm_6_reg , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_11_lpi_1_dfm_6_1_reg
      , FpIntToFloat_17U_5U_10U_else_i_abs_0_11_lpi_1_dfm_7};
  wire [16:0] nl_cvt_11_leading_sign_17_0_2_rg_mantissa;
  assign nl_cvt_11_leading_sign_17_0_2_rg_mantissa = {cvt_11_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16
      , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_11_lpi_1_dfm_6_reg , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_11_lpi_1_dfm_6_1_reg
      , FpIntToFloat_17U_5U_10U_else_i_abs_0_11_lpi_1_dfm_7};
  wire [16:0] nl_cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg_a;
  assign nl_cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg_a = {cvt_12_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16
      , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_12_lpi_1_dfm_7_reg , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_12_lpi_1_dfm_7_1_reg
      , FpIntToFloat_17U_5U_10U_else_i_abs_0_12_lpi_1_dfm_8};
  wire [16:0] nl_cvt_12_leading_sign_17_0_3_rg_mantissa;
  assign nl_cvt_12_leading_sign_17_0_3_rg_mantissa = {cvt_12_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16
      , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_12_lpi_1_dfm_7_reg , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_12_lpi_1_dfm_7_1_reg
      , FpIntToFloat_17U_5U_10U_else_i_abs_0_12_lpi_1_dfm_8};
  wire [16:0] nl_cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a;
  assign nl_cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a = {cvt_13_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16
      , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_13_lpi_1_dfm_6_reg , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_13_lpi_1_dfm_6_1_reg
      , FpIntToFloat_17U_5U_10U_else_i_abs_0_13_lpi_1_dfm_7};
  wire [16:0] nl_cvt_13_leading_sign_17_0_2_rg_mantissa;
  assign nl_cvt_13_leading_sign_17_0_2_rg_mantissa = {cvt_13_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16
      , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_13_lpi_1_dfm_6_reg , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_13_lpi_1_dfm_6_1_reg
      , FpIntToFloat_17U_5U_10U_else_i_abs_0_13_lpi_1_dfm_7};
  wire [16:0] nl_cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg_a;
  assign nl_cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg_a = {cvt_14_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16
      , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_14_lpi_1_dfm_7_reg , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_14_lpi_1_dfm_7_1_reg
      , FpIntToFloat_17U_5U_10U_else_i_abs_0_14_lpi_1_dfm_8};
  wire [16:0] nl_cvt_14_leading_sign_17_0_3_rg_mantissa;
  assign nl_cvt_14_leading_sign_17_0_3_rg_mantissa = {cvt_14_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16
      , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_14_lpi_1_dfm_7_reg , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_14_lpi_1_dfm_7_1_reg
      , FpIntToFloat_17U_5U_10U_else_i_abs_0_14_lpi_1_dfm_8};
  wire [16:0] nl_cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg_a;
  assign nl_cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg_a = {cvt_15_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16
      , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_15_lpi_1_dfm_7_reg , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_15_lpi_1_dfm_7_1_reg
      , FpIntToFloat_17U_5U_10U_else_i_abs_0_15_lpi_1_dfm_8};
  wire [16:0] nl_cvt_15_leading_sign_17_0_3_rg_mantissa;
  assign nl_cvt_15_leading_sign_17_0_3_rg_mantissa = {cvt_15_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16
      , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_15_lpi_1_dfm_7_reg , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_15_lpi_1_dfm_7_1_reg
      , FpIntToFloat_17U_5U_10U_else_i_abs_0_15_lpi_1_dfm_8};
  wire [16:0] nl_cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_rg_a;
  assign nl_cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_rg_a = {cvt_16_FpIntToFloat_17U_5U_10U_else_i_abs_conc_7_16
      , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_lpi_1_dfm_8_reg , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_lpi_1_dfm_8_1_reg
      , FpIntToFloat_17U_5U_10U_else_i_abs_0_lpi_1_dfm_9};
  wire [16:0] nl_cvt_16_leading_sign_17_0_4_rg_mantissa;
  assign nl_cvt_16_leading_sign_17_0_4_rg_mantissa = {cvt_16_FpIntToFloat_17U_5U_10U_else_i_abs_conc_7_16
      , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_lpi_1_dfm_8_reg , reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_lpi_1_dfm_8_1_reg
      , FpIntToFloat_17U_5U_10U_else_i_abs_0_lpi_1_dfm_9};
  wire [23:0] nl_cvt_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_a;
  assign nl_cvt_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_a = {1'b1 , (chn_idata_data_sva_1_27_0_1[22:0])};
  wire [3:0] nl_cvt_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_s;
  assign nl_cvt_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_s = {FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_2_sva_2
      , (~ (chn_idata_data_sva_1_27_0_1[23]))};
  wire [5:0] nl_cvt_1_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg_s;
  assign nl_cvt_1_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg_s = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_1_sva_2
      + 5'b11111;
  wire [23:0] nl_cvt_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_a;
  assign nl_cvt_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_a = {1'b1 ,
      (chn_idata_data_sva_1_59_31_1[23:1])};
  wire [3:0] nl_cvt_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s;
  assign nl_cvt_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s = {FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_3_sva_2
      , (~ (chn_idata_data_sva_1_59_31_1[24]))};
  wire [5:0] nl_cvt_2_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg_s;
  assign nl_cvt_2_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg_s = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_2_sva_2
      + 5'b11111;
  wire [23:0] nl_cvt_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_a;
  assign nl_cvt_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_a = {1'b1 ,
      (chn_idata_data_sva_1_91_63_1[23:1])};
  wire [3:0] nl_cvt_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s;
  assign nl_cvt_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s = {FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_4_sva_2
      , (~ (chn_idata_data_sva_1_91_63_1[24]))};
  wire [5:0] nl_cvt_3_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg_s;
  assign nl_cvt_3_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg_s = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_3_sva_2
      + 5'b11111;
  wire [23:0] nl_cvt_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a;
  assign nl_cvt_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a = {1'b1 ,
      (chn_idata_data_sva_1_123_95_1[23:1])};
  wire [3:0] nl_cvt_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s;
  assign nl_cvt_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s = {FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_5_sva_2
      , (~ (chn_idata_data_sva_1_123_95_1[24]))};
  wire [5:0] nl_cvt_4_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s;
  assign nl_cvt_4_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_4_sva_2
      + 5'b11111;
  wire [23:0] nl_cvt_5_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_a;
  assign nl_cvt_5_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_a = {1'b1 ,
      (chn_idata_data_sva_1_155_127_1[23:1])};
  wire [3:0] nl_cvt_5_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s;
  assign nl_cvt_5_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s = {FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_6_sva_2
      , (~ (chn_idata_data_sva_1_155_127_1[24]))};
  wire [5:0] nl_cvt_5_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg_s;
  assign nl_cvt_5_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg_s = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_5_sva_2
      + 5'b11111;
  wire [23:0] nl_cvt_6_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a;
  assign nl_cvt_6_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a = {1'b1 ,
      (chn_idata_data_sva_1_187_159_1[23:1])};
  wire [3:0] nl_cvt_6_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s;
  assign nl_cvt_6_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s = {FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_7_sva_2
      , (~ (chn_idata_data_sva_1_187_159_1[24]))};
  wire [5:0] nl_cvt_6_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s;
  assign nl_cvt_6_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_6_sva_2
      + 5'b11111;
  wire [23:0] nl_cvt_7_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a;
  assign nl_cvt_7_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a = {1'b1 ,
      (chn_idata_data_sva_1_219_191_1[23:1])};
  wire [3:0] nl_cvt_7_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s;
  assign nl_cvt_7_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s = {FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_8_sva_2
      , (~ (chn_idata_data_sva_1_219_191_1[24]))};
  wire [5:0] nl_cvt_7_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s;
  assign nl_cvt_7_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_7_sva_2
      + 5'b11111;
  wire [23:0] nl_cvt_8_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_a;
  assign nl_cvt_8_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_a = {1'b1 ,
      (chn_idata_data_sva_1_251_223_1[23:1])};
  wire [3:0] nl_cvt_8_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s;
  assign nl_cvt_8_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s = {FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_9_sva_2
      , (~ (chn_idata_data_sva_1_251_223_1[24]))};
  wire [5:0] nl_cvt_8_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg_s;
  assign nl_cvt_8_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg_s = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_8_sva_2
      + 5'b11111;
  wire [23:0] nl_cvt_9_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_a;
  assign nl_cvt_9_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_a = {1'b1 ,
      (chn_idata_data_sva_1_283_255_1[23:1])};
  wire [3:0] nl_cvt_9_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s;
  assign nl_cvt_9_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s = {FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_10_sva_2
      , (~ (chn_idata_data_sva_1_283_255_1[24]))};
  wire [5:0] nl_cvt_9_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg_s;
  assign nl_cvt_9_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg_s = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_9_sva_2
      + 5'b11111;
  wire [23:0] nl_cvt_10_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a;
  assign nl_cvt_10_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a = {1'b1
      , (chn_idata_data_sva_1_315_287_1[23:1])};
  wire [3:0] nl_cvt_10_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s;
  assign nl_cvt_10_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s = {FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_11_sva_2
      , (~ (chn_idata_data_sva_1_315_287_1[24]))};
  wire [5:0] nl_cvt_10_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s;
  assign nl_cvt_10_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_10_sva_2
      + 5'b11111;
  wire [23:0] nl_cvt_11_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a;
  assign nl_cvt_11_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a = {1'b1
      , (chn_idata_data_sva_1_347_319_1[23:1])};
  wire [3:0] nl_cvt_11_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s;
  assign nl_cvt_11_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s = {FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_12_sva_2
      , (~ (chn_idata_data_sva_1_347_319_1[24]))};
  wire [5:0] nl_cvt_11_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s;
  assign nl_cvt_11_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_11_sva_2
      + 5'b11111;
  wire [23:0] nl_cvt_12_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_a;
  assign nl_cvt_12_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_a = {1'b1
      , (chn_idata_data_sva_1_379_351_1[23:1])};
  wire [3:0] nl_cvt_12_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s;
  assign nl_cvt_12_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s = {FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_13_sva_2
      , (~ (chn_idata_data_sva_1_379_351_1[24]))};
  wire [5:0] nl_cvt_12_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg_s;
  assign nl_cvt_12_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg_s = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_12_sva_2
      + 5'b11111;
  wire [23:0] nl_cvt_13_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a;
  assign nl_cvt_13_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a = {1'b1
      , (chn_idata_data_sva_1_411_383_1[23:1])};
  wire [3:0] nl_cvt_13_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s;
  assign nl_cvt_13_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s = {FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_14_sva_2
      , (~ (chn_idata_data_sva_1_411_383_1[24]))};
  wire [5:0] nl_cvt_13_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s;
  assign nl_cvt_13_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_13_sva_2
      + 5'b11111;
  wire [23:0] nl_cvt_14_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_a;
  assign nl_cvt_14_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_a = {1'b1
      , (chn_idata_data_sva_1_443_415_1[23:1])};
  wire [3:0] nl_cvt_14_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s;
  assign nl_cvt_14_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s = {FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_15_sva_2
      , (~ (chn_idata_data_sva_1_443_415_1[24]))};
  wire [5:0] nl_cvt_14_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg_s;
  assign nl_cvt_14_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg_s = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_14_sva_2
      + 5'b11111;
  wire [23:0] nl_cvt_15_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_a;
  assign nl_cvt_15_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_a = {1'b1
      , (chn_idata_data_sva_1_475_447_1[23:1])};
  wire [3:0] nl_cvt_15_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s;
  assign nl_cvt_15_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s = {FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_16_sva_2
      , (~ (chn_idata_data_sva_1_475_447_1[24]))};
  wire [5:0] nl_cvt_15_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg_s;
  assign nl_cvt_15_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg_s = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_15_sva_2
      + 5'b11111;
  wire [23:0] nl_cvt_16_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_4_rg_a;
  assign nl_cvt_16_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_4_rg_a = {1'b1
      , (chn_idata_data_sva_1_507_479_1[23:1])};
  wire [3:0] nl_cvt_16_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_4_rg_s;
  assign nl_cvt_16_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_4_rg_s = {FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_2
      , (~ (chn_idata_data_sva_1_507_479_1[24]))};
  wire [5:0] nl_cvt_16_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_4_rg_s;
  assign nl_cvt_16_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_4_rg_s = FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva_2
      + 5'b11111;
  wire [271:0] nl_NV_NVDLA_SDP_CORE_c_core_chn_out_rsci_inst_chn_out_rsci_d;
  assign nl_NV_NVDLA_SDP_CORE_c_core_chn_out_rsci_inst_chn_out_rsci_d = {chn_out_rsci_d_271
      , chn_out_rsci_d_270 , chn_out_rsci_d_269 , chn_out_rsci_d_268 , chn_out_rsci_d_267
      , chn_out_rsci_d_266 , chn_out_rsci_d_265 , chn_out_rsci_d_264 , chn_out_rsci_d_263
      , chn_out_rsci_d_262 , chn_out_rsci_d_261 , chn_out_rsci_d_260 , chn_out_rsci_d_259
      , chn_out_rsci_d_258 , chn_out_rsci_d_257 , chn_out_rsci_d_256 , chn_out_rsci_d_255
      , chn_out_rsci_d_254 , chn_out_rsci_d_253_250 , chn_out_rsci_d_249_241 , chn_out_rsci_d_240
      , chn_out_rsci_d_239 , chn_out_rsci_d_238 , chn_out_rsci_d_237_234 , chn_out_rsci_d_233_225
      , chn_out_rsci_d_224 , chn_out_rsci_d_223 , chn_out_rsci_d_222 , chn_out_rsci_d_221_218
      , chn_out_rsci_d_217_209 , chn_out_rsci_d_208 , chn_out_rsci_d_207 , chn_out_rsci_d_206
      , chn_out_rsci_d_205_202 , chn_out_rsci_d_201_193 , chn_out_rsci_d_192 , chn_out_rsci_d_191
      , chn_out_rsci_d_190 , chn_out_rsci_d_189_186 , chn_out_rsci_d_185_177 , chn_out_rsci_d_176
      , chn_out_rsci_d_175 , chn_out_rsci_d_174 , chn_out_rsci_d_173_170 , chn_out_rsci_d_169_161
      , chn_out_rsci_d_160 , chn_out_rsci_d_159 , chn_out_rsci_d_158 , chn_out_rsci_d_157_154
      , chn_out_rsci_d_153_145 , chn_out_rsci_d_144 , chn_out_rsci_d_143 , chn_out_rsci_d_142
      , chn_out_rsci_d_141_138 , chn_out_rsci_d_137_129 , chn_out_rsci_d_128 , chn_out_rsci_d_127
      , chn_out_rsci_d_126 , chn_out_rsci_d_125_122 , chn_out_rsci_d_121_113 , chn_out_rsci_d_112
      , chn_out_rsci_d_111 , chn_out_rsci_d_110 , chn_out_rsci_d_109_106 , chn_out_rsci_d_105_97
      , chn_out_rsci_d_96 , chn_out_rsci_d_95 , chn_out_rsci_d_94 , chn_out_rsci_d_93_90
      , chn_out_rsci_d_89_81 , chn_out_rsci_d_80 , chn_out_rsci_d_79 , chn_out_rsci_d_78
      , chn_out_rsci_d_77_74 , chn_out_rsci_d_73_65 , chn_out_rsci_d_64 , chn_out_rsci_d_63
      , chn_out_rsci_d_62 , chn_out_rsci_d_61_58 , chn_out_rsci_d_57_49 , chn_out_rsci_d_48
      , chn_out_rsci_d_47 , chn_out_rsci_d_46 , chn_out_rsci_d_45_42 , chn_out_rsci_d_41_33
      , chn_out_rsci_d_32 , chn_out_rsci_d_31 , chn_out_rsci_d_30 , chn_out_rsci_d_29_26
      , chn_out_rsci_d_25_17 , chn_out_rsci_d_16 , chn_out_rsci_d_15 , chn_out_rsci_d_14
      , chn_out_rsci_d_13_10 , chn_out_rsci_d_9_1 , chn_out_rsci_d_0};
  SDP_C_mgc_in_wire_v1 #(.rscid(32'sd2),
  .width(32'sd32)) cfg_offset_rsci (
      .d(cfg_offset_rsci_d),
      .z(cfg_offset_rsc_z)
    );
  SDP_C_mgc_in_wire_v1 #(.rscid(32'sd3),
  .width(32'sd16)) cfg_scale_rsci (
      .d(cfg_scale_rsci_d),
      .z(cfg_scale_rsc_z)
    );
  SDP_C_mgc_in_wire_v1 #(.rscid(32'sd4),
  .width(32'sd6)) cfg_truncate_rsci (
      .d(cfg_truncate_rsci_d),
      .z(cfg_truncate_rsc_z)
    );
  SDP_C_mgc_in_wire_v1 #(.rscid(32'sd5),
  .width(32'sd2)) cfg_proc_precision_rsci (
      .d(cfg_proc_precision_rsci_d),
      .z(cfg_proc_precision_rsc_z)
    );
  SDP_C_mgc_in_wire_v1 #(.rscid(32'sd6),
  .width(32'sd2)) cfg_out_precision_rsci (
      .d(cfg_out_precision_rsci_d),
      .z(cfg_out_precision_rsc_z)
    );
  SDP_C_mgc_in_wire_v1 #(.rscid(32'sd7),
  .width(32'sd1)) cfg_mode_eql_rsci (
      .d(cfg_mode_eql_rsci_d),
      .z(cfg_mode_eql_rsc_z)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd49),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd49)) cvt_4_IntShiftRightSat_49U_6U_17U_i_rshift_2_rg (
      .a(IntMulExt_33U_16U_49U_return_4_sva_1),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRightSat_49U_6U_17U_i_4_sva_mx0w1)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd49),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd49)) cvt_6_IntShiftRightSat_49U_6U_17U_i_rshift_2_rg (
      .a(IntMulExt_33U_16U_49U_return_6_sva_1),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRightSat_49U_6U_17U_i_6_sva_mx0w1)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd49),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd49)) cvt_8_IntShiftRightSat_49U_6U_17U_i_rshift_3_rg (
      .a(IntMulExt_33U_16U_49U_return_8_sva_1),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRightSat_49U_6U_17U_i_8_sva_mx0w1)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd49),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd49)) cvt_7_IntShiftRightSat_49U_6U_17U_i_rshift_2_rg (
      .a(IntMulExt_33U_16U_49U_return_7_sva_1),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRightSat_49U_6U_17U_i_7_sva_mx0w1)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd49),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd49)) cvt_10_IntShiftRightSat_49U_6U_17U_i_rshift_2_rg (
      .a(IntMulExt_33U_16U_49U_return_10_sva_1),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRightSat_49U_6U_17U_i_10_sva_mx0w1)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd49),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd49)) cvt_12_IntShiftRightSat_49U_6U_17U_i_rshift_3_rg (
      .a(IntMulExt_33U_16U_49U_return_12_sva_1),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRightSat_49U_6U_17U_i_12_sva_mx0w1)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd49),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd49)) cvt_11_IntShiftRightSat_49U_6U_17U_i_rshift_2_rg (
      .a(IntMulExt_33U_16U_49U_return_11_sva_1),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRightSat_49U_6U_17U_i_11_sva_mx0w1)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd49),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd49)) cvt_14_IntShiftRightSat_49U_6U_17U_i_rshift_3_rg (
      .a(IntMulExt_33U_16U_49U_return_14_sva_1),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRightSat_49U_6U_17U_i_14_sva_mx0w1)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd49),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd49)) cvt_16_IntShiftRightSat_49U_6U_17U_i_rshift_4_rg (
      .a(IntMulExt_33U_16U_49U_return_sva_1),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRightSat_49U_6U_17U_i_sva_mx0w1)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd49),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd49)) cvt_15_IntShiftRightSat_49U_6U_17U_i_rshift_3_rg (
      .a(IntMulExt_33U_16U_49U_return_15_sva_1),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRightSat_49U_6U_17U_i_15_sva_mx0w1)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd49),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd49)) cvt_13_IntShiftRightSat_49U_6U_17U_i_rshift_2_rg (
      .a(IntMulExt_33U_16U_49U_return_13_sva_1),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRightSat_49U_6U_17U_i_13_sva_mx0w1)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd49),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd49)) cvt_1_IntShiftRightSat_49U_6U_17U_i_rshift_rg (
      .a(IntMulExt_33U_16U_49U_return_1_sva_2),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRightSat_49U_6U_17U_i_1_sva_mx0w0)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd49),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd49)) cvt_2_IntShiftRightSat_49U_6U_17U_i_rshift_1_rg (
      .a(IntMulExt_33U_16U_49U_return_2_sva_2),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRightSat_49U_6U_17U_i_2_sva_mx0w0)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd49),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd49)) cvt_3_IntShiftRightSat_49U_6U_17U_i_rshift_1_rg (
      .a(IntMulExt_33U_16U_49U_return_3_sva_2),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRightSat_49U_6U_17U_i_3_sva_mx0w0)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd49),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd49)) cvt_5_IntShiftRightSat_49U_6U_17U_i_rshift_1_rg (
      .a(IntMulExt_33U_16U_49U_return_5_sva_2),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRightSat_49U_6U_17U_i_5_sva_mx0w0)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd49),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd49)) cvt_9_IntShiftRightSat_49U_6U_17U_i_rshift_1_rg (
      .a(IntMulExt_33U_16U_49U_return_9_sva_2),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRightSat_49U_6U_17U_i_9_sva_mx0w0)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) cvt_2_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg (
      .a(nl_cvt_2_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg_a[111:0]),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) cvt_4_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg (
      .a(nl_cvt_4_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a[111:0]),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) cvt_3_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg (
      .a(nl_cvt_3_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg_a[111:0]),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) cvt_6_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg (
      .a(nl_cvt_6_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a[111:0]),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) cvt_8_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg (
      .a(nl_cvt_8_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg_a[111:0]),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) cvt_7_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg (
      .a(nl_cvt_7_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a[111:0]),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) cvt_5_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg (
      .a(nl_cvt_5_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg_a[111:0]),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) cvt_10_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg (
      .a(nl_cvt_10_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a[111:0]),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) cvt_12_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg (
      .a(nl_cvt_12_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg_a[111:0]),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) cvt_11_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg (
      .a(nl_cvt_11_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a[111:0]),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) cvt_14_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg (
      .a(nl_cvt_14_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg_a[111:0]),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) cvt_16_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_4_rg (
      .a(nl_cvt_16_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_4_rg_a[111:0]),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) cvt_15_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg (
      .a(nl_cvt_15_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_3_rg_a[111:0]),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) cvt_13_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg (
      .a(nl_cvt_13_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_2_rg_a[111:0]),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) cvt_9_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg (
      .a(nl_cvt_9_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_1_rg_a[111:0]),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd112),
  .signd_a(32'sd1),
  .width_s(32'sd6),
  .width_z(32'sd112)) cvt_1_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_rg (
      .a(nl_cvt_1_IntShiftRight_49U_6U_17U_mbits_fixed_rshift_rg_a[111:0]),
      .s(cfg_truncate_1_sva_2),
      .z(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva)
    );
  SDP_C_mgc_shift_br_v4 #(.width_a(32'sd42),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd75)) cvt_1_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_rg (
      .a(nl_cvt_1_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_rg_a[41:0]),
      .s(nl_cvt_1_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_rg_s[5:0]),
      .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva)
    );
  SDP_C_mgc_shift_br_v4 #(.width_a(32'sd42),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd75)) cvt_2_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg
      (
      .a(nl_cvt_2_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_a[41:0]),
      .s(nl_cvt_2_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s[5:0]),
      .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva)
    );
  SDP_C_mgc_shift_br_v4 #(.width_a(32'sd42),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd75)) cvt_3_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg
      (
      .a(nl_cvt_3_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_a[41:0]),
      .s(nl_cvt_3_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s[5:0]),
      .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva)
    );
  SDP_C_mgc_shift_br_v4 #(.width_a(32'sd42),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd75)) cvt_4_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg
      (
      .a(nl_cvt_4_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a[41:0]),
      .s(nl_cvt_4_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s[5:0]),
      .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva)
    );
  SDP_C_mgc_shift_br_v4 #(.width_a(32'sd42),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd75)) cvt_5_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg
      (
      .a(nl_cvt_5_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_a[41:0]),
      .s(nl_cvt_5_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s[5:0]),
      .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva)
    );
  SDP_C_mgc_shift_br_v4 #(.width_a(32'sd42),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd75)) cvt_6_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg
      (
      .a(nl_cvt_6_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a[41:0]),
      .s(nl_cvt_6_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s[5:0]),
      .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva)
    );
  SDP_C_mgc_shift_br_v4 #(.width_a(32'sd42),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd75)) cvt_7_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg
      (
      .a(nl_cvt_7_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a[41:0]),
      .s(nl_cvt_7_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s[5:0]),
      .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva)
    );
  SDP_C_mgc_shift_br_v4 #(.width_a(32'sd42),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd75)) cvt_8_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg
      (
      .a(nl_cvt_8_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_a[41:0]),
      .s(nl_cvt_8_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s[5:0]),
      .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva)
    );
  SDP_C_mgc_shift_br_v4 #(.width_a(32'sd42),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd75)) cvt_9_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg
      (
      .a(nl_cvt_9_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_a[41:0]),
      .s(nl_cvt_9_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_1_rg_s[5:0]),
      .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva)
    );
  SDP_C_mgc_shift_br_v4 #(.width_a(32'sd42),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd75)) cvt_10_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg
      (
      .a(nl_cvt_10_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a[41:0]),
      .s(nl_cvt_10_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s[5:0]),
      .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva)
    );
  SDP_C_mgc_shift_br_v4 #(.width_a(32'sd42),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd75)) cvt_11_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg
      (
      .a(nl_cvt_11_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a[41:0]),
      .s(nl_cvt_11_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s[5:0]),
      .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva)
    );
  SDP_C_mgc_shift_br_v4 #(.width_a(32'sd42),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd75)) cvt_12_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg
      (
      .a(nl_cvt_12_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_a[41:0]),
      .s(nl_cvt_12_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s[5:0]),
      .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva)
    );
  SDP_C_mgc_shift_br_v4 #(.width_a(32'sd42),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd75)) cvt_13_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg
      (
      .a(nl_cvt_13_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_a[41:0]),
      .s(nl_cvt_13_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_2_rg_s[5:0]),
      .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva)
    );
  SDP_C_mgc_shift_br_v4 #(.width_a(32'sd42),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd75)) cvt_14_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg
      (
      .a(nl_cvt_14_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_a[41:0]),
      .s(nl_cvt_14_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s[5:0]),
      .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva)
    );
  SDP_C_mgc_shift_br_v4 #(.width_a(32'sd42),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd75)) cvt_15_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg
      (
      .a(nl_cvt_15_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_a[41:0]),
      .s(nl_cvt_15_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_3_rg_s[5:0]),
      .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva)
    );
  SDP_C_mgc_shift_br_v4 #(.width_a(32'sd42),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd75)) cvt_16_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_4_rg
      (
      .a(nl_cvt_16_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_4_rg_a[41:0]),
      .s(nl_cvt_16_IntSignedShiftRight_12U_6U_26U_mbits_fixed_rshift_4_rg_s[5:0]),
      .z(IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd17),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd17)) cvt_1_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_rg (
      .a(nl_cvt_1_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_rg_a[16:0]),
      .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_16),
      .z(FpIntToFloat_17U_5U_10U_else_int_mant_1_sva)
    );
  SDP_C_leading_sign_17_0 cvt_1_leading_sign_17_0_rg (
      .mantissa(nl_cvt_1_leading_sign_17_0_rg_mantissa[16:0]),
      .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_16)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd17),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd17)) cvt_2_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg (
      .a(nl_cvt_2_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg_a[16:0]),
      .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_17),
      .z(FpIntToFloat_17U_5U_10U_else_int_mant_2_sva)
    );
  SDP_C_leading_sign_17_0 cvt_2_leading_sign_17_0_1_rg (
      .mantissa(nl_cvt_2_leading_sign_17_0_1_rg_mantissa[16:0]),
      .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_17)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd17),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd17)) cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg (
      .a(nl_cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg_a[16:0]),
      .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_18),
      .z(cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp)
    );
  SDP_C_leading_sign_17_0 cvt_3_leading_sign_17_0_1_rg (
      .mantissa(nl_cvt_3_leading_sign_17_0_1_rg_mantissa[16:0]),
      .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_18)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd17),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd17)) cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg (
      .a(nl_cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a[16:0]),
      .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_19),
      .z(cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp)
    );
  SDP_C_leading_sign_17_0 cvt_4_leading_sign_17_0_2_rg (
      .mantissa(nl_cvt_4_leading_sign_17_0_2_rg_mantissa[16:0]),
      .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_19)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd17),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd17)) cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg (
      .a(nl_cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg_a[16:0]),
      .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_20),
      .z(cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp)
    );
  SDP_C_leading_sign_17_0 cvt_5_leading_sign_17_0_1_rg (
      .mantissa(nl_cvt_5_leading_sign_17_0_1_rg_mantissa[16:0]),
      .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_20)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd17),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd17)) cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg (
      .a(nl_cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a[16:0]),
      .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_21),
      .z(cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp)
    );
  SDP_C_leading_sign_17_0 cvt_6_leading_sign_17_0_2_rg (
      .mantissa(nl_cvt_6_leading_sign_17_0_2_rg_mantissa[16:0]),
      .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_21)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd17),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd17)) cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg (
      .a(nl_cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a[16:0]),
      .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_22),
      .z(cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp)
    );
  SDP_C_leading_sign_17_0 cvt_7_leading_sign_17_0_2_rg (
      .mantissa(nl_cvt_7_leading_sign_17_0_2_rg_mantissa[16:0]),
      .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_22)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd17),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd17)) cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg (
      .a(nl_cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg_a[16:0]),
      .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_23),
      .z(cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp)
    );
  SDP_C_leading_sign_17_0 cvt_8_leading_sign_17_0_3_rg (
      .mantissa(nl_cvt_8_leading_sign_17_0_3_rg_mantissa[16:0]),
      .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_23)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd17),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd17)) cvt_9_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg (
      .a(nl_cvt_9_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_rg_a[16:0]),
      .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_24),
      .z(FpIntToFloat_17U_5U_10U_else_int_mant_9_sva)
    );
  SDP_C_leading_sign_17_0 cvt_9_leading_sign_17_0_1_rg (
      .mantissa(nl_cvt_9_leading_sign_17_0_1_rg_mantissa[16:0]),
      .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_24)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd17),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd17)) cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg (
      .a(nl_cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a[16:0]),
      .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_25),
      .z(cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp)
    );
  SDP_C_leading_sign_17_0 cvt_10_leading_sign_17_0_2_rg (
      .mantissa(nl_cvt_10_leading_sign_17_0_2_rg_mantissa[16:0]),
      .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_25)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd17),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd17)) cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg (
      .a(nl_cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a[16:0]),
      .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_26),
      .z(cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp)
    );
  SDP_C_leading_sign_17_0 cvt_11_leading_sign_17_0_2_rg (
      .mantissa(nl_cvt_11_leading_sign_17_0_2_rg_mantissa[16:0]),
      .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_26)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd17),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd17)) cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg (
      .a(nl_cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg_a[16:0]),
      .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_27),
      .z(cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp)
    );
  SDP_C_leading_sign_17_0 cvt_12_leading_sign_17_0_3_rg (
      .mantissa(nl_cvt_12_leading_sign_17_0_3_rg_mantissa[16:0]),
      .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_27)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd17),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd17)) cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg (
      .a(nl_cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_rg_a[16:0]),
      .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_28),
      .z(cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp)
    );
  SDP_C_leading_sign_17_0 cvt_13_leading_sign_17_0_2_rg (
      .mantissa(nl_cvt_13_leading_sign_17_0_2_rg_mantissa[16:0]),
      .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_28)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd17),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd17)) cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg (
      .a(nl_cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg_a[16:0]),
      .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_29),
      .z(cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp)
    );
  SDP_C_leading_sign_17_0 cvt_14_leading_sign_17_0_3_rg (
      .mantissa(nl_cvt_14_leading_sign_17_0_3_rg_mantissa[16:0]),
      .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_29)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd17),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd17)) cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg (
      .a(nl_cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_rg_a[16:0]),
      .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_30),
      .z(cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp)
    );
  SDP_C_leading_sign_17_0 cvt_15_leading_sign_17_0_3_rg (
      .mantissa(nl_cvt_15_leading_sign_17_0_3_rg_mantissa[16:0]),
      .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_30)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd17),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd17)) cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_rg (
      .a(nl_cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_rg_a[16:0]),
      .s(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_31),
      .z(cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_tmp)
    );
  SDP_C_leading_sign_17_0 cvt_16_leading_sign_17_0_4_rg (
      .mantissa(nl_cvt_16_leading_sign_17_0_4_rg_mantissa[16:0]),
      .rtn(libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_31)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd24)) cvt_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg (
      .a(nl_cvt_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_a[23:0]),
      .s(nl_cvt_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_rg_s[3:0]),
      .z(cvt_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_itm)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_1_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg (
      .a(1'b1),
      .s(nl_cvt_1_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_rg_s[4:0]),
      .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_1_sva)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_1_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_rg (
      .a(1'b1),
      .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_1_sva_2),
      .z(FpMantDecShiftRight_23U_8U_10U_least_mask_1_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd24)) cvt_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg (
      .a(nl_cvt_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_a[23:0]),
      .s(nl_cvt_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s[3:0]),
      .z(cvt_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_itm)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_2_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg
      (
      .a(1'b1),
      .s(nl_cvt_2_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg_s[4:0]),
      .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_2_sva)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_2_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_1_rg
      (
      .a(1'b1),
      .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_2_sva_2),
      .z(FpMantDecShiftRight_23U_8U_10U_least_mask_2_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd24)) cvt_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg (
      .a(nl_cvt_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_a[23:0]),
      .s(nl_cvt_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s[3:0]),
      .z(cvt_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_itm)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_3_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg
      (
      .a(1'b1),
      .s(nl_cvt_3_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg_s[4:0]),
      .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_3_sva)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_3_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_1_rg
      (
      .a(1'b1),
      .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_3_sva_2),
      .z(FpMantDecShiftRight_23U_8U_10U_least_mask_3_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd24)) cvt_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg (
      .a(nl_cvt_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a[23:0]),
      .s(nl_cvt_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s[3:0]),
      .z(cvt_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_4_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg
      (
      .a(1'b1),
      .s(nl_cvt_4_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s[4:0]),
      .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_4_sva)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_4_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_2_rg
      (
      .a(1'b1),
      .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_4_sva_2),
      .z(FpMantDecShiftRight_23U_8U_10U_least_mask_4_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd24)) cvt_5_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg (
      .a(nl_cvt_5_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_a[23:0]),
      .s(nl_cvt_5_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s[3:0]),
      .z(cvt_5_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_itm)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_5_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg
      (
      .a(1'b1),
      .s(nl_cvt_5_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg_s[4:0]),
      .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_5_sva)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_5_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_1_rg
      (
      .a(1'b1),
      .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_5_sva_2),
      .z(FpMantDecShiftRight_23U_8U_10U_least_mask_5_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd24)) cvt_6_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg (
      .a(nl_cvt_6_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a[23:0]),
      .s(nl_cvt_6_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s[3:0]),
      .z(cvt_6_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_6_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg
      (
      .a(1'b1),
      .s(nl_cvt_6_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s[4:0]),
      .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_6_sva)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_6_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_2_rg
      (
      .a(1'b1),
      .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_6_sva_2),
      .z(FpMantDecShiftRight_23U_8U_10U_least_mask_6_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd24)) cvt_7_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg (
      .a(nl_cvt_7_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a[23:0]),
      .s(nl_cvt_7_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s[3:0]),
      .z(cvt_7_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_7_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg
      (
      .a(1'b1),
      .s(nl_cvt_7_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s[4:0]),
      .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_7_sva)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_7_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_2_rg
      (
      .a(1'b1),
      .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_7_sva_2),
      .z(FpMantDecShiftRight_23U_8U_10U_least_mask_7_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd24)) cvt_8_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg (
      .a(nl_cvt_8_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_a[23:0]),
      .s(nl_cvt_8_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s[3:0]),
      .z(cvt_8_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_itm)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_8_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg
      (
      .a(1'b1),
      .s(nl_cvt_8_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg_s[4:0]),
      .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_8_sva)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_8_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_3_rg
      (
      .a(1'b1),
      .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_8_sva_2),
      .z(FpMantDecShiftRight_23U_8U_10U_least_mask_8_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd24)) cvt_9_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg (
      .a(nl_cvt_9_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_a[23:0]),
      .s(nl_cvt_9_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_rg_s[3:0]),
      .z(cvt_9_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_itm)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_9_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg
      (
      .a(1'b1),
      .s(nl_cvt_9_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_1_rg_s[4:0]),
      .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_9_sva)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_9_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_1_rg
      (
      .a(1'b1),
      .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_9_sva_2),
      .z(FpMantDecShiftRight_23U_8U_10U_least_mask_9_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd24)) cvt_10_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg (
      .a(nl_cvt_10_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a[23:0]),
      .s(nl_cvt_10_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s[3:0]),
      .z(cvt_10_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_10_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg
      (
      .a(1'b1),
      .s(nl_cvt_10_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s[4:0]),
      .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_10_sva)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_10_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_2_rg
      (
      .a(1'b1),
      .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_10_sva_2),
      .z(FpMantDecShiftRight_23U_8U_10U_least_mask_10_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd24)) cvt_11_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg (
      .a(nl_cvt_11_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a[23:0]),
      .s(nl_cvt_11_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s[3:0]),
      .z(cvt_11_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_11_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg
      (
      .a(1'b1),
      .s(nl_cvt_11_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s[4:0]),
      .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_11_sva)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_11_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_2_rg
      (
      .a(1'b1),
      .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_11_sva_2),
      .z(FpMantDecShiftRight_23U_8U_10U_least_mask_11_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd24)) cvt_12_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg (
      .a(nl_cvt_12_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_a[23:0]),
      .s(nl_cvt_12_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s[3:0]),
      .z(cvt_12_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_itm)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_12_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg
      (
      .a(1'b1),
      .s(nl_cvt_12_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg_s[4:0]),
      .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_12_sva)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_12_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_3_rg
      (
      .a(1'b1),
      .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_12_sva_2),
      .z(FpMantDecShiftRight_23U_8U_10U_least_mask_12_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd24)) cvt_13_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg (
      .a(nl_cvt_13_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_a[23:0]),
      .s(nl_cvt_13_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_rg_s[3:0]),
      .z(cvt_13_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_13_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg
      (
      .a(1'b1),
      .s(nl_cvt_13_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_2_rg_s[4:0]),
      .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_13_sva)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_13_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_2_rg
      (
      .a(1'b1),
      .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_13_sva_2),
      .z(FpMantDecShiftRight_23U_8U_10U_least_mask_13_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd24)) cvt_14_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg (
      .a(nl_cvt_14_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_a[23:0]),
      .s(nl_cvt_14_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s[3:0]),
      .z(cvt_14_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_itm)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_14_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg
      (
      .a(1'b1),
      .s(nl_cvt_14_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg_s[4:0]),
      .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_14_sva)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_14_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_3_rg
      (
      .a(1'b1),
      .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_14_sva_2),
      .z(FpMantDecShiftRight_23U_8U_10U_least_mask_14_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd24)) cvt_15_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg (
      .a(nl_cvt_15_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_a[23:0]),
      .s(nl_cvt_15_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_rg_s[3:0]),
      .z(cvt_15_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_itm)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_15_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg
      (
      .a(1'b1),
      .s(nl_cvt_15_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_3_rg_s[4:0]),
      .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_15_sva)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_15_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_3_rg
      (
      .a(1'b1),
      .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_15_sva_2),
      .z(FpMantDecShiftRight_23U_8U_10U_least_mask_15_sva)
    );
  SDP_C_mgc_shift_r_v4 #(.width_a(32'sd24),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd24)) cvt_16_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_4_rg (
      .a(nl_cvt_16_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_4_rg_a[23:0]),
      .s(nl_cvt_16_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_4_rg_s[3:0]),
      .z(cvt_16_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_4_itm)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_16_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_4_rg
      (
      .a(1'b1),
      .s(nl_cvt_16_FpMantDecShiftRight_23U_8U_10U_guard_mask_lshift_4_rg_s[4:0]),
      .z(FpMantDecShiftRight_23U_8U_10U_guard_mask_sva)
    );
  SDP_C_mgc_shift_l_v4 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd24)) cvt_16_FpMantDecShiftRight_23U_8U_10U_least_mask_lshift_4_rg
      (
      .a(1'b1),
      .s(FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva_2),
      .z(FpMantDecShiftRight_23U_8U_10U_least_mask_sva)
    );
  NV_NVDLA_SDP_CORE_c_core_chn_in_rsci NV_NVDLA_SDP_CORE_c_core_chn_in_rsci_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_in_rsc_z(chn_in_rsc_z),
      .chn_in_rsc_vz(chn_in_rsc_vz),
      .chn_in_rsc_lz(chn_in_rsc_lz),
      .chn_in_rsci_oswt(chn_in_rsci_oswt),
      .core_wen(core_wen),
      .chn_in_rsci_iswt0(chn_in_rsci_iswt0),
      .chn_in_rsci_bawt(chn_in_rsci_bawt),
      .chn_in_rsci_wen_comp(chn_in_rsci_wen_comp),
      .chn_in_rsci_ld_core_psct(chn_in_rsci_ld_core_psct),
      .chn_in_rsci_d_mxwt(chn_in_rsci_d_mxwt),
      .core_wten(core_wten)
    );
  NV_NVDLA_SDP_CORE_c_core_chn_out_rsci NV_NVDLA_SDP_CORE_c_core_chn_out_rsci_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_out_rsc_z(chn_out_rsc_z),
      .chn_out_rsc_vz(chn_out_rsc_vz),
      .chn_out_rsc_lz(chn_out_rsc_lz),
      .chn_out_rsci_oswt(chn_out_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_out_rsci_iswt0(chn_out_rsci_iswt0),
      .chn_out_rsci_bawt(chn_out_rsci_bawt),
      .chn_out_rsci_wen_comp(chn_out_rsci_wen_comp),
      .chn_out_rsci_ld_core_psct(reg_chn_out_rsci_ld_core_psct_cse),
      .chn_out_rsci_d(nl_NV_NVDLA_SDP_CORE_c_core_chn_out_rsci_inst_chn_out_rsci_d[271:0])
    );
  NV_NVDLA_SDP_CORE_c_core_staller NV_NVDLA_SDP_CORE_c_core_staller_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .chn_in_rsci_wen_comp(chn_in_rsci_wen_comp),
      .core_wten(core_wten),
      .chn_out_rsci_wen_comp(chn_out_rsci_wen_comp)
    );
  NV_NVDLA_SDP_CORE_c_core_core_fsm NV_NVDLA_SDP_CORE_c_core_core_fsm_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign and_15 = and_dcpl_4 & main_stage_v_1 & cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_2
      & (~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_st_2
      | cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_2));
  assign shift_0_prb = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_2_sva_2)
      , (chn_idata_data_sva_1_27_0_1[23])}) + 5'b1)), and_15);
// assert(shift > 0) - ../include/nvdla_float.h: line 286
// PSL cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln286_assert_shift_gt_0 : assert { shift_0_prb } @rose(nvdla_core_clk);
  assign and_19 = and_dcpl_4 & main_stage_v_1 & cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2
      & (~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_st_2
      | cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2));
  assign shift_0_prb_1 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_3_sva_2)
      , (chn_idata_data_sva_1_59_31_1[24])}) + 5'b1)), and_19);
// assert(shift > 0) - ../include/nvdla_float.h: line 286
// PSL cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln286_assert_shift_gt_0_1 : assert { shift_0_prb_1 } @rose(nvdla_core_clk);
  assign and_23 = and_dcpl_4 & main_stage_v_1 & cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2
      & (~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_st_2
      | cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2));
  assign shift_0_prb_2 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_4_sva_2)
      , (chn_idata_data_sva_1_91_63_1[24])}) + 5'b1)), and_23);
// assert(shift > 0) - ../include/nvdla_float.h: line 286
// PSL cvt_3_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln286_assert_shift_gt_0_1 : assert { shift_0_prb_2 } @rose(nvdla_core_clk);
  assign and_27 = and_dcpl_4 & main_stage_v_1 & cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
      & (~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_st_2
      | cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2));
  assign shift_0_prb_3 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_5_sva_2)
      , (chn_idata_data_sva_1_123_95_1[24])}) + 5'b1)), and_27);
// assert(shift > 0) - ../include/nvdla_float.h: line 286
// PSL cvt_4_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln286_assert_shift_gt_0_2 : assert { shift_0_prb_3 } @rose(nvdla_core_clk);
  assign and_32 = and_dcpl_3 & main_stage_v_1 & cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2
      & (~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_st_2
      | cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2))
      & or_5189_cse;
  assign shift_0_prb_4 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_6_sva_2)
      , (chn_idata_data_sva_1_155_127_1[24])}) + 5'b1)), and_32);
// assert(shift > 0) - ../include/nvdla_float.h: line 286
// PSL cvt_5_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln286_assert_shift_gt_0_1 : assert { shift_0_prb_4 } @rose(nvdla_core_clk);
  assign and_37 = and_dcpl_3 & main_stage_v_1 & cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
      & (~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_st_2
      | cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2))
      & or_5189_cse;
  assign shift_0_prb_5 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_7_sva_2)
      , (chn_idata_data_sva_1_187_159_1[24])}) + 5'b1)), and_37);
// assert(shift > 0) - ../include/nvdla_float.h: line 286
// PSL cvt_6_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln286_assert_shift_gt_0_2 : assert { shift_0_prb_5 } @rose(nvdla_core_clk);
  assign and_41 = and_dcpl_4 & main_stage_v_1 & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_st_2)
      & cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
      & (~ cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2);
  assign shift_0_prb_6 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_8_sva_2)
      , (chn_idata_data_sva_1_219_191_1[24])}) + 5'b1)), and_41);
// assert(shift > 0) - ../include/nvdla_float.h: line 286
// PSL cvt_7_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln286_assert_shift_gt_0_2 : assert { shift_0_prb_6 } @rose(nvdla_core_clk);
  assign and_45 = and_dcpl_4 & main_stage_v_1 & cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2
      & (~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_st_2
      | cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2));
  assign shift_0_prb_7 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_9_sva_2)
      , (chn_idata_data_sva_1_251_223_1[24])}) + 5'b1)), and_45);
// assert(shift > 0) - ../include/nvdla_float.h: line 286
// PSL cvt_8_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln286_assert_shift_gt_0_3 : assert { shift_0_prb_7 } @rose(nvdla_core_clk);
  assign and_49 = and_dcpl_4 & main_stage_v_1 & cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2
      & (~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_st_2
      | cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2));
  assign shift_0_prb_8 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_10_sva_2)
      , (chn_idata_data_sva_1_283_255_1[24])}) + 5'b1)), and_49);
// assert(shift > 0) - ../include/nvdla_float.h: line 286
// PSL cvt_9_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln286_assert_shift_gt_0_1 : assert { shift_0_prb_8 } @rose(nvdla_core_clk);
  assign and_54 = and_dcpl_3 & main_stage_v_1 & cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
      & (~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_st_2
      | cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2))
      & or_5189_cse;
  assign shift_0_prb_9 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_11_sva_2)
      , (chn_idata_data_sva_1_315_287_1[24])}) + 5'b1)), and_54);
// assert(shift > 0) - ../include/nvdla_float.h: line 286
// PSL cvt_10_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln286_assert_shift_gt_0_2 : assert { shift_0_prb_9 } @rose(nvdla_core_clk);
  assign and_58 = and_dcpl_4 & main_stage_v_1 & cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
      & (~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_st_2
      | cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2));
  assign shift_0_prb_10 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_12_sva_2)
      , (chn_idata_data_sva_1_347_319_1[24])}) + 5'b1)), and_58);
// assert(shift > 0) - ../include/nvdla_float.h: line 286
// PSL cvt_11_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln286_assert_shift_gt_0_2 : assert { shift_0_prb_10 } @rose(nvdla_core_clk);
  assign and_62 = and_dcpl_4 & main_stage_v_1 & cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2
      & (~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_st_2
      | cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2));
  assign shift_0_prb_11 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_13_sva_2)
      , (chn_idata_data_sva_1_379_351_1[24])}) + 5'b1)), and_62);
// assert(shift > 0) - ../include/nvdla_float.h: line 286
// PSL cvt_12_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln286_assert_shift_gt_0_3 : assert { shift_0_prb_11 } @rose(nvdla_core_clk);
  assign and_67 = and_dcpl_3 & main_stage_v_1 & cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
      & (~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_st_2
      | cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2))
      & or_5189_cse;
  assign shift_0_prb_12 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_14_sva_2)
      , (chn_idata_data_sva_1_411_383_1[24])}) + 5'b1)), and_67);
// assert(shift > 0) - ../include/nvdla_float.h: line 286
// PSL cvt_13_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln286_assert_shift_gt_0_2 : assert { shift_0_prb_12 } @rose(nvdla_core_clk);
  assign and_71 = and_dcpl_4 & main_stage_v_1 & cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2
      & (~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_st_2
      | cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2));
  assign shift_0_prb_13 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_15_sva_2)
      , (chn_idata_data_sva_1_443_415_1[24])}) + 5'b1)), and_71);
// assert(shift > 0) - ../include/nvdla_float.h: line 286
// PSL cvt_14_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln286_assert_shift_gt_0_3 : assert { shift_0_prb_13 } @rose(nvdla_core_clk);
  assign and_75 = and_dcpl_4 & main_stage_v_1 & cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2
      & (~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_st_2
      | cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2));
  assign shift_0_prb_14 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_16_sva_2)
      , (chn_idata_data_sva_1_475_447_1[24])}) + 5'b1)), and_75);
// assert(shift > 0) - ../include/nvdla_float.h: line 286
// PSL cvt_15_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln286_assert_shift_gt_0_3 : assert { shift_0_prb_14 } @rose(nvdla_core_clk);
  assign and_79 = and_dcpl_4 & main_stage_v_1 & cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_4_svs_st_2
      & (~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_2
      | cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_st_2));
  assign shift_0_prb_15 = MUX1HOT_s_1_1_2(readslicef_5_1_4((({1'b1 , (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_2)
      , (chn_idata_data_sva_1_507_479_1[24])}) + 5'b1)), and_79);
// assert(shift > 0) - ../include/nvdla_float.h: line 286
// PSL cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln286_assert_shift_gt_0_4 : assert { shift_0_prb_15 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iMantWidth >= oMantWidth) - ../include/nvdla_float.h: line 669
// PSL cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln669_assert_iMantWidth_ge_oMantWidth : assert { iMantWidth_oMantWidth_prb } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iExpoWidth >= oExpoWidth) - ../include/nvdla_float.h: line 670
// PSL cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth : assert { iExpoWidth_oExpoWidth_prb } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_1 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iMantWidth >= oMantWidth) - ../include/nvdla_float.h: line 669
// PSL cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln669_assert_iMantWidth_ge_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_1 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_1 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iExpoWidth >= oExpoWidth) - ../include/nvdla_float.h: line 670
// PSL cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_1 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_2 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iMantWidth >= oMantWidth) - ../include/nvdla_float.h: line 669
// PSL cvt_3_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln669_assert_iMantWidth_ge_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_2 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_2 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iExpoWidth >= oExpoWidth) - ../include/nvdla_float.h: line 670
// PSL cvt_3_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_2 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_3 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iMantWidth >= oMantWidth) - ../include/nvdla_float.h: line 669
// PSL cvt_4_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln669_assert_iMantWidth_ge_oMantWidth_2 : assert { iMantWidth_oMantWidth_prb_3 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_3 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iExpoWidth >= oExpoWidth) - ../include/nvdla_float.h: line 670
// PSL cvt_4_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_2 : assert { iExpoWidth_oExpoWidth_prb_3 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_4 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iMantWidth >= oMantWidth) - ../include/nvdla_float.h: line 669
// PSL cvt_5_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln669_assert_iMantWidth_ge_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_4 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_4 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iExpoWidth >= oExpoWidth) - ../include/nvdla_float.h: line 670
// PSL cvt_5_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_4 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_5 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iMantWidth >= oMantWidth) - ../include/nvdla_float.h: line 669
// PSL cvt_6_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln669_assert_iMantWidth_ge_oMantWidth_2 : assert { iMantWidth_oMantWidth_prb_5 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_5 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iExpoWidth >= oExpoWidth) - ../include/nvdla_float.h: line 670
// PSL cvt_6_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_2 : assert { iExpoWidth_oExpoWidth_prb_5 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_6 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iMantWidth >= oMantWidth) - ../include/nvdla_float.h: line 669
// PSL cvt_7_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln669_assert_iMantWidth_ge_oMantWidth_2 : assert { iMantWidth_oMantWidth_prb_6 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_6 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iExpoWidth >= oExpoWidth) - ../include/nvdla_float.h: line 670
// PSL cvt_7_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_2 : assert { iExpoWidth_oExpoWidth_prb_6 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_7 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iMantWidth >= oMantWidth) - ../include/nvdla_float.h: line 669
// PSL cvt_8_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln669_assert_iMantWidth_ge_oMantWidth_3 : assert { iMantWidth_oMantWidth_prb_7 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_7 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iExpoWidth >= oExpoWidth) - ../include/nvdla_float.h: line 670
// PSL cvt_8_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_3 : assert { iExpoWidth_oExpoWidth_prb_7 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_8 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iMantWidth >= oMantWidth) - ../include/nvdla_float.h: line 669
// PSL cvt_9_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln669_assert_iMantWidth_ge_oMantWidth_1 : assert { iMantWidth_oMantWidth_prb_8 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_8 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iExpoWidth >= oExpoWidth) - ../include/nvdla_float.h: line 670
// PSL cvt_9_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_1 : assert { iExpoWidth_oExpoWidth_prb_8 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_9 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iMantWidth >= oMantWidth) - ../include/nvdla_float.h: line 669
// PSL cvt_10_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln669_assert_iMantWidth_ge_oMantWidth_2 : assert { iMantWidth_oMantWidth_prb_9 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_9 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iExpoWidth >= oExpoWidth) - ../include/nvdla_float.h: line 670
// PSL cvt_10_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_2 : assert { iExpoWidth_oExpoWidth_prb_9 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_10 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iMantWidth >= oMantWidth) - ../include/nvdla_float.h: line 669
// PSL cvt_11_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln669_assert_iMantWidth_ge_oMantWidth_2 : assert { iMantWidth_oMantWidth_prb_10 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_10 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iExpoWidth >= oExpoWidth) - ../include/nvdla_float.h: line 670
// PSL cvt_11_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_2 : assert { iExpoWidth_oExpoWidth_prb_10 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_11 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iMantWidth >= oMantWidth) - ../include/nvdla_float.h: line 669
// PSL cvt_12_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln669_assert_iMantWidth_ge_oMantWidth_3 : assert { iMantWidth_oMantWidth_prb_11 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_11 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iExpoWidth >= oExpoWidth) - ../include/nvdla_float.h: line 670
// PSL cvt_12_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_3 : assert { iExpoWidth_oExpoWidth_prb_11 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_12 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iMantWidth >= oMantWidth) - ../include/nvdla_float.h: line 669
// PSL cvt_13_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln669_assert_iMantWidth_ge_oMantWidth_2 : assert { iMantWidth_oMantWidth_prb_12 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_12 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iExpoWidth >= oExpoWidth) - ../include/nvdla_float.h: line 670
// PSL cvt_13_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_2 : assert { iExpoWidth_oExpoWidth_prb_12 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_13 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iMantWidth >= oMantWidth) - ../include/nvdla_float.h: line 669
// PSL cvt_14_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln669_assert_iMantWidth_ge_oMantWidth_3 : assert { iMantWidth_oMantWidth_prb_13 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_13 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iExpoWidth >= oExpoWidth) - ../include/nvdla_float.h: line 670
// PSL cvt_14_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_3 : assert { iExpoWidth_oExpoWidth_prb_13 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_14 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iMantWidth >= oMantWidth) - ../include/nvdla_float.h: line 669
// PSL cvt_15_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln669_assert_iMantWidth_ge_oMantWidth_3 : assert { iMantWidth_oMantWidth_prb_14 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_14 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iExpoWidth >= oExpoWidth) - ../include/nvdla_float.h: line 670
// PSL cvt_15_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_3 : assert { iExpoWidth_oExpoWidth_prb_14 } @rose(nvdla_core_clk);
  assign iMantWidth_oMantWidth_prb_15 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iMantWidth >= oMantWidth) - ../include/nvdla_float.h: line 669
// PSL cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln669_assert_iMantWidth_ge_oMantWidth_4 : assert { iMantWidth_oMantWidth_prb_15 } @rose(nvdla_core_clk);
  assign iExpoWidth_oExpoWidth_prb_15 = cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1;
// assert(iExpoWidth >= oExpoWidth) - ../include/nvdla_float.h: line 670
// PSL cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4 : assert { iExpoWidth_oExpoWidth_prb_15 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth > mWidth) - ../include/nvdla_int.h: line 281
// PSL cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln281_assert_oWidth_gt_mWidth : assert { oWidth_mWidth_prb } @rose(nvdla_core_clk);
  assign oWidth_aWidth_bWidth_prb = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth >= aWidth+bWidth) - ../include/nvdla_int.h: line 346
// PSL cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth : assert { oWidth_aWidth_bWidth_prb } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth : assert { oWidth_iWidth_prb } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_1 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1 : assert { oWidth_iWidth_prb_1 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_1 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth > mWidth) - ../include/nvdla_int.h: line 281
// PSL cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln281_assert_oWidth_gt_mWidth_1 : assert { oWidth_mWidth_prb_1 } @rose(nvdla_core_clk);
  assign oWidth_aWidth_bWidth_prb_1 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth >= aWidth+bWidth) - ../include/nvdla_int.h: line 346
// PSL cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1 : assert { oWidth_aWidth_bWidth_prb_1 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_2 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_2 : assert { oWidth_iWidth_prb_2 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_3 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_3 : assert { oWidth_iWidth_prb_3 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_2 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth > mWidth) - ../include/nvdla_int.h: line 281
// PSL cvt_3_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln281_assert_oWidth_gt_mWidth_1 : assert { oWidth_mWidth_prb_2 } @rose(nvdla_core_clk);
  assign oWidth_aWidth_bWidth_prb_2 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth >= aWidth+bWidth) - ../include/nvdla_int.h: line 346
// PSL cvt_3_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1 : assert { oWidth_aWidth_bWidth_prb_2 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_4 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_3_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_2 : assert { oWidth_iWidth_prb_4 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_5 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_3_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_3 : assert { oWidth_iWidth_prb_5 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_3 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth > mWidth) - ../include/nvdla_int.h: line 281
// PSL cvt_4_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln281_assert_oWidth_gt_mWidth_2 : assert { oWidth_mWidth_prb_3 } @rose(nvdla_core_clk);
  assign oWidth_aWidth_bWidth_prb_3 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth >= aWidth+bWidth) - ../include/nvdla_int.h: line 346
// PSL cvt_4_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_2 : assert { oWidth_aWidth_bWidth_prb_3 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_6 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_4_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_4 : assert { oWidth_iWidth_prb_6 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_7 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_4_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_5 : assert { oWidth_iWidth_prb_7 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_4 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth > mWidth) - ../include/nvdla_int.h: line 281
// PSL cvt_5_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln281_assert_oWidth_gt_mWidth_1 : assert { oWidth_mWidth_prb_4 } @rose(nvdla_core_clk);
  assign oWidth_aWidth_bWidth_prb_4 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth >= aWidth+bWidth) - ../include/nvdla_int.h: line 346
// PSL cvt_5_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1 : assert { oWidth_aWidth_bWidth_prb_4 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_8 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_5_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_2 : assert { oWidth_iWidth_prb_8 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_9 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_5_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_3 : assert { oWidth_iWidth_prb_9 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_5 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth > mWidth) - ../include/nvdla_int.h: line 281
// PSL cvt_6_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln281_assert_oWidth_gt_mWidth_2 : assert { oWidth_mWidth_prb_5 } @rose(nvdla_core_clk);
  assign oWidth_aWidth_bWidth_prb_5 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth >= aWidth+bWidth) - ../include/nvdla_int.h: line 346
// PSL cvt_6_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_2 : assert { oWidth_aWidth_bWidth_prb_5 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_10 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_6_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_4 : assert { oWidth_iWidth_prb_10 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_11 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_6_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_5 : assert { oWidth_iWidth_prb_11 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_6 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth > mWidth) - ../include/nvdla_int.h: line 281
// PSL cvt_7_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln281_assert_oWidth_gt_mWidth_2 : assert { oWidth_mWidth_prb_6 } @rose(nvdla_core_clk);
  assign oWidth_aWidth_bWidth_prb_6 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth >= aWidth+bWidth) - ../include/nvdla_int.h: line 346
// PSL cvt_7_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_2 : assert { oWidth_aWidth_bWidth_prb_6 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_12 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_7_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_4 : assert { oWidth_iWidth_prb_12 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_13 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_7_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_5 : assert { oWidth_iWidth_prb_13 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_7 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth > mWidth) - ../include/nvdla_int.h: line 281
// PSL cvt_8_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln281_assert_oWidth_gt_mWidth_3 : assert { oWidth_mWidth_prb_7 } @rose(nvdla_core_clk);
  assign oWidth_aWidth_bWidth_prb_7 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth >= aWidth+bWidth) - ../include/nvdla_int.h: line 346
// PSL cvt_8_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_3 : assert { oWidth_aWidth_bWidth_prb_7 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_14 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_8_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_6 : assert { oWidth_iWidth_prb_14 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_15 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_8_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_7 : assert { oWidth_iWidth_prb_15 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_8 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth > mWidth) - ../include/nvdla_int.h: line 281
// PSL cvt_9_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln281_assert_oWidth_gt_mWidth_1 : assert { oWidth_mWidth_prb_8 } @rose(nvdla_core_clk);
  assign oWidth_aWidth_bWidth_prb_8 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth >= aWidth+bWidth) - ../include/nvdla_int.h: line 346
// PSL cvt_9_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1 : assert { oWidth_aWidth_bWidth_prb_8 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_16 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_9_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_2 : assert { oWidth_iWidth_prb_16 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_17 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_9_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_3 : assert { oWidth_iWidth_prb_17 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_9 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth > mWidth) - ../include/nvdla_int.h: line 281
// PSL cvt_10_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln281_assert_oWidth_gt_mWidth_2 : assert { oWidth_mWidth_prb_9 } @rose(nvdla_core_clk);
  assign oWidth_aWidth_bWidth_prb_9 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth >= aWidth+bWidth) - ../include/nvdla_int.h: line 346
// PSL cvt_10_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_2 : assert { oWidth_aWidth_bWidth_prb_9 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_18 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_10_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_4 : assert { oWidth_iWidth_prb_18 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_19 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_10_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_5 : assert { oWidth_iWidth_prb_19 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_10 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth > mWidth) - ../include/nvdla_int.h: line 281
// PSL cvt_11_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln281_assert_oWidth_gt_mWidth_2 : assert { oWidth_mWidth_prb_10 } @rose(nvdla_core_clk);
  assign oWidth_aWidth_bWidth_prb_10 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth >= aWidth+bWidth) - ../include/nvdla_int.h: line 346
// PSL cvt_11_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_2 : assert { oWidth_aWidth_bWidth_prb_10 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_20 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_11_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_4 : assert { oWidth_iWidth_prb_20 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_21 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_11_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_5 : assert { oWidth_iWidth_prb_21 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_11 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth > mWidth) - ../include/nvdla_int.h: line 281
// PSL cvt_12_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln281_assert_oWidth_gt_mWidth_3 : assert { oWidth_mWidth_prb_11 } @rose(nvdla_core_clk);
  assign oWidth_aWidth_bWidth_prb_11 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth >= aWidth+bWidth) - ../include/nvdla_int.h: line 346
// PSL cvt_12_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_3 : assert { oWidth_aWidth_bWidth_prb_11 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_22 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_12_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_6 : assert { oWidth_iWidth_prb_22 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_23 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_12_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_7 : assert { oWidth_iWidth_prb_23 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_12 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth > mWidth) - ../include/nvdla_int.h: line 281
// PSL cvt_13_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln281_assert_oWidth_gt_mWidth_2 : assert { oWidth_mWidth_prb_12 } @rose(nvdla_core_clk);
  assign oWidth_aWidth_bWidth_prb_12 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth >= aWidth+bWidth) - ../include/nvdla_int.h: line 346
// PSL cvt_13_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_2 : assert { oWidth_aWidth_bWidth_prb_12 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_24 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_13_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_4 : assert { oWidth_iWidth_prb_24 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_25 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_13_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_5 : assert { oWidth_iWidth_prb_25 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_13 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth > mWidth) - ../include/nvdla_int.h: line 281
// PSL cvt_14_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln281_assert_oWidth_gt_mWidth_3 : assert { oWidth_mWidth_prb_13 } @rose(nvdla_core_clk);
  assign oWidth_aWidth_bWidth_prb_13 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth >= aWidth+bWidth) - ../include/nvdla_int.h: line 346
// PSL cvt_14_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_3 : assert { oWidth_aWidth_bWidth_prb_13 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_26 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_14_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_6 : assert { oWidth_iWidth_prb_26 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_27 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_14_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_7 : assert { oWidth_iWidth_prb_27 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_14 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth > mWidth) - ../include/nvdla_int.h: line 281
// PSL cvt_15_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln281_assert_oWidth_gt_mWidth_3 : assert { oWidth_mWidth_prb_14 } @rose(nvdla_core_clk);
  assign oWidth_aWidth_bWidth_prb_14 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth >= aWidth+bWidth) - ../include/nvdla_int.h: line 346
// PSL cvt_15_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_3 : assert { oWidth_aWidth_bWidth_prb_14 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_28 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_15_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_6 : assert { oWidth_iWidth_prb_28 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_29 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_15_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_7 : assert { oWidth_iWidth_prb_29 } @rose(nvdla_core_clk);
  assign oWidth_mWidth_prb_15 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth > mWidth) - ../include/nvdla_int.h: line 281
// PSL cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln281_assert_oWidth_gt_mWidth_4 : assert { oWidth_mWidth_prb_15 } @rose(nvdla_core_clk);
  assign oWidth_aWidth_bWidth_prb_15 = cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1;
// assert(oWidth >= aWidth+bWidth) - ../include/nvdla_int.h: line 346
// PSL cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_4 : assert { oWidth_aWidth_bWidth_prb_15 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_30 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_8 : assert { oWidth_iWidth_prb_30 } @rose(nvdla_core_clk);
  assign oWidth_iWidth_prb_31 = cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1_sig_mx0w1;
// assert(oWidth <= iWidth) - ../include/nvdla_int.h: line 402
// PSL cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_9 : assert { oWidth_iWidth_prb_31 } @rose(nvdla_core_clk);
  assign cvt_or_cse = cvt_asn_319 | (cvt_else_equal_tmp & (~ cfg_mode_eql_1_sva_6)
      & cvt_unequal_tmp_21);
  assign chn_out_and_cse = core_wen & (~ or_dcpl_4);
  assign or_5189_cse = (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt;
  assign and_3024_cse = ((~ cvt_unequal_tmp_21) | cfg_mode_eql_1_sva_6 | (cfg_out_precision_1_sva_6!=2'b11))
      & or_5189_cse & and_dcpl_1742;
  assign cvt_or_2_cse = cvt_asn_319 | (cvt_else_equal_tmp_3_mx0 & (~ cfg_mode_eql_1_sva_6)
      & cvt_unequal_tmp_21);
  assign cvt_or_6_cse = cvt_asn_319 | (cvt_else_equal_tmp_9_mx1 & (~ cfg_mode_eql_1_sva_6)
      & cvt_unequal_tmp_21);
  assign cvt_or_10_cse = cvt_asn_319 | (cvt_else_equal_tmp_15_mx0 & (~ cfg_mode_eql_1_sva_6)
      & cvt_unequal_tmp_21);
  assign cvt_or_12_cse = cvt_asn_319 | (cvt_else_equal_tmp_18_mx0 & (~ cfg_mode_eql_1_sva_6)
      & cvt_unequal_tmp_21);
  assign cvt_or_14_cse = cvt_asn_319 | (cvt_else_equal_tmp_21_mx1 & cvt_and_147_m1c);
  assign cvt_or_18_cse = cvt_asn_319 | (cvt_else_equal_tmp_27_mx0 & (~ cfg_mode_eql_1_sva_6)
      & cvt_unequal_tmp_21);
  assign cvt_or_20_cse = cvt_asn_319 | (cvt_else_equal_tmp_30_mx0 & (~ cfg_mode_eql_1_sva_6)
      & cvt_unequal_tmp_21);
  assign cvt_or_22_cse = cvt_asn_319 | (cvt_else_equal_tmp_33_mx1 & (~ cfg_mode_eql_1_sva_6)
      & cvt_unequal_tmp_21);
  assign cvt_or_24_cse = cvt_asn_319 | (cvt_else_equal_tmp_36_mx0 & (~ cfg_mode_eql_1_sva_6)
      & cvt_unequal_tmp_21);
  assign cvt_or_26_cse = cvt_asn_319 | (cvt_else_equal_tmp_39_mx1 & (~ cfg_mode_eql_1_sva_6)
      & cvt_unequal_tmp_21);
  assign mux_2354_nl = MUX_s_1_2_2(mux_tmp_2347, (~ or_tmp_4095), cfg_proc_precision_1_sva_st_90[1]);
  assign mux_2355_nl = MUX_s_1_2_2((mux_2354_nl), mux_tmp_2347, cfg_proc_precision_1_sva_st_90[0]);
  assign and_3063_cse = ((~ (mux_2355_nl)) | (~ cvt_unequal_tmp_21) | cfg_mode_eql_1_sva_6)
      & or_5189_cse & and_dcpl_1742;
  assign cvt_or_28_cse = cvt_asn_319 | (cvt_else_equal_tmp_42_mx0 & (~ cfg_mode_eql_1_sva_6)
      & cvt_unequal_tmp_21);
  assign or_5254_cse = (cfg_proc_precision_1_sva_st_108!=2'b10);
  assign cvt_or_30_cse = cvt_asn_319 | (cvt_else_equal_tmp_45_mx1 & cvt_unequal_tmp_21
      & (~ cfg_mode_eql_1_sva_6));
  assign chn_out_and_32_cse = core_wen & ((main_stage_v_3 & cvt_unequal_tmp_21 &
      or_5189_cse) | and_dcpl_98);
  assign chn_out_and_77_cse = core_wen & ((cfg_mode_eql_1_sva_6 & main_stage_v_3
      & or_5189_cse) | and_dcpl_102);
  assign nor_8_cse = ~((cfg_proc_precision_1_sva_st_64!=2'b10));
  assign and_2239_cse = cfg_mode_eql_1_sva_4 & main_stage_v_1;
  assign mux_12_nl = MUX_s_1_2_2(main_stage_v_1, chn_in_rsci_bawt, or_5189_cse);
  assign chn_idata_data_and_1_cse = core_wen & (~ and_dcpl_93) & (mux_12_nl);
  assign or_183_cse_1 = (reg_cfg_proc_precision_1_sva_st_40_cse!=2'b10);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse = core_wen & (~ and_dcpl_93) &
      (~ mux_tmp_6);
  assign IntMulExt_33U_16U_49U_and_11_cse = core_wen & (~ and_dcpl_93) & mux_133_cse;
  assign IntMulExt_33U_16U_49U_and_1_cse = core_wen & (and_550_cse | IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1);
  assign cfg_proc_precision_and_11_cse = core_wen & (~ and_dcpl_93) & mux_tmp_114;
  assign chn_idata_data_and_16_cse = core_wen & (~ and_dcpl_93) & mux_tmp_161;
  assign and_637_rgt = or_5189_cse & (~ IsNaN_8U_23U_land_1_lpi_1_dfm_3);
  assign nand_219_cse = ~((cfg_proc_precision_1_sva_st_65[1]) & (cfg_out_precision_1_sva_st_149[0]));
  assign nor_2047_cse = ~((cfg_out_precision_1_sva_st_154!=2'b01) | (~ main_stage_v_1)
      | (cfg_proc_precision_1_sva_st_64!=2'b10));
  assign and_639_rgt = or_5189_cse & (~ IsNaN_8U_23U_land_2_lpi_1_dfm_3);
  assign nor_2046_nl = ~((~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b01)
      | (cfg_proc_precision_1_sva_st_65!=2'b10));
  assign mux_163_nl = MUX_s_1_2_2((nor_2046_nl), nor_2047_cse, or_5189_cse);
  assign FpFloatToInt_16U_5U_10U_shift_and_1_cse = core_wen & (~ and_dcpl_93) & (mux_163_nl);
  assign and_641_rgt = or_5189_cse & (~ IsNaN_8U_23U_land_3_lpi_1_dfm_3);
  assign and_643_rgt = or_5189_cse & (~ IsNaN_8U_23U_land_4_lpi_1_dfm_3);
  assign nor_1099_cse = ~(IsNaN_8U_23U_IsNaN_8U_23U_nand_4_itm_2 | IsNaN_8U_23U_nor_4_itm_2);
  assign and_646_rgt = or_tmp_2469 & or_5189_cse;
  assign nor_2040_cse = ~((~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt);
  assign or_300_cse = (cfg_out_precision_1_sva_st_113!=2'b01);
  assign or_303_cse = nor_2040_cse | (cfg_out_precision_1_sva_st_154!=2'b01) | (~
      main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign or_306_cse = (cfg_out_precision_1_sva_st_154!=2'b01) | (~ main_stage_v_1)
      | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_166_cse = MUX_s_1_2_2(or_tmp_306, or_306_cse, or_5189_cse);
  assign and_648_rgt = or_5189_cse & (~ IsNaN_8U_23U_land_6_lpi_1_dfm_3);
  assign or_309_cse = (cfg_out_precision_1_sva_st_149!=2'b01);
  assign mux_169_nl = MUX_s_1_2_2(mux_166_cse, or_303_cse, or_309_cse);
  assign FpFloatToInt_16U_5U_10U_shift_and_5_cse = core_wen & (~ and_dcpl_93) & (~
      (mux_169_nl));
  assign and_650_rgt = or_5189_cse & (~ IsNaN_8U_23U_land_7_lpi_1_dfm_3);
  assign and_652_rgt = or_5189_cse & (~ IsNaN_8U_23U_land_8_lpi_1_dfm_3);
  assign and_654_rgt = or_5189_cse & (~ IsNaN_8U_23U_land_9_lpi_1_dfm_3);
  assign nor_45_cse = ~((cfg_out_precision_1_sva_st_149!=2'b01));
  assign mux_175_nl = MUX_s_1_2_2(or_303_cse, mux_166_cse, nor_45_cse);
  assign FpFloatToInt_16U_5U_10U_shift_and_8_cse = core_wen & (~ and_dcpl_93) & (~
      (mux_175_nl));
  assign and_656_rgt = or_5189_cse & (~ IsNaN_8U_23U_land_10_lpi_1_dfm_3);
  assign and_658_rgt = or_5189_cse & (~ IsNaN_8U_23U_land_11_lpi_1_dfm_3);
  assign and_660_rgt = or_5189_cse & (~ IsNaN_8U_23U_land_12_lpi_1_dfm_3);
  assign and_662_rgt = or_5189_cse & (~ IsNaN_8U_23U_land_13_lpi_1_dfm_3);
  assign and_664_rgt = or_5189_cse & (~ IsNaN_8U_23U_land_14_lpi_1_dfm_3);
  assign and_666_rgt = or_5189_cse & (~ IsNaN_8U_23U_land_15_lpi_1_dfm_3);
  assign and_668_rgt = or_5189_cse & (~ IsNaN_8U_23U_land_lpi_1_dfm_3);
  assign nor_50_cse = ~((cfg_proc_precision_1_sva_st_65!=2'b10));
  assign nor_2026_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ mux_tmp_200));
  assign mux_201_cse = MUX_s_1_2_2((nor_2026_nl), mux_tmp_200, cfg_proc_precision_1_sva_st_101[0]);
  assign or_400_cse_1 = (cfg_proc_precision_1_sva_st_101!=2'b10);
  assign and_2237_cse = main_stage_v_2 & or_4862_cse;
  assign or_419_cse = (~ cvt_unequal_tmp_19) | cfg_mode_eql_1_sva_4 | (cfg_out_precision_1_sva_st_154!=2'b00);
  assign or_423_cse = (~ cvt_unequal_tmp_20) | cfg_mode_eql_1_sva_5 | (cfg_out_precision_1_sva_st_113!=2'b00);
  assign or_425_cse = (cfg_out_precision_1_sva_st_113!=2'b00);
  assign IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_27_cse =
      and_dcpl_204 | and_dcpl_4;
  assign FpIntToFloat_17U_5U_10U_else_i_abs_and_cse = core_wen & ((or_5189_cse &
      (~ cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_nor_tmp) & ((cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_acc_tmp[16])
      | cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_and_1_tmp)) | and_dcpl_209) &
      (~ mux_tmp_245);
  assign nor_57_cse = ~((cfg_out_precision_1_sva_st_113!=2'b10));
  assign or_451_cse = (~ cvt_unequal_tmp_20) | cfg_mode_eql_1_sva_5;
  assign and_676_cse = and_tmp_12 & or_5189_cse;
  assign IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse =
      and_676_cse | and_685_rgt;
  assign nor_2011_cse = ~((cfg_out_precision_1_sva_st_154!=2'b00) | (~ mux_tmp_259));
  assign or_461_cse = (cfg_out_precision_1_sva_st_149!=2'b00);
  assign FpIntToFloat_17U_5U_10U_else_i_abs_and_13_cse = core_wen & ((or_5189_cse
      & (~ cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp) & ((cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[16])
      | cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp)) | and_dcpl_217) &
      not_tmp_249;
  assign nor_63_cse = ~((cfg_out_precision_1_sva_st_149!=2'b10));
  assign nor_2004_cse = ~((cfg_out_precision_1_sva_st_154!=2'b10) | (~ and_1386_cse));
  assign nor_2005_cse = ~(nor_2040_cse | (cfg_out_precision_1_sva_st_154!=2'b10)
      | (~ and_1386_cse));
  assign mux_273_nl = MUX_s_1_2_2(and_1078_cse, and_1386_cse, or_5189_cse);
  assign IntShiftRightSat_49U_6U_17U_if_and_cse = core_wen & (~ and_dcpl_93) & (mux_273_nl);
  assign and_685_rgt = or_dcpl_15 & or_5189_cse;
  assign FpIntToFloat_17U_5U_10U_else_i_abs_and_15_cse = core_wen & ((or_5189_cse
      & (~ cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp) & (cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp
      | (cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[16]))) | and_dcpl_224)
      & not_tmp_269;
  assign or_513_cse = (~ cvt_unequal_tmp_19) | cfg_mode_eql_1_sva_4;
  assign nor_1980_cse = ~((cfg_out_precision_1_sva_st_154!=2'b00) | (~ mux_tmp_305));
  assign or_3063_cse = nor_tmp_636 | (cfg_out_precision_1_sva_st_154!=2'b10) | or_dcpl_15;
  assign and_696_nl = and_676_cse & and_dcpl_228 & (~ cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp)
      & or_dcpl_108;
  assign and_699_nl = and_676_cse & or_dcpl_109 & and_dcpl_228;
  assign mux_1750_nl = MUX_s_1_2_2(or_3696_cse, (~ mux_tmp_321), main_stage_v_2);
  assign mux_1751_nl = MUX_s_1_2_2((mux_1750_nl), or_3696_cse, or_5189_cse);
  assign mux_1752_nl = MUX_s_1_2_2(or_3063_cse, (mux_1751_nl), nor_63_cse);
  assign FpIntToFloat_17U_5U_10U_else_if_mux1h_9_rgt = MUX1HOT_v_15_3_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_4_sva[15:1]),
      IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_mx0w0, ({5'b0 , FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_10_itm_mx0w0}),
      {(and_696_nl) , (and_699_nl) , (mux_1752_nl)});
  assign or_4550_cse = (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign and_2257_cse = or_183_cse_1 & or_4550_cse & or_5189_cse & (cfg_out_precision_1_sva_st_154==2'b10)
      & core_wen;
  assign nor_2150_cse = ~((reg_cfg_proc_precision_1_sva_st_40_cse!=2'b10));
  assign or_4559_cse = nor_2150_cse | (cfg_out_precision_1_sva_st_154[0]);
  assign nor_2326_cse = ~((cfg_out_precision_1_sva_st_154[1]) | (~ or_tmp_3763));
  assign mux_2172_nl = MUX_s_1_2_2(nor_2326_cse, or_tmp_3763, or_4559_cse);
  assign mux_2173_nl = MUX_s_1_2_2(or_tmp_3763, (mux_2172_nl), or_183_cse_1);
  assign mux_2174_nl = MUX_s_1_2_2((mux_2173_nl), or_tmp_3763, nor_8_cse);
  assign and_2259_cse = (~((mux_2174_nl) | nor_2040_cse)) & core_wen;
  assign and_704_rgt = or_dcpl_109 & or_5189_cse;
  assign and_2230_cse = main_stage_v_2 & mux_1126_cse;
  assign and_711_nl = and_676_cse & and_dcpl_228 & (~ cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp)
      & or_dcpl_110;
  assign and_714_nl = and_676_cse & or_dcpl_111 & and_dcpl_228;
  assign or_3070_nl = nor_tmp_636 | (cfg_out_precision_1_sva_st_154[0]) | not_tmp_2254;
  assign mux_2170_nl = MUX_s_1_2_2(or_tmp_2960, (~ mux_tmp_455), main_stage_v_2);
  assign mux_1757_nl = MUX_s_1_2_2((mux_2170_nl), or_tmp_2960, or_5189_cse);
  assign mux_1758_nl = MUX_s_1_2_2((mux_1757_nl), (or_3070_nl), or_578_cse);
  assign FpIntToFloat_17U_5U_10U_else_if_mux1h_12_rgt = MUX1HOT_v_15_3_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_5_sva[15:1]),
      IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_mx0w0, ({5'b0 , FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_13_itm_mx0w0}),
      {(and_711_nl) , (and_714_nl) , (mux_1758_nl)});
  assign and_719_rgt = or_dcpl_111 & or_5189_cse;
  assign or_578_cse = (cfg_out_precision_1_sva_st_149!=2'b10);
  assign nor_1958_nl = ~((cfg_proc_precision_1_sva_st_64[1]) | (~ or_183_cse_1));
  assign mux_344_cse = MUX_s_1_2_2((nor_1958_nl), or_183_cse_1, cfg_proc_precision_1_sva_st_64[0]);
  assign and_174_cse = main_stage_v_2 & mux_382_cse;
  assign mux_1760_nl = MUX_s_1_2_2(or_3696_cse, (~ and_tmp_225), main_stage_v_2);
  assign mux_1761_cse = MUX_s_1_2_2((mux_1760_nl), or_3696_cse, or_5189_cse);
  assign mux_1762_cse = MUX_s_1_2_2(or_3063_cse, mux_1761_cse, nor_63_cse);
  assign and_726_nl = and_676_cse & and_dcpl_228 & (~ cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp)
      & or_dcpl_113;
  assign and_729_nl = and_676_cse & or_dcpl_114 & and_dcpl_228;
  assign FpIntToFloat_17U_5U_10U_else_if_mux1h_15_rgt = MUX1HOT_v_15_3_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_6_sva[15:1]),
      IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_mx0w0, ({5'b0 , FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_16_itm_mx0w0}),
      {(and_726_nl) , (and_729_nl) , mux_1762_cse});
  assign mux_2177_nl = MUX_s_1_2_2(nor_2326_cse, or_tmp_3763, cfg_out_precision_1_sva_st_154[0]);
  assign mux_2178_nl = MUX_s_1_2_2((mux_2177_nl), or_tmp_3763, nor_2150_cse);
  assign mux_2179_nl = MUX_s_1_2_2((mux_2178_nl), or_tmp_3763, nor_8_cse);
  assign and_2275_cse = (~((mux_2179_nl) | nor_2040_cse)) & core_wen;
  assign and_734_rgt = or_dcpl_114 & or_5189_cse;
  assign and_178_itm = main_stage_v_2 & and_tmp_79;
  assign mux_378_nl = MUX_s_1_2_2(and_178_itm, and_tmp_19, or_5189_cse);
  assign IntShiftRightSat_49U_6U_17U_if_and_3_cse = core_wen & (~ and_dcpl_93) &
      (mux_378_nl);
  assign or_4536_cse = IntShiftRightSat_49U_6U_17U_lor_8_lpi_1_dfm | cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2;
  assign nor_1939_nl = ~((cfg_proc_precision_1_sva_st_65[1]) | (~ mux_tmp_345));
  assign mux_382_cse = MUX_s_1_2_2((nor_1939_nl), mux_tmp_345, cfg_proc_precision_1_sva_st_65[0]);
  assign and_741_nl = and_676_cse & and_dcpl_228 & (~ cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp)
      & or_dcpl_115;
  assign and_744_nl = and_676_cse & or_dcpl_116 & and_dcpl_228;
  assign FpIntToFloat_17U_5U_10U_else_if_mux1h_18_rgt = MUX1HOT_v_15_3_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_7_sva[15:1]),
      IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_mx0w0, ({5'b0 , FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_19_itm_mx0w0}),
      {(and_741_nl) , (and_744_nl) , mux_1762_cse});
  assign and_749_rgt = or_dcpl_116 & or_5189_cse;
  assign or_4535_cse = IntShiftRightSat_49U_6U_17U_lor_9_lpi_1_dfm | cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_svs_st_2;
  assign nor_1917_nl = ~((cfg_proc_precision_1_sva_st_65[1]) | (~ mux_tmp_416));
  assign mux_417_cse = MUX_s_1_2_2((nor_1917_nl), mux_tmp_416, cfg_proc_precision_1_sva_st_65[0]);
  assign nor_1898_cse = ~((cfg_out_precision_1_sva_st_154!=2'b00) | (~ mux_tmp_435));
  assign and_756_nl = and_676_cse & and_dcpl_228 & (~ cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp)
      & or_dcpl_119;
  assign and_759_nl = and_676_cse & or_dcpl_120 & and_dcpl_228;
  assign mux_1772_nl = MUX_s_1_2_2(mux_1761_cse, or_3063_cse, or_578_cse);
  assign FpIntToFloat_17U_5U_10U_else_if_mux1h_21_rgt = MUX1HOT_v_15_3_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_8_sva[15:1]),
      IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_mx0w0, ({5'b0 , FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_22_itm_mx0w0}),
      {(and_756_nl) , (and_759_nl) , (mux_1772_nl)});
  assign and_766_rgt = or_dcpl_120 & or_5189_cse;
  assign FpIntToFloat_17U_5U_10U_else_i_abs_and_22_cse = core_wen & ((or_5189_cse
      & (~ cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp) & ((cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[16])
      | cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp)) | and_dcpl_301) &
      not_tmp_520;
  assign nor_1875_nl = ~((cfg_proc_precision_1_sva_st_64[1]) | (~ mux_tmp_317));
  assign mux_474_cse = MUX_s_1_2_2((nor_1875_nl), mux_tmp_317, cfg_proc_precision_1_sva_st_64[0]);
  assign mux_2171_nl = MUX_s_1_2_2(or_3696_cse, (~ mux_1142_cse), main_stage_v_2);
  assign mux_1779_cse = MUX_s_1_2_2((mux_2171_nl), or_3696_cse, or_5189_cse);
  assign and_780_nl = and_676_cse & and_dcpl_228 & (~ cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp)
      & or_dcpl_124;
  assign and_783_nl = and_676_cse & or_dcpl_125 & and_dcpl_228;
  assign mux_1780_nl = MUX_s_1_2_2(mux_1779_cse, or_3063_cse, or_578_cse);
  assign FpIntToFloat_17U_5U_10U_else_if_mux1h_27_rgt = MUX1HOT_v_15_3_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_10_sva[15:1]),
      IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_mx0w0, ({5'b0 , FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_28_itm_mx0w0}),
      {(and_780_nl) , (and_783_nl) , (mux_1780_nl)});
  assign and_787_rgt = or_dcpl_125 & or_5189_cse;
  assign and_794_nl = and_676_cse & and_dcpl_228 & (~ cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp)
      & or_dcpl_126;
  assign and_797_nl = and_676_cse & or_dcpl_127 & and_dcpl_228;
  assign mux_1785_nl = MUX_s_1_2_2(or_3063_cse, mux_1779_cse, nor_63_cse);
  assign FpIntToFloat_17U_5U_10U_else_if_mux1h_30_rgt = MUX1HOT_v_15_3_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_11_sva[15:1]),
      IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_mx0w0, ({5'b0 , FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_31_itm_mx0w0}),
      {(and_794_nl) , (and_797_nl) , (mux_1785_nl)});
  assign and_801_rgt = or_dcpl_127 & or_5189_cse;
  assign or_3151_cse = (cfg_out_precision_1_sva_st_149!=2'b10) | (~ mux_1142_cse);
  assign and_808_nl = and_676_cse & and_dcpl_228 & (~ cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp)
      & or_dcpl_130;
  assign and_811_nl = and_676_cse & or_dcpl_131 & and_dcpl_228;
  assign mux_1788_nl = MUX_s_1_2_2(or_3696_cse, or_3151_cse, nor_tmp_636);
  assign FpIntToFloat_17U_5U_10U_else_if_mux1h_33_rgt = MUX1HOT_v_15_3_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_12_sva[15:1]),
      IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_mx0w0, ({5'b0 , FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_34_itm_mx0w0}),
      {(and_808_nl) , (and_811_nl) , (mux_1788_nl)});
  assign nor_2300_nl = ~((cfg_out_precision_1_sva_st_154[1]) | (~ or_tmp_3379));
  assign mux_2193_nl = MUX_s_1_2_2((nor_2300_nl), or_tmp_3379, or_4559_cse);
  assign mux_2195_nl = MUX_s_1_2_2(or_tmp_3379, (mux_2193_nl), or_183_cse_1);
  assign mux_2196_nl = MUX_s_1_2_2((mux_2195_nl), or_tmp_3379, nor_8_cse);
  assign and_2317_cse = (~((mux_2196_nl) | nor_2040_cse)) & core_wen;
  assign and_816_rgt = or_dcpl_131 & or_5189_cse;
  assign and_823_nl = and_676_cse & and_dcpl_228 & (~ cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp)
      & or_dcpl_132;
  assign and_826_nl = and_676_cse & or_dcpl_133 & and_dcpl_228;
  assign nand_51_nl = ~((cfg_out_precision_1_sva_st_149[1]) & (~ or_tmp_3025));
  assign mux_1790_nl = MUX_s_1_2_2(or_3696_cse, (nand_51_nl), nor_tmp_636);
  assign mux_1791_nl = MUX_s_1_2_2((mux_1790_nl), or_3063_cse, nor_151_cse);
  assign FpIntToFloat_17U_5U_10U_else_if_mux1h_36_rgt = MUX1HOT_v_15_3_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_13_sva[15:1]),
      IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_mx0w0, ({5'b0 , FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_37_itm_mx0w0}),
      {(and_823_nl) , (and_826_nl) , (mux_1791_nl)});
  assign and_830_rgt = or_dcpl_133 & or_5189_cse;
  assign IntShiftRightSat_49U_6U_17U_o_and_90_cse = core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
      & mux_tmp_161;
  assign nor_1772_cse = ~((cfg_out_precision_1_sva_st_154!=2'b00) | (~ mux_tmp_634));
  assign FpIntToFloat_17U_5U_10U_not_1_nl = ~ (fsm_output[0]);
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_63_nl = MUX_v_10_2_2(10'b0000000000,
      FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_40_itm_mx0w0, (FpIntToFloat_17U_5U_10U_not_1_nl));
  assign or_3170_nl = (cfg_out_precision_1_sva_st_154[0]) | main_stage_v_2 | not_tmp_270;
  assign mux_1794_nl = MUX_s_1_2_2((or_3170_nl), or_tmp_3032, or_5189_cse);
  assign nand_225_nl = ~(main_stage_v_2 & (cfg_out_precision_1_sva_st_149==2'b10)
      & mux_1142_cse);
  assign mux_1796_nl = MUX_s_1_2_2(not_tmp_270, or_3151_cse, main_stage_v_2);
  assign mux_1797_nl = MUX_s_1_2_2((mux_1796_nl), (nand_225_nl), cfg_out_precision_1_sva_st_154[0]);
  assign mux_1798_nl = MUX_s_1_2_2((mux_1797_nl), or_tmp_3032, or_5189_cse);
  assign mux_1799_nl = MUX_s_1_2_2((mux_1798_nl), (mux_1794_nl), nor_151_cse);
  assign or_4348_nl = (mux_1799_nl) | (fsm_output[0]);
  assign and_840_nl = and_676_cse & and_dcpl_363 & or_dcpl_136 & (~ cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp);
  assign and_843_nl = and_676_cse & and_dcpl_363 & or_dcpl_137;
  assign FpIntToFloat_17U_5U_10U_else_i_abs_mux1h_17_rgt = MUX1HOT_v_15_3_2(({5'b0
      , (FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_63_nl)}), (FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_14_sva[15:1]),
      IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_mx0w0, {(or_4348_nl) , (and_840_nl)
      , (and_843_nl)});
  assign and_849_rgt = or_dcpl_137 & or_5189_cse;
  assign nor_1761_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ mux_1463_cse));
  assign mux_660_cse = MUX_s_1_2_2((nor_1761_nl), mux_1463_cse, cfg_proc_precision_1_sva_st_101[0]);
  assign and_856_nl = and_676_cse & and_dcpl_228 & (~ cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp)
      & or_dcpl_139;
  assign and_859_nl = and_676_cse & or_dcpl_140 & and_dcpl_228;
  assign or_3196_nl = (cfg_out_precision_1_sva_st_149[0]) | (~((cfg_out_precision_1_sva_st_149[1])
      & and_tmp_225));
  assign mux_1807_nl = MUX_s_1_2_2(or_3696_cse, (or_3196_nl), nor_tmp_636);
  assign mux_1808_nl = MUX_s_1_2_2((mux_1807_nl), or_3063_cse, nor_151_cse);
  assign FpIntToFloat_17U_5U_10U_else_if_mux1h_41_rgt = MUX1HOT_v_15_3_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_15_sva[15:1]),
      IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_mx0w0, ({5'b0 , FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_43_itm_mx0w0}),
      {(and_856_nl) , (and_859_nl) , (mux_1808_nl)});
  assign and_866_rgt = or_dcpl_140 & or_5189_cse;
  assign and_873_nl = and_676_cse & and_dcpl_228 & (~ cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_nor_20_tmp)
      & or_dcpl_143;
  assign and_876_nl = and_676_cse & or_dcpl_144 & and_dcpl_228;
  assign or_3220_nl = main_stage_v_2 | (cfg_out_precision_1_sva_st_154!=2'b10) |
      or_dcpl_15;
  assign mux_1814_nl = MUX_s_1_2_2(or_3696_cse, (~ mux_tmp_1813), main_stage_v_2);
  assign mux_1815_nl = MUX_s_1_2_2((mux_1814_nl), (or_3220_nl), or_578_cse);
  assign mux_1816_nl = MUX_s_1_2_2((mux_1815_nl), or_3696_cse, or_5189_cse);
  assign mux_1817_nl = MUX_s_1_2_2((mux_1816_nl), or_3063_cse, nor_151_cse);
  assign FpIntToFloat_17U_5U_10U_else_if_mux1h_44_rgt = MUX1HOT_v_15_3_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_sva[15:1]),
      IntShiftRightSat_49U_6U_17U_o_15_1_sva_mx0w0, ({5'b0 , FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_46_itm_mx0w0}),
      {(and_873_nl) , (and_876_nl) , (mux_1817_nl)});
  assign and_881_rgt = or_dcpl_144 & or_5189_cse;
  assign nor_1683_nl = ~((cfg_proc_precision_1_sva_st_89[1]) | (~ mux_tmp_766));
  assign mux_767_cse = MUX_s_1_2_2((nor_1683_nl), mux_tmp_766, cfg_proc_precision_1_sva_st_89[0]);
  assign nor_1674_nl = ~((cfg_proc_precision_1_sva_st_89[1]) | (~ mux_tmp_765));
  assign mux_786_cse_1 = MUX_s_1_2_2((nor_1674_nl), mux_tmp_765, cfg_proc_precision_1_sva_st_89[0]);
  assign nor_151_cse = ~((cfg_proc_precision_1_sva_st_101!=2'b10));
  assign mux_796_nl = MUX_s_1_2_2(and_tmp_94, and_1386_cse, or_5189_cse);
  assign cfg_proc_precision_and_24_cse = core_wen & (~ and_dcpl_93) & (mux_796_nl);
  assign mux_800_nl = MUX_s_1_2_2(and_2237_cse, and_tmp_11, or_5189_cse);
  assign cfg_proc_precision_and_27_cse = core_wen & (~ and_dcpl_93) & (mux_800_nl);
  assign FpFloatToInt_16U_5U_10U_internal_int_and_cse = core_wen & (and_dcpl_407
      | and_dcpl_409 | and_dcpl_411);
  assign nor_1056_cse = ~((~ cvt_1_FpFloatToInt_16U_5U_10U_if_acc_itm_11_1) | (cfg_out_precision_1_sva_st_149!=2'b01));
  assign nor_1672_cse = ~((cfg_proc_precision_1_sva_st_66!=2'b10));
  assign or_1157_cse = (cfg_out_precision_1_sva_6!=2'b01);
  assign nor_1666_cse = ~((~ main_stage_v_2) | cfg_mode_eql_1_sva_5);
  assign nor_1669_cse = ~((cfg_out_precision_1_sva_st_113!=2'b01) | (~ main_stage_v_2)
      | cfg_mode_eql_1_sva_5);
  assign or_1159_cse = (cfg_proc_precision_1_sva_st_66!=2'b10);
  assign and_896_rgt = ((~ cvt_1_FpFloatToInt_16U_5U_10U_if_acc_itm_11_1) | (cfg_out_precision_1_sva_st_149[1])
      | (cfg_proc_precision_1_sva_st_65[0]) | nand_219_cse) & and_dcpl_408;
  assign and_900_rgt = nor_1056_cse & (cfg_proc_precision_1_sva_st_65[1]) & and_dcpl_417;
  assign nor_1664_cse = ~((cfg_proc_precision_1_sva_st_65!=2'b10) | (cfg_out_precision_1_sva_st_113!=2'b01));
  assign or_1176_cse = (cfg_out_precision_1_sva_6!=2'b01) | cfg_mode_eql_1_sva_6;
  assign mux_813_cse = MUX_s_1_2_2(cfg_mode_eql_1_sva_6, or_1176_cse, nor_1672_cse);
  assign nor_1659_nl = ~((cfg_out_precision_1_sva_st_113!=2'b01) | (~ main_stage_v_2)
      | cvt_unequal_tmp_20 | cfg_mode_eql_1_sva_5);
  assign mux_816_nl = MUX_s_1_2_2(nor_1626_cse, (nor_1659_nl), nor_50_cse);
  assign nor_1661_nl = ~((cfg_out_precision_1_sva_6!=2'b01) | (~ main_stage_v_3)
      | cvt_unequal_tmp_21 | cfg_mode_eql_1_sva_6);
  assign mux_817_nl = MUX_s_1_2_2(nor_1630_cse, (nor_1661_nl), nor_1672_cse);
  assign mux_818_nl = MUX_s_1_2_2((mux_817_nl), (mux_816_nl), or_5189_cse);
  assign FpFloatToInt_16U_5U_10U_if_and_cse = core_wen & (~ and_dcpl_93) & (mux_818_nl);
  assign IsNaN_5U_10U_aelse_or_cse = ((~ or_4862_cse) & or_5189_cse) | and_dcpl_424;
  assign IsNaN_5U_10U_aelse_and_cse = core_wen & IsNaN_5U_10U_aelse_or_cse;
  assign or_1196_cse = cvt_unequal_tmp_20 | (cfg_out_precision_1_sva_st_113!=2'b01);
  assign or_1202_cse = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_16!=5'b00000);
  assign nand_207_cse = ~((cfg_out_precision_1_sva_6[1]) & or_1159_cse);
  assign mux_827_cse = MUX_s_1_2_2(or_1159_cse, (~ or_1159_cse), or_1157_cse);
  assign or_1198_cse = (cfg_out_precision_1_sva_st_113!=2'b10);
  assign nor_2099_cse = ~(cvt_unequal_tmp_20 | nor_2285_cse);
  assign nor_213_cse = ~((cfg_proc_precision_1_sva_st_90!=2'b10));
  assign nl_cvt_2_FpMantRNE_17U_11U_else_acc_1_nl = (FpIntToFloat_17U_5U_10U_else_int_mant_2_sva[15:6])
      + conv_u2u_1_10(FpMantRNE_17U_11U_else_carry_2_sva);
  assign cvt_2_FpMantRNE_17U_11U_else_acc_1_nl = nl_cvt_2_FpMantRNE_17U_11U_else_acc_1_nl[9:0];
  assign FpIntToFloat_17U_5U_10U_if_not_179_nl = ~ cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_4_nl = MUX_v_10_2_2(10'b0000000000,
      (cvt_2_FpMantRNE_17U_11U_else_acc_1_nl), (FpIntToFloat_17U_5U_10U_if_not_179_nl));
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_1_nl = MUX_v_10_2_2((FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_4_nl),
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_6_lpi_1_dfm_8, and_dcpl_408);
  assign FpFloatToInt_16U_5U_10U_and_33_nl = (~ (chn_idata_data_sva_2_79_63_1[0]))
      & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_1_m1c & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_34_nl = (chn_idata_data_sva_2_79_63_1[0]) &
      FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_1_m1c & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_3_nl = cvt_2_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1
      & (~ IsNaN_5U_10U_land_2_lpi_1_dfm_mx0w0) & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_nl = IsNaN_5U_10U_land_2_lpi_1_dfm_mx0w0
      & and_dcpl_433;
  assign and_916_nl = (or_dcpl_151 | (cfg_out_precision_1_sva_st_113[0])) & and_dcpl_420;
  assign and_921_nl = and_tmp_50 & (cfg_out_precision_1_sva_st_113==2'b00) & cvt_unequal_tmp_20
      & or_5189_cse;
  assign nor_2100_nl = ~(nor_2219_cse | (cfg_out_precision_1_sva_st_113!=2'b10));
  assign mux_1828_nl = MUX_s_1_2_2((nor_2100_nl), nor_2099_cse, nor_50_cse);
  assign nor_2101_nl = ~(nor_213_cse | (cfg_out_precision_1_sva_6[0]) | nand_207_cse);
  assign mux_1830_nl = MUX_s_1_2_2(mux_827_cse, (nor_2101_nl), cvt_unequal_tmp_21);
  assign mux_1831_nl = MUX_s_1_2_2((mux_1830_nl), (mux_1828_nl), or_5189_cse);
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_1_rgt = MUX1HOT_v_15_7_2((FpFloatToInt_16U_5U_10U_internal_int_24_1_2_sva[14:0]),
      (FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_2_sva[15:1]), (FpFloatToInt_16U_5U_10U_if_qr_2_lpi_1_dfm_mx0[15:1]),
      15'b100000000000000, IntSaturation_17U_16U_o_15_1_2_lpi_1_dfm_6, IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_2,
      ({5'b0 , (FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_1_nl)}), {(FpFloatToInt_16U_5U_10U_and_33_nl)
      , (FpFloatToInt_16U_5U_10U_and_34_nl) , (FpFloatToInt_16U_5U_10U_and_3_nl)
      , (FpFloatToInt_16U_5U_10U_o_int_and_nl) , (and_916_nl) , (and_921_nl) , (mux_1831_nl)});
  assign nor_2285_cse = ~((cfg_out_precision_1_sva_st_113!=2'b01));
  assign or_4709_cse = cvt_unequal_tmp_20 | nor_2285_cse;
  assign nor_2219_cse = ~((cfg_proc_precision_1_sva_st_89!=2'b10));
  assign and_2360_cse = (cfg_proc_precision_1_sva_st_65==2'b10);
  assign or_4714_cse = (cfg_proc_precision_1_sva_st_89!=2'b10);
  assign IsNaN_5U_10U_aelse_or_1_cse = and_dcpl_408 | and_dcpl_420;
  assign IsNaN_5U_10U_aelse_and_1_cse = core_wen & IsNaN_5U_10U_aelse_or_1_cse;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_2_nl = MUX_v_10_2_2(FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_10_itm_mx0w0,
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_10_lpi_1_dfm_8, and_dcpl_408);
  assign FpFloatToInt_16U_5U_10U_and_35_nl = (~ (chn_idata_data_sva_2_111_95_1[0]))
      & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_2_m1c & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_36_nl = (chn_idata_data_sva_2_111_95_1[0]) &
      FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_2_m1c & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_5_nl = cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1
      & (~ IsNaN_5U_10U_land_3_lpi_1_dfm_4) & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_29_nl = IsNaN_5U_10U_land_3_lpi_1_dfm_4
      & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_2_rgt = MUX1HOT_v_15_7_2((FpFloatToInt_16U_5U_10U_internal_int_24_1_3_sva[14:0]),
      (FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_3_sva[15:1]), (FpFloatToInt_16U_5U_10U_if_qr_3_lpi_1_dfm_mx0[15:1]),
      15'b100000000000000, IntSaturation_17U_16U_o_15_1_3_lpi_1_dfm_6, IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_2,
      ({5'b0 , (FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_2_nl)}), {(FpFloatToInt_16U_5U_10U_and_35_nl)
      , (FpFloatToInt_16U_5U_10U_and_36_nl) , (FpFloatToInt_16U_5U_10U_and_5_nl)
      , (FpFloatToInt_16U_5U_10U_o_int_and_29_nl) , and_dcpl_425 , and_dcpl_446 ,
      not_tmp_2422});
  assign nor_2284_nl = ~((cfg_proc_precision_1_sva_st_65[0]) | (~((cfg_proc_precision_1_sva_st_65[1])
      & cvt_unequal_tmp_20)));
  assign mux_2225_nl = MUX_s_1_2_2((nor_2284_nl), cvt_unequal_tmp_20, cfg_out_precision_1_sva_st_113[0]);
  assign or_4718_nl = (~((~ (cfg_out_precision_1_sva_st_113[0])) | (cfg_proc_precision_1_sva_st_65!=2'b10)))
      | cvt_unequal_tmp_20;
  assign mux_2226_nl = MUX_s_1_2_2((or_4718_nl), (mux_2225_nl), cfg_out_precision_1_sva_st_113[1]);
  assign and_2365_cse = (mux_2226_nl) & or_5189_cse & core_wen;
  assign and_2369_cse = (and_2360_cse | cvt_unequal_tmp_20 | ((cfg_out_precision_1_sva_st_113==2'b10)))
      & or_5189_cse & core_wen;
  assign nor_1049_nl = ~(nor_1589_cse | nor_183_cse | nor_213_cse | (cfg_out_precision_1_sva_6[0])
      | nand_207_cse);
  assign mux_1851_cse = MUX_s_1_2_2(mux_827_cse, (nor_1049_nl), cvt_unequal_tmp_21);
  assign nor_1048_cse = ~(nor_2219_cse | nor_151_cse | (cfg_out_precision_1_sva_st_113!=2'b10));
  assign mux_1849_cse = MUX_s_1_2_2(nor_1048_cse, nor_2099_cse, nor_50_cse);
  assign mux_1852_cse = MUX_s_1_2_2(mux_1851_cse, mux_1849_cse, or_5189_cse);
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_3_nl = MUX_v_10_2_2(FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_46_itm_mx0w0,
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_8_lpi_1_dfm_8, and_dcpl_408);
  assign FpFloatToInt_16U_5U_10U_and_61_nl = (~ chn_idata_data_sva_2_511_1) & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_15_m1c
      & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_62_nl = chn_idata_data_sva_2_511_1 & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_15_m1c
      & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_31_nl = cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_itm_11_1
      & (~ IsNaN_5U_10U_land_lpi_1_dfm_4) & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_27_nl = IsNaN_5U_10U_land_lpi_1_dfm_4
      & and_dcpl_433;
  assign and_945_nl = ((~ and_tmp_225) | (cfg_out_precision_1_sva_st_113[0])) & and_dcpl_420;
  assign and_949_nl = mux_tmp_1813 & or_5189_cse & and_dcpl_458;
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_4_rgt = MUX1HOT_v_15_7_2((FpFloatToInt_16U_5U_10U_internal_int_24_1_sva[14:0]),
      (FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_sva[15:1]), (FpFloatToInt_16U_5U_10U_if_qr_lpi_1_dfm_mx0[15:1]),
      15'b100000000000000, IntSaturation_17U_16U_o_15_1_lpi_1_dfm_9, IntShiftRightSat_49U_6U_17U_o_15_1_sva_2,
      ({5'b0 , (FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_3_nl)}), {(FpFloatToInt_16U_5U_10U_and_61_nl)
      , (FpFloatToInt_16U_5U_10U_and_62_nl) , (FpFloatToInt_16U_5U_10U_and_31_nl)
      , (FpFloatToInt_16U_5U_10U_o_int_and_27_nl) , (and_945_nl) , (and_949_nl) ,
      mux_1852_cse});
  assign and_2371_nl = cvt_unequal_tmp_20 & (nor_2219_cse | nor_151_cse | (cfg_out_precision_1_sva_st_113!=2'b10));
  assign mux_2227_nl = MUX_s_1_2_2((and_2371_nl), or_4709_cse, nor_50_cse);
  assign and_2372_cse = (mux_2227_nl) & or_5189_cse & core_wen;
  assign and_2380_cse = ((or_4714_cse & (cfg_out_precision_1_sva_st_113==2'b10) &
      or_400_cse_1) | and_2360_cse | cvt_unequal_tmp_20) & or_5189_cse & core_wen;
  assign and_2156_nl = cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1 & nor_2285_cse;
  assign mux_1859_nl = MUX_s_1_2_2((~ or_4862_cse), or_4862_cse, and_2156_nl);
  assign and_954_rgt = (mux_1859_nl) & and_dcpl_408;
  assign and_956_rgt = cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1 & (cfg_proc_precision_1_sva_st_65[1])
      & and_dcpl_417;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_4_nl = MUX_v_10_2_2(FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_13_itm_mx0w0,
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_11_lpi_1_dfm_8, and_dcpl_408);
  assign FpFloatToInt_16U_5U_10U_and_39_nl = (~ (chn_idata_data_sva_2_175_159_1[0]))
      & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_4_m1c & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_40_nl = (chn_idata_data_sva_2_175_159_1[0])
      & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_4_m1c & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_9_nl = cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1
      & (~ IsNaN_5U_10U_land_5_lpi_1_dfm_4) & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_26_nl = IsNaN_5U_10U_land_5_lpi_1_dfm_4
      & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_5_rgt = MUX1HOT_v_15_7_2((FpFloatToInt_16U_5U_10U_internal_int_24_1_5_sva[14:0]),
      (FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_5_sva[15:1]), (FpFloatToInt_16U_5U_10U_if_qr_5_lpi_1_dfm_mx0[15:1]),
      15'b100000000000000, IntSaturation_17U_16U_o_15_1_5_lpi_1_dfm_6, IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_2,
      ({5'b0 , (FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_4_nl)}), {(FpFloatToInt_16U_5U_10U_and_39_nl)
      , (FpFloatToInt_16U_5U_10U_and_40_nl) , (FpFloatToInt_16U_5U_10U_and_9_nl)
      , (FpFloatToInt_16U_5U_10U_o_int_and_26_nl) , and_dcpl_425 , and_dcpl_446 ,
      not_tmp_2422});
  assign nor_1624_cse = ~(chn_idata_data_sva_2_511_1 | (~ main_stage_v_2) | cvt_unequal_tmp_20
      | cfg_mode_eql_1_sva_5);
  assign nor_1630_cse = ~((~ main_stage_v_3) | cvt_unequal_tmp_21 | cfg_mode_eql_1_sva_6);
  assign nor_1629_cse = ~((cfg_out_precision_1_sva_6!=2'b01));
  assign nor_1626_cse = ~((~ main_stage_v_2) | cvt_unequal_tmp_20 | cfg_mode_eql_1_sva_5);
  assign and_957_rgt = or_dcpl_147 & or_5189_cse;
  assign nor_1040_nl = ~(nor_2219_cse | nor_151_cse | (~ (cfg_out_precision_1_sva_st_149[1]))
      | (cfg_out_precision_1_sva_st_113!=2'b10));
  assign mux_1864_cse = MUX_s_1_2_2((nor_1040_nl), nor_2099_cse, nor_50_cse);
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_5_nl = MUX_v_10_2_2(FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_43_itm_mx0w0,
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_7_lpi_1_dfm_8, and_dcpl_408);
  assign FpFloatToInt_16U_5U_10U_and_59_nl = (~ (chn_idata_data_sva_2_495_479_1[0]))
      & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_14_m1c & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_60_nl = (chn_idata_data_sva_2_495_479_1[0])
      & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_14_m1c & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_29_nl = cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1
      & (~ IsNaN_5U_10U_land_15_lpi_1_dfm_mx0w0) & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_25_nl = IsNaN_5U_10U_land_15_lpi_1_dfm_mx0w0
      & and_dcpl_433;
  assign and_961_nl = ((~ and_tmp_225) | or_dcpl_160) & and_dcpl_420;
  assign and_966_nl = and_dcpl_473 & (~ (cfg_out_precision_1_sva_st_149[1])) & (~
      (cfg_out_precision_1_sva_st_113[0])) & cvt_unequal_tmp_20;
  assign mux_1867_nl = MUX_s_1_2_2(mux_1851_cse, mux_1864_cse, or_5189_cse);
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_6_rgt = MUX1HOT_v_15_7_2((FpFloatToInt_16U_5U_10U_internal_int_24_1_15_sva[14:0]),
      (FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_15_sva[15:1]), (FpFloatToInt_16U_5U_10U_if_qr_15_lpi_1_dfm_mx0[15:1]),
      15'b100000000000000, IntSaturation_17U_16U_o_15_1_15_lpi_1_dfm_8, IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_2,
      ({5'b0 , (FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_5_nl)}), {(FpFloatToInt_16U_5U_10U_and_59_nl)
      , (FpFloatToInt_16U_5U_10U_and_60_nl) , (FpFloatToInt_16U_5U_10U_and_29_nl)
      , (FpFloatToInt_16U_5U_10U_o_int_and_25_nl) , (and_961_nl) , (and_966_nl) ,
      (mux_1867_nl)});
  assign or_4745_nl = cvt_unequal_tmp_20 | (cfg_out_precision_1_sva_st_113[0]);
  assign mux_2230_cse = MUX_s_1_2_2((or_4745_nl), cvt_unequal_tmp_20, cfg_out_precision_1_sva_st_113[1]);
  assign or_4749_cse = nor_2219_cse | nor_151_cse | (~ (cfg_out_precision_1_sva_st_149[1]))
      | (cfg_out_precision_1_sva_st_113[0]);
  assign and_2388_cse = cvt_unequal_tmp_20 & or_4749_cse;
  assign mux_2231_nl = MUX_s_1_2_2(and_2388_cse, mux_2230_cse, nor_50_cse);
  assign and_2389_cse = (mux_2231_nl) & or_5189_cse & core_wen;
  assign or_4755_nl = cvt_unequal_tmp_20 | (~ or_4749_cse);
  assign mux_2232_nl = MUX_s_1_2_2(and_2388_cse, (or_4755_nl), cfg_out_precision_1_sva_st_113[1]);
  assign and_2393_cse = ((mux_2232_nl) | and_2360_cse) & or_5189_cse & core_wen;
  assign and_976_cse = (or_dcpl_163 | and_1021_cse | (cfg_out_precision_1_sva_st_113[0]))
      & and_dcpl_420;
  assign and_978_cse = and_tmp_225 & and_dcpl_481;
  assign nor_1033_nl = ~(nor_183_cse | nor_213_cse | (cfg_out_precision_1_sva_6[0])
      | nand_207_cse);
  assign mux_1881_cse = MUX_s_1_2_2(mux_827_cse, (nor_1033_nl), cvt_unequal_tmp_21);
  assign mux_1882_cse = MUX_s_1_2_2(mux_1881_cse, mux_1849_cse, or_5189_cse);
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_6_nl = MUX_v_10_2_2(FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_16_itm_mx0w0,
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_12_lpi_1_dfm_8, and_dcpl_408);
  assign FpFloatToInt_16U_5U_10U_and_41_nl = (~ (chn_idata_data_sva_2_207_191_1[0]))
      & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_5_m1c & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_42_nl = (chn_idata_data_sva_2_207_191_1[0])
      & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_5_m1c & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_11_nl = cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1
      & (~ IsNaN_5U_10U_land_6_lpi_1_dfm_4) & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_24_nl = IsNaN_5U_10U_land_6_lpi_1_dfm_4
      & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_7_rgt = MUX1HOT_v_15_7_2((FpFloatToInt_16U_5U_10U_internal_int_24_1_6_sva[14:0]),
      (FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_6_sva[15:1]), (FpFloatToInt_16U_5U_10U_if_qr_6_lpi_1_dfm_mx0[15:1]),
      15'b100000000000000, IntSaturation_17U_16U_o_15_1_6_lpi_1_dfm_7, IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_2,
      ({5'b0 , (FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_6_nl)}), {(FpFloatToInt_16U_5U_10U_and_41_nl)
      , (FpFloatToInt_16U_5U_10U_and_42_nl) , (FpFloatToInt_16U_5U_10U_and_11_nl)
      , (FpFloatToInt_16U_5U_10U_o_int_and_24_nl) , and_976_cse , and_978_cse , mux_1882_cse});
  assign and_2395_nl = cvt_unequal_tmp_20 & (~(or_4714_cse & (~(nor_151_cse | (cfg_out_precision_1_sva_st_113!=2'b10)))));
  assign mux_2233_nl = MUX_s_1_2_2((and_2395_nl), or_4709_cse, nor_50_cse);
  assign and_2396_cse = (mux_2233_nl) & or_5189_cse & core_wen;
  assign and_2402_cse = ((or_400_cse_1 & (cfg_out_precision_1_sva_st_113[1]) & (~(nor_2219_cse
      | (cfg_out_precision_1_sva_st_113[0])))) | and_2360_cse | cvt_unequal_tmp_20)
      & or_5189_cse & core_wen;
  assign and_2154_nl = cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1 & nor_45_cse;
  assign mux_1886_nl = MUX_s_1_2_2((~ or_4862_cse), or_4862_cse, and_2154_nl);
  assign and_984_rgt = (mux_1886_nl) & and_dcpl_408;
  assign and_986_rgt = cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1 & (cfg_proc_precision_1_sva_st_65[1])
      & and_dcpl_417;
  assign FpFloatToInt_16U_5U_10U_and_57_nl = (~ (chn_idata_data_sva_2_463_447_1[0]))
      & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_13_m1c & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_58_nl = (chn_idata_data_sva_2_463_447_1[0])
      & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_13_m1c & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_27_nl = cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1
      & (~ IsNaN_5U_10U_land_14_lpi_1_dfm_5) & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_23_nl = IsNaN_5U_10U_land_14_lpi_1_dfm_5
      & and_dcpl_433;
  assign mux_1888_nl = MUX_s_1_2_2(or_4862_cse, (~ or_4862_cse), nor_2285_cse);
  assign nor_2142_nl = ~(cvt_unequal_tmp_20 | (mux_1888_nl));
  assign mux_1832_nl = MUX_s_1_2_2((~ or_1159_cse), or_1159_cse, or_1157_cse);
  assign nor_2143_nl = ~(cvt_unequal_tmp_21 | (mux_1832_nl));
  assign mux_1889_nl = MUX_s_1_2_2((nor_2143_nl), (nor_2142_nl), or_5189_cse);
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_8_rgt = MUX1HOT_v_15_6_2((FpFloatToInt_16U_5U_10U_internal_int_24_1_14_sva[14:0]),
      (FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_14_sva[15:1]), (FpFloatToInt_16U_5U_10U_if_qr_14_lpi_1_dfm_mx0[15:1]),
      15'b100000000000000, IntSaturation_17U_16U_o_15_1_14_lpi_1_dfm_8, ({5'b0 ,
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_lpi_1_dfm_9}), {(FpFloatToInt_16U_5U_10U_and_57_nl)
      , (FpFloatToInt_16U_5U_10U_and_58_nl) , (FpFloatToInt_16U_5U_10U_and_27_nl)
      , (FpFloatToInt_16U_5U_10U_o_int_and_23_nl) , and_dcpl_420 , (mux_1889_nl)});
  assign and_2153_nl = cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1 & nor_45_cse;
  assign mux_1892_nl = MUX_s_1_2_2((~ or_4862_cse), or_4862_cse, and_2153_nl);
  assign and_987_rgt = (mux_1892_nl) & and_dcpl_408;
  assign and_989_rgt = cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1 & (cfg_proc_precision_1_sva_st_65[1])
      & and_dcpl_417;
  assign nor_183_cse = ~((cfg_proc_precision_1_sva_st_102!=2'b10));
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_7_nl = MUX_v_10_2_2(FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_19_itm_mx0w0,
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_13_lpi_1_dfm_8, and_dcpl_408);
  assign FpFloatToInt_16U_5U_10U_and_43_nl = (~ (chn_idata_data_sva_2_239_223_1[0]))
      & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_6_m1c & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_44_nl = (chn_idata_data_sva_2_239_223_1[0])
      & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_6_m1c & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_13_nl = cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1
      & (~ IsNaN_5U_10U_land_7_lpi_1_dfm_5) & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_22_nl = IsNaN_5U_10U_land_7_lpi_1_dfm_5
      & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_9_rgt = MUX1HOT_v_15_7_2((FpFloatToInt_16U_5U_10U_internal_int_24_1_7_sva[14:0]),
      (FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_7_sva[15:1]), (FpFloatToInt_16U_5U_10U_if_qr_7_lpi_1_dfm_mx0[15:1]),
      15'b100000000000000, IntSaturation_17U_16U_o_15_1_7_lpi_1_dfm_7, IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_2,
      ({5'b0 , (FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_7_nl)}), {(FpFloatToInt_16U_5U_10U_and_43_nl)
      , (FpFloatToInt_16U_5U_10U_and_44_nl) , (FpFloatToInt_16U_5U_10U_and_13_nl)
      , (FpFloatToInt_16U_5U_10U_o_int_and_22_nl) , and_976_cse , and_978_cse , mux_1882_cse});
  assign nor_1589_cse = ~((cfg_proc_precision_1_sva_st_108!=2'b10));
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_8_nl = MUX_v_10_2_2(FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_37_itm_mx0w0,
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_5_lpi_1_dfm_8, and_dcpl_408);
  assign FpFloatToInt_16U_5U_10U_and_55_nl = (~ (chn_idata_data_sva_2_431_415_1[0]))
      & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_12_m1c & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_56_nl = (chn_idata_data_sva_2_431_415_1[0])
      & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_12_m1c & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_25_nl = cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1
      & (~ IsNaN_5U_10U_land_13_lpi_1_dfm_4) & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_21_nl = IsNaN_5U_10U_land_13_lpi_1_dfm_4
      & and_dcpl_433;
  assign and_999_nl = ((~ mux_tmp_455) | or_dcpl_160) & and_dcpl_420;
  assign and_1004_nl = and_dcpl_499 & (~ (cfg_out_precision_1_sva_st_149[1])) & (~
      (cfg_out_precision_1_sva_st_113[0])) & cvt_unequal_tmp_20 & or_400_cse_1;
  assign mux_1909_nl = MUX_s_1_2_2(mux_1881_cse, mux_1864_cse, or_5189_cse);
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_10_rgt = MUX1HOT_v_15_7_2((FpFloatToInt_16U_5U_10U_internal_int_24_1_13_sva[14:0]),
      (FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_13_sva[15:1]), (FpFloatToInt_16U_5U_10U_if_qr_13_lpi_1_dfm_mx0[15:1]),
      15'b100000000000000, IntSaturation_17U_16U_o_15_1_13_lpi_1_dfm_7, IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_2,
      ({5'b0 , (FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_8_nl)}), {(FpFloatToInt_16U_5U_10U_and_55_nl)
      , (FpFloatToInt_16U_5U_10U_and_56_nl) , (FpFloatToInt_16U_5U_10U_and_25_nl)
      , (FpFloatToInt_16U_5U_10U_o_int_and_21_nl) , (and_999_nl) , (and_1004_nl)
      , (mux_1909_nl)});
  assign nor_2269_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ or_4714_cse));
  assign mux_2236_nl = MUX_s_1_2_2((nor_2269_nl), or_4714_cse, cfg_proc_precision_1_sva_st_101[0]);
  assign or_4788_cse = (cfg_out_precision_1_sva_st_113[0]) | (~((cfg_out_precision_1_sva_st_149[1])
      & (mux_2236_nl)));
  assign and_2422_cse = cvt_unequal_tmp_20 & or_4788_cse;
  assign and_2151_nl = cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1 & nor_45_cse;
  assign mux_1916_nl = MUX_s_1_2_2((~ or_4862_cse), or_4862_cse, and_2151_nl);
  assign and_1009_rgt = (mux_1916_nl) & and_dcpl_408;
  assign and_1011_rgt = cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1 & (cfg_proc_precision_1_sva_st_65[1])
      & and_dcpl_417;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_9_nl = MUX_v_10_2_2(FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_22_itm_mx0w0,
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_14_lpi_1_dfm_8, and_dcpl_408);
  assign FpFloatToInt_16U_5U_10U_and_45_nl = (~ (chn_idata_data_sva_2_271_255_1[0]))
      & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_7_m1c & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_46_nl = (chn_idata_data_sva_2_271_255_1[0])
      & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_7_m1c & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_15_nl = cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1
      & (~ IsNaN_5U_10U_land_8_lpi_1_dfm_4) & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_20_nl = IsNaN_5U_10U_land_8_lpi_1_dfm_4
      & and_dcpl_433;
  assign and_1013_nl = (or_3774_cse | (cfg_out_precision_1_sva_st_113[0])) & and_dcpl_420;
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_11_rgt = MUX1HOT_v_15_7_2((FpFloatToInt_16U_5U_10U_internal_int_24_1_8_sva[14:0]),
      (FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_8_sva[15:1]), (FpFloatToInt_16U_5U_10U_if_qr_8_lpi_1_dfm_mx0[15:1]),
      15'b100000000000000, IntSaturation_17U_16U_o_15_1_8_lpi_1_dfm_8, IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_2,
      ({5'b0 , (FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_9_nl)}), {(FpFloatToInt_16U_5U_10U_and_45_nl)
      , (FpFloatToInt_16U_5U_10U_and_46_nl) , (FpFloatToInt_16U_5U_10U_and_15_nl)
      , (FpFloatToInt_16U_5U_10U_o_int_and_20_nl) , (and_1013_nl) , and_978_cse ,
      mux_1852_cse});
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_10_nl = MUX_v_10_2_2(FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_34_itm_mx0w0,
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_4_lpi_1_dfm_8, and_dcpl_408);
  assign FpFloatToInt_16U_5U_10U_and_53_nl = (~ (chn_idata_data_sva_2_399_383_1[0]))
      & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_11_m1c & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_54_nl = (chn_idata_data_sva_2_399_383_1[0])
      & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_11_m1c & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_23_nl = cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1
      & (~ IsNaN_5U_10U_land_12_lpi_1_dfm_4) & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_19_nl = IsNaN_5U_10U_land_12_lpi_1_dfm_4
      & and_dcpl_433;
  assign and_1023_nl = (or_3817_cse | (cfg_out_precision_1_sva_st_113[0])) & and_dcpl_420;
  assign and_1027_nl = mux_1142_cse & (~ (cfg_out_precision_1_sva_st_149[1])) & (~
      (cfg_out_precision_1_sva_st_113[0])) & cvt_unequal_tmp_20 & or_5189_cse;
  assign and_2149_nl = (cfg_out_precision_1_sva_st_149[1]) & nor_1048_cse;
  assign mux_1930_nl = MUX_s_1_2_2((and_2149_nl), nor_2099_cse, nor_50_cse);
  assign mux_1933_nl = MUX_s_1_2_2(mux_1851_cse, (mux_1930_nl), or_5189_cse);
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_12_rgt = MUX1HOT_v_15_7_2((FpFloatToInt_16U_5U_10U_internal_int_24_1_12_sva[14:0]),
      (FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_12_sva[15:1]), (FpFloatToInt_16U_5U_10U_if_qr_12_lpi_1_dfm_mx0[15:1]),
      15'b100000000000000, IntSaturation_17U_16U_o_15_1_12_lpi_1_dfm_8, IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_2,
      ({5'b0 , (FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_10_nl)}), {(FpFloatToInt_16U_5U_10U_and_53_nl)
      , (FpFloatToInt_16U_5U_10U_and_54_nl) , (FpFloatToInt_16U_5U_10U_and_23_nl)
      , (FpFloatToInt_16U_5U_10U_o_int_and_19_nl) , (and_1023_nl) , (and_1027_nl)
      , (mux_1933_nl)});
  assign nl_cvt_9_FpMantRNE_17U_11U_else_acc_1_nl = (FpIntToFloat_17U_5U_10U_else_int_mant_9_sva[15:6])
      + conv_u2u_1_10(FpMantRNE_17U_11U_else_carry_9_sva);
  assign cvt_9_FpMantRNE_17U_11U_else_acc_1_nl = nl_cvt_9_FpMantRNE_17U_11U_else_acc_1_nl[9:0];
  assign FpIntToFloat_17U_5U_10U_if_not_200_nl = ~ cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_25_nl = MUX_v_10_2_2(10'b0000000000,
      (cvt_9_FpMantRNE_17U_11U_else_acc_1_nl), (FpIntToFloat_17U_5U_10U_if_not_200_nl));
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_11_nl = MUX_v_10_2_2((FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_25_nl),
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_15_lpi_1_dfm_8, and_dcpl_408);
  assign FpFloatToInt_16U_5U_10U_and_47_nl = (~ (chn_idata_data_sva_2_303_287_1[0]))
      & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_8_m1c & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_48_nl = (chn_idata_data_sva_2_303_287_1[0])
      & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_8_m1c & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_17_nl = cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1
      & (~ IsNaN_5U_10U_land_9_lpi_1_dfm_4) & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_18_nl = IsNaN_5U_10U_land_9_lpi_1_dfm_4
      & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_13_rgt = MUX1HOT_v_15_7_2((FpFloatToInt_16U_5U_10U_internal_int_24_1_9_sva[14:0]),
      (FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_9_sva[15:1]), (FpFloatToInt_16U_5U_10U_if_qr_9_lpi_1_dfm_mx0[15:1]),
      15'b100000000000000, IntSaturation_17U_16U_o_15_1_9_lpi_1_dfm_6, IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_2,
      ({5'b0 , (FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_11_nl)}), {(FpFloatToInt_16U_5U_10U_and_47_nl)
      , (FpFloatToInt_16U_5U_10U_and_48_nl) , (FpFloatToInt_16U_5U_10U_and_17_nl)
      , (FpFloatToInt_16U_5U_10U_o_int_and_18_nl) , and_dcpl_425 , and_dcpl_446 ,
      not_tmp_2422});
  assign and_1038_cse = ((~ mux_tmp_455) | and_1021_cse | (cfg_out_precision_1_sva_st_113[0]))
      & and_dcpl_420;
  assign and_1039_cse = mux_1142_cse & and_dcpl_481;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_12_nl = MUX_v_10_2_2(FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_31_itm_mx0w0,
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_3_lpi_1_dfm_8, and_dcpl_408);
  assign FpFloatToInt_16U_5U_10U_and_51_nl = (~ (chn_idata_data_sva_2_367_351_1[0]))
      & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_10_m1c & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_52_nl = (chn_idata_data_sva_2_367_351_1[0])
      & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_10_m1c & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_21_nl = cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1
      & (~ IsNaN_5U_10U_land_11_lpi_1_dfm_4) & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_17_nl = IsNaN_5U_10U_land_11_lpi_1_dfm_4
      & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_14_rgt = MUX1HOT_v_15_7_2((FpFloatToInt_16U_5U_10U_internal_int_24_1_11_sva[14:0]),
      (FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_11_sva[15:1]), (FpFloatToInt_16U_5U_10U_if_qr_11_lpi_1_dfm_mx0[15:1]),
      15'b100000000000000, IntSaturation_17U_16U_o_15_1_11_lpi_1_dfm_7, IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_2,
      ({5'b0 , (FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_12_nl)}), {(FpFloatToInt_16U_5U_10U_and_51_nl)
      , (FpFloatToInt_16U_5U_10U_and_52_nl) , (FpFloatToInt_16U_5U_10U_and_21_nl)
      , (FpFloatToInt_16U_5U_10U_o_int_and_17_nl) , and_1038_cse , and_1039_cse ,
      mux_1882_cse});
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_13_nl = MUX_v_10_2_2(FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_28_itm_mx0w0,
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_2_lpi_1_dfm_8, and_dcpl_408);
  assign FpFloatToInt_16U_5U_10U_and_49_nl = (~ (chn_idata_data_sva_2_335_319_1[0]))
      & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_9_m1c & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_50_nl = (chn_idata_data_sva_2_335_319_1[0])
      & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_9_m1c & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_and_19_nl = cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1
      & (~ IsNaN_5U_10U_land_10_lpi_1_dfm_4) & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_and_16_nl = IsNaN_5U_10U_land_10_lpi_1_dfm_4
      & and_dcpl_433;
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_15_rgt = MUX1HOT_v_15_7_2((FpFloatToInt_16U_5U_10U_internal_int_24_1_10_sva[14:0]),
      (FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_10_sva[15:1]), (FpFloatToInt_16U_5U_10U_if_qr_10_lpi_1_dfm_mx0[15:1]),
      15'b100000000000000, IntSaturation_17U_16U_o_15_1_10_lpi_1_dfm_7, IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_2,
      ({5'b0 , (FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_13_nl)}), {(FpFloatToInt_16U_5U_10U_and_49_nl)
      , (FpFloatToInt_16U_5U_10U_and_50_nl) , (FpFloatToInt_16U_5U_10U_and_19_nl)
      , (FpFloatToInt_16U_5U_10U_o_int_and_16_nl) , and_1038_cse , and_1039_cse ,
      mux_1882_cse});
  assign mux_938_nl = MUX_s_1_2_2(main_stage_v_3, main_stage_v_2, or_5189_cse);
  assign cfg_out_precision_and_32_cse = core_wen & (~ and_dcpl_93) & (mux_938_nl);
  assign nor_1556_cse = ~((~ main_stage_v_2) | (~ cvt_unequal_tmp_20) | cfg_mode_eql_1_sva_5);
  assign IntShiftRightSat_49U_6U_17U_o_and_cse = core_wen & (~ and_dcpl_93);
  assign cvt_else_and_cse = core_wen & (~ (fsm_output[0]));
  assign mux_948_nl = MUX_s_1_2_2(mux_tmp_947, mux_tmp_945, or_5189_cse);
  assign cvt_else_and_24_cse = cvt_else_and_cse & (~(or_dcpl_178 | (~ main_stage_v_3)))
      & (~ (mux_948_nl));
  assign reg_cvt_else_cvt_else_nor_4_cse = ~((~ mux_tmp_986) | and_dcpl_535 | (~
      main_stage_v_3));
  assign cvt_else_and_10_cse = core_wen & reg_cvt_else_cvt_else_nor_4_cse;
  assign mux_989_cse = MUX_s_1_2_2(and_1386_cse, mux_1142_cse, main_stage_v_2);
  assign mux_984_nl = MUX_s_1_2_2((~ or_5379_cse), mux_tmp_944, or_183_cse_1);
  assign mux_985_nl = MUX_s_1_2_2((mux_984_nl), mux_1142_cse, main_stage_v_2);
  assign nor_1536_nl = ~((cfg_proc_precision_1_sva_st_108[1]) | (~ mux_tmp_987));
  assign mux_988_nl = MUX_s_1_2_2((nor_1536_nl), mux_tmp_987, cfg_proc_precision_1_sva_st_108[0]);
  assign mux_990_nl = MUX_s_1_2_2(mux_989_cse, (mux_988_nl), main_stage_v_3);
  assign mux_991_nl = MUX_s_1_2_2((mux_990_nl), (mux_985_nl), or_5189_cse);
  assign cvt_else_and_34_cse = cvt_else_and_cse & (~((~ mux_tmp_987) | and_1059_cse
      | (~ main_stage_v_3))) & (~ (mux_991_nl));
  assign cvt_else_and_19_cse = core_wen & (~(or_dcpl_195 | and_1059_cse | (~ main_stage_v_3)));
  assign nor_1523_nl = ~((cfg_out_precision_1_sva_st_113!=2'b00) | (~ main_stage_v_2)
      | (~ cvt_unequal_tmp_20) | cfg_mode_eql_1_sva_5);
  assign mux_1001_nl = MUX_s_1_2_2((nor_1523_nl), nor_1556_cse, nor_50_cse);
  assign nor_1524_nl = ~((~ main_stage_v_3) | (~ cvt_unequal_tmp_21) | cfg_mode_eql_1_sva_6);
  assign nor_1525_nl = ~((cfg_out_precision_1_sva_6!=2'b00) | (~ main_stage_v_3)
      | (~ cvt_unequal_tmp_21) | cfg_mode_eql_1_sva_6);
  assign mux_1002_nl = MUX_s_1_2_2((nor_1525_nl), (nor_1524_nl), nor_1672_cse);
  assign mux_1003_nl = MUX_s_1_2_2((mux_1002_nl), (mux_1001_nl), or_5189_cse);
  assign IntShiftRightSat_49U_6U_17U_o_and_103_cse = core_wen & (~ and_dcpl_93) &
      (mux_1003_nl);
  assign and_1069_m1c = cvt_1_FpMantRNE_17U_11U_else_and_tmp & cvt_unequal_tmp_20
      & or_5189_cse;
  assign nl_cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_nl = (~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_16)
      + 5'b1;
  assign cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_nl = nl_cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_nl[4:0];
  assign FpIntToFloat_17U_5U_10U_o_expo_or_15_nl = ((~ cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_1_itm_4)
      & and_1069_m1c) | ((~ cvt_1_FpMantRNE_17U_11U_else_and_tmp) & cvt_unequal_tmp_20
      & or_5189_cse);
  assign FpIntToFloat_17U_5U_10U_o_expo_and_31_nl = cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_1_itm_4
      & and_1069_m1c;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_1_itm = MUX1HOT_v_5_3_2((~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_16),
      (cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_nl), ({1'b0 , FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_9_3_0_1}),
      {(FpIntToFloat_17U_5U_10U_o_expo_or_15_nl) , (FpIntToFloat_17U_5U_10U_o_expo_and_31_nl)
      , (~ mux_1966_itm)});
  assign or_4862_cse = (cfg_proc_precision_1_sva_st_65!=2'b10);
  assign or_1587_cse = (~ cvt_unequal_tmp_20) | (cfg_out_precision_1_sva_st_113!=2'b10)
      | cfg_mode_eql_1_sva_5;
  assign or_3538_cse = (cfg_proc_precision_1_sva_st_90!=2'b10);
  assign and_1078_cse = main_stage_v_2 & and_tmp_50;
  assign and_1077_rgt = (or_dcpl_151 | (~ main_stage_v_2)) & or_1159_cse & or_3538_cse
      & and_dcpl_103;
  assign and_1080_m1c = or_5189_cse & cvt_unequal_tmp_20 & cvt_2_FpMantRNE_17U_11U_else_and_1_tmp;
  assign or_1596_cse = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_17!=5'b00000);
  assign nl_cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl = (~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_17)
      + 5'b1;
  assign cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl = nl_cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl[4:0];
  assign FpIntToFloat_17U_5U_10U_o_expo_or_14_nl = ((~ cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4)
      & and_1080_m1c) | (or_5189_cse & cvt_unequal_tmp_20 & (~ cvt_2_FpMantRNE_17U_11U_else_and_1_tmp));
  assign FpIntToFloat_17U_5U_10U_o_expo_and_29_nl = cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4
      & and_1080_m1c;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_3_itm = MUX1HOT_v_5_3_2((~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_17),
      (cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl), ({1'b0 , FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_9_3_0_1}),
      {(FpIntToFloat_17U_5U_10U_o_expo_or_14_nl) , (FpIntToFloat_17U_5U_10U_o_expo_and_29_nl)
      , (~ mux_1966_itm)});
  assign nor_1500_cse = ~(nor_213_cse | nor_1672_cse | (~ main_stage_v_3) | (~ cvt_unequal_tmp_21)
      | cfg_mode_eql_1_sva_6 | (cfg_out_precision_1_sva_6!=2'b10) | (cfg_out_precision_1_sva_st_144!=2'b10));
  assign nor_1498_nl = ~(nor_2219_cse | (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | (~ cvt_unequal_tmp_20) | cfg_mode_eql_1_sva_5 | (cfg_out_precision_1_sva_st_113!=2'b10)
      | nor_50_cse);
  assign mux_1027_nl = MUX_s_1_2_2(nor_1500_cse, (nor_1498_nl), or_5189_cse);
  assign FpIntToFloat_17U_5U_10U_is_inf_and_14_cse = core_wen & (~ and_dcpl_93) &
      (mux_1027_nl);
  assign and_1084_m1c = or_5189_cse & cvt_unequal_tmp_20 & cvt_3_FpMantRNE_17U_11U_else_and_1_tmp;
  assign or_1625_cse = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_18!=5'b00000);
  assign nl_cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl = (~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_18)
      + 5'b1;
  assign cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl = nl_cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl[4:0];
  assign FpIntToFloat_17U_5U_10U_o_expo_or_13_nl = ((~ cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4)
      & and_1084_m1c) | (or_5189_cse & cvt_unequal_tmp_20 & (~ cvt_3_FpMantRNE_17U_11U_else_and_1_tmp));
  assign FpIntToFloat_17U_5U_10U_o_expo_and_27_nl = cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4
      & and_1084_m1c;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_5_itm = MUX1HOT_v_5_3_2((~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_18),
      (cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl), ({1'b0 , FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_9_3_0_1}),
      {(FpIntToFloat_17U_5U_10U_o_expo_or_13_nl) , (FpIntToFloat_17U_5U_10U_o_expo_and_27_nl)
      , (~ mux_1966_itm)});
  assign nor_1488_cse = ~((~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt
      | (~ main_stage_v_3) | (cfg_out_precision_1_sva_st_144!=2'b00) | (~ mux_tmp_986));
  assign nor_1489_cse = ~((~ main_stage_v_3) | (cfg_out_precision_1_sva_st_144!=2'b00)
      | (~ mux_tmp_986));
  assign or_4524_cse = (cfg_proc_precision_rsci_d!=2'b10);
  assign and_2186_cse = or_4524_cse & chn_in_rsci_bawt;
  assign or_3542_cse = (cfg_proc_precision_1_sva_st_102!=2'b10);
  assign and_1091_rgt = ((~ and_tmp_50) | and_1021_cse | (~ main_stage_v_2)) & or_1159_cse
      & or_3538_cse & or_3542_cse & and_dcpl_103;
  assign mux_1050_nl = MUX_s_1_2_2(mux_tmp_1049, (~ or_tmp_1650), cfg_proc_precision_1_sva_st_64[1]);
  assign mux_1051_nl = MUX_s_1_2_2((mux_1050_nl), mux_tmp_1049, cfg_proc_precision_1_sva_st_64[0]);
  assign mux_1052_nl = MUX_s_1_2_2(and_tmp_171, and_2186_cse, or_5189_cse);
  assign mux_1053_cse = MUX_s_1_2_2((mux_1052_nl), (mux_1051_nl), main_stage_v_1);
  assign and_1093_m1c = cvt_4_FpMantRNE_17U_11U_else_and_2_tmp & cvt_unequal_tmp_20
      & or_5189_cse;
  assign or_1659_cse_1 = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_19!=5'b00000);
  assign nl_cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl = (~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_19)
      + 5'b1;
  assign cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl = nl_cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl[4:0];
  assign FpIntToFloat_17U_5U_10U_o_expo_or_12_nl = ((~ cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4)
      & and_1093_m1c) | ((~ cvt_4_FpMantRNE_17U_11U_else_and_2_tmp) & cvt_unequal_tmp_20
      & or_5189_cse);
  assign FpIntToFloat_17U_5U_10U_o_expo_and_25_nl = cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4
      & and_1093_m1c;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_7_itm = MUX1HOT_v_5_3_2((~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_19),
      (cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl), ({1'b0 , FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_9_3_0_1}),
      {(FpIntToFloat_17U_5U_10U_o_expo_or_12_nl) , (FpIntToFloat_17U_5U_10U_o_expo_and_25_nl)
      , (~ mux_1966_itm)});
  assign and_1097_m1c = or_5189_cse & cvt_unequal_tmp_20 & cvt_5_FpMantRNE_17U_11U_else_and_1_tmp;
  assign or_1693_cse = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_20!=5'b00000);
  assign nl_cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl = (~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_20)
      + 5'b1;
  assign cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl = nl_cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl[4:0];
  assign FpIntToFloat_17U_5U_10U_o_expo_or_11_nl = ((~ cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4)
      & and_1097_m1c) | (or_5189_cse & cvt_unequal_tmp_20 & (~ cvt_5_FpMantRNE_17U_11U_else_and_1_tmp));
  assign FpIntToFloat_17U_5U_10U_o_expo_and_23_nl = cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4
      & and_1097_m1c;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_9_itm = MUX1HOT_v_5_3_2((~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_20),
      (cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl), ({1'b0 , FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_9_3_0_1}),
      {(FpIntToFloat_17U_5U_10U_o_expo_or_11_nl) , (FpIntToFloat_17U_5U_10U_o_expo_and_23_nl)
      , (~ mux_1966_itm)});
  assign and_1104_rgt = (or_dcpl_163 | and_1021_cse | (~ main_stage_v_2)) & or_1159_cse
      & or_3538_cse & or_3542_cse & and_dcpl_103;
  assign FpIntToFloat_17U_5U_10U_is_inf_FpIntToFloat_17U_5U_10U_is_inf_or_15_cse
      = (and_tmp_225 & and_dcpl_401) | and_1104_rgt;
  assign nor_1463_nl = ~(main_stage_v_2 | (~ mux_tmp_960));
  assign mux_1071_cse = MUX_s_1_2_2((nor_1463_nl), mux_tmp_961, or_1587_cse);
  assign and_1106_m1c = or_5189_cse & cvt_unequal_tmp_20 & cvt_6_FpMantRNE_17U_11U_else_and_2_tmp;
  assign or_1720_cse_1 = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_21!=5'b00000);
  assign nl_cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl = (~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_21)
      + 5'b1;
  assign cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl = nl_cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl[4:0];
  assign FpIntToFloat_17U_5U_10U_o_expo_or_10_nl = ((~ cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4)
      & and_1106_m1c) | (or_5189_cse & cvt_unequal_tmp_20 & (~ cvt_6_FpMantRNE_17U_11U_else_and_2_tmp));
  assign FpIntToFloat_17U_5U_10U_o_expo_and_21_nl = cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4
      & and_1106_m1c;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_11_itm = MUX1HOT_v_5_3_2((~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_21),
      (cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl), ({1'b0 , FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_9_3_0_1}),
      {(FpIntToFloat_17U_5U_10U_o_expo_or_10_nl) , (FpIntToFloat_17U_5U_10U_o_expo_and_21_nl)
      , (~ mux_1966_itm)});
  assign and_1115_m1c = or_5189_cse & cvt_unequal_tmp_20 & cvt_7_FpMantRNE_17U_11U_else_and_2_tmp;
  assign or_1752_cse_1 = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_22!=5'b00000);
  assign nl_cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl = (~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_22)
      + 5'b1;
  assign cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl = nl_cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl[4:0];
  assign FpIntToFloat_17U_5U_10U_o_expo_or_9_nl = ((~ cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4)
      & and_1115_m1c) | (or_5189_cse & cvt_unequal_tmp_20 & (~ cvt_7_FpMantRNE_17U_11U_else_and_2_tmp));
  assign FpIntToFloat_17U_5U_10U_o_expo_and_19_nl = cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4
      & and_1115_m1c;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_13_itm = MUX1HOT_v_5_3_2((~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_22),
      (cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl), ({1'b0 , FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_9_3_0_1}),
      {(FpIntToFloat_17U_5U_10U_o_expo_or_9_nl) , (FpIntToFloat_17U_5U_10U_o_expo_and_19_nl)
      , (~ mux_1966_itm)});
  assign and_1119_m1c = or_5189_cse & cvt_unequal_tmp_20 & cvt_8_FpMantRNE_17U_11U_else_and_3_tmp;
  assign or_1789_cse_1 = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_23!=5'b00000);
  assign nl_cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl = (~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_23)
      + 5'b1;
  assign cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl = nl_cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl[4:0];
  assign FpIntToFloat_17U_5U_10U_o_expo_or_8_nl = ((~ cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4)
      & and_1119_m1c) | (or_5189_cse & cvt_unequal_tmp_20 & (~ cvt_8_FpMantRNE_17U_11U_else_and_3_tmp));
  assign FpIntToFloat_17U_5U_10U_o_expo_and_17_nl = cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4
      & and_1119_m1c;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_15_itm = MUX1HOT_v_5_3_2((~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_23),
      (cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl), ({1'b0 , FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_9_3_0_1}),
      {(FpIntToFloat_17U_5U_10U_o_expo_or_8_nl) , (FpIntToFloat_17U_5U_10U_o_expo_and_17_nl)
      , (~ mux_1966_itm)});
  assign nor_1434_nl = ~((cfg_proc_precision_1_sva_st_65[1]) | (~ or_4714_cse));
  assign mux_1126_cse = MUX_s_1_2_2((nor_1434_nl), or_4714_cse, cfg_proc_precision_1_sva_st_65[0]);
  assign and_1123_m1c = cvt_9_FpMantRNE_17U_11U_else_and_1_tmp & cvt_unequal_tmp_20
      & or_5189_cse;
  assign or_1829_cse = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_24!=5'b00000);
  assign nl_cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl = (~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_24)
      + 5'b1;
  assign cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl = nl_cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl[4:0];
  assign FpIntToFloat_17U_5U_10U_o_expo_or_7_nl = ((~ cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4)
      & and_1123_m1c) | ((~ cvt_9_FpMantRNE_17U_11U_else_and_1_tmp) & cvt_unequal_tmp_20
      & or_5189_cse);
  assign FpIntToFloat_17U_5U_10U_o_expo_and_15_nl = cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4
      & and_1123_m1c;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_17_itm = MUX1HOT_v_5_3_2((~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_24),
      (cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_3_nl), ({1'b0 , FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_9_3_0_1}),
      {(FpIntToFloat_17U_5U_10U_o_expo_or_7_nl) , (FpIntToFloat_17U_5U_10U_o_expo_and_15_nl)
      , (~ mux_1966_itm)});
  assign FpIntToFloat_17U_5U_10U_is_inf_or_cse = (mux_1142_cse & and_dcpl_401) |
      and_dcpl_617;
  assign and_1132_m1c = or_5189_cse & cvt_unequal_tmp_20 & cvt_10_FpMantRNE_17U_11U_else_and_2_tmp;
  assign or_1851_cse_1 = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_25!=5'b00000);
  assign nl_cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl = (~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_25)
      + 5'b1;
  assign cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl = nl_cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl[4:0];
  assign FpIntToFloat_17U_5U_10U_o_expo_or_6_nl = ((~ cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4)
      & and_1132_m1c) | (or_5189_cse & cvt_unequal_tmp_20 & (~ cvt_10_FpMantRNE_17U_11U_else_and_2_tmp));
  assign FpIntToFloat_17U_5U_10U_o_expo_and_13_nl = cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4
      & and_1132_m1c;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_19_itm = MUX1HOT_v_5_3_2((~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_25),
      (cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl), ({1'b0 , FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_9_3_0_1}),
      {(FpIntToFloat_17U_5U_10U_o_expo_or_6_nl) , (FpIntToFloat_17U_5U_10U_o_expo_and_13_nl)
      , (~ mux_1966_itm)});
  assign nor_1415_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ mux_tmp_455));
  assign mux_1142_cse = MUX_s_1_2_2((nor_1415_nl), mux_tmp_455, cfg_proc_precision_1_sva_st_101[0]);
  assign and_1141_m1c = cvt_11_FpMantRNE_17U_11U_else_and_2_tmp & cvt_unequal_tmp_20
      & or_5189_cse;
  assign or_1892_cse_1 = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_26!=5'b00000);
  assign nl_cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl = (~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_26)
      + 5'b1;
  assign cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl = nl_cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl[4:0];
  assign FpIntToFloat_17U_5U_10U_o_expo_or_5_nl = ((~ cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4)
      & and_1141_m1c) | ((~ cvt_11_FpMantRNE_17U_11U_else_and_2_tmp) & cvt_unequal_tmp_20
      & or_5189_cse);
  assign FpIntToFloat_17U_5U_10U_o_expo_and_11_nl = cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4
      & and_1141_m1c;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_21_itm = MUX1HOT_v_5_3_2((~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_26),
      (cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl), ({1'b0 , FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_9_3_0_1}),
      {(FpIntToFloat_17U_5U_10U_o_expo_or_5_nl) , (FpIntToFloat_17U_5U_10U_o_expo_and_11_nl)
      , (~ mux_1966_itm)});
  assign or_1919_cse = cfg_mode_eql_1_sva_6 | (cfg_out_precision_1_sva_6[0]);
  assign and_1145_m1c = cvt_12_FpMantRNE_17U_11U_else_and_3_tmp & cvt_unequal_tmp_20
      & or_5189_cse;
  assign or_1925_cse_1 = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_27!=5'b00000);
  assign nl_cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl = (~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_27)
      + 5'b1;
  assign cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl = nl_cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl[4:0];
  assign FpIntToFloat_17U_5U_10U_o_expo_or_4_nl = ((~ cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4)
      & and_1145_m1c) | ((~ cvt_12_FpMantRNE_17U_11U_else_and_3_tmp) & cvt_unequal_tmp_20
      & or_5189_cse);
  assign FpIntToFloat_17U_5U_10U_o_expo_and_9_nl = cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4
      & and_1145_m1c;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_23_itm = MUX1HOT_v_5_3_2((~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_27),
      (cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl), ({1'b0 , FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_9_3_0_1}),
      {(FpIntToFloat_17U_5U_10U_o_expo_or_4_nl) , (FpIntToFloat_17U_5U_10U_o_expo_and_9_nl)
      , (~ mux_1966_itm)});
  assign and_283_cse = main_stage_v_3 & mux_tmp_987;
  assign FpIntToFloat_17U_5U_10U_is_inf_and_8_cse = core_wen & ((and_dcpl_499 & and_dcpl_626)
      | and_dcpl_631);
  assign and_1155_m1c = cvt_13_FpMantRNE_17U_11U_else_and_2_tmp & cvt_unequal_tmp_20
      & or_5189_cse;
  assign nl_cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl = (~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_28)
      + 5'b1;
  assign cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl = nl_cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl[4:0];
  assign FpIntToFloat_17U_5U_10U_o_expo_or_3_nl = ((~ cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4)
      & and_1155_m1c) | ((~ cvt_13_FpMantRNE_17U_11U_else_and_2_tmp) & cvt_unequal_tmp_20
      & or_5189_cse);
  assign FpIntToFloat_17U_5U_10U_o_expo_and_7_nl = cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4
      & and_1155_m1c;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_25_itm = MUX1HOT_v_5_3_2((~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_28),
      (cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_5_nl), ({1'b0 , FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_9_3_0_1}),
      {(FpIntToFloat_17U_5U_10U_o_expo_or_3_nl) , (FpIntToFloat_17U_5U_10U_o_expo_and_7_nl)
      , (~ mux_1966_itm)});
  assign or_5038_cse = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_28!=5'b00000);
  assign and_1159_m1c = or_5189_cse & cvt_unequal_tmp_20 & cvt_14_FpMantRNE_17U_11U_else_and_3_tmp;
  assign nl_cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl = (~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_29)
      + 5'b1;
  assign cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl = nl_cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl[4:0];
  assign FpIntToFloat_17U_5U_10U_o_expo_or_2_nl = ((~ cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4)
      & and_1159_m1c) | (or_5189_cse & cvt_unequal_tmp_20 & (~ cvt_14_FpMantRNE_17U_11U_else_and_3_tmp));
  assign FpIntToFloat_17U_5U_10U_o_expo_and_5_nl = cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4
      & and_1159_m1c;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_27_itm = MUX1HOT_v_5_3_2((~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_29),
      (cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl), ({1'b0 , FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_9_3_0_1}),
      {(FpIntToFloat_17U_5U_10U_o_expo_or_2_nl) , (FpIntToFloat_17U_5U_10U_o_expo_and_5_nl)
      , (~ mux_1966_itm)});
  assign or_5053_cse = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_29!=5'b00000);
  assign mux_2000_nl = MUX_s_1_2_2((cfg_out_precision_1_sva_6[1]), (cfg_out_precision_1_sva_st_149[1]),
      or_5189_cse);
  assign IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_mux_rgt = MUX_v_15_2_2(IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_2,
      ({5'b0 , FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_40_itm_mx0w0}),
      mux_2000_nl);
  assign FpIntToFloat_17U_5U_10U_is_inf_and_10_cse = core_wen & ((and_dcpl_473 &
      and_dcpl_626) | and_dcpl_648);
  assign and_1172_m1c = or_5189_cse & cvt_unequal_tmp_20 & cvt_15_FpMantRNE_17U_11U_else_and_3_tmp;
  assign nl_cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl = (~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_30)
      + 5'b1;
  assign cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl = nl_cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl[4:0];
  assign FpIntToFloat_17U_5U_10U_o_expo_or_1_nl = ((~ cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4)
      & and_1172_m1c) | (or_5189_cse & cvt_unequal_tmp_20 & (~ cvt_15_FpMantRNE_17U_11U_else_and_3_tmp));
  assign FpIntToFloat_17U_5U_10U_o_expo_and_3_nl = cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4
      & and_1172_m1c;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_29_itm = MUX1HOT_v_5_3_2((~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_30),
      (cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_7_nl), ({1'b0 , FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_9_3_0_1}),
      {(FpIntToFloat_17U_5U_10U_o_expo_or_1_nl) , (FpIntToFloat_17U_5U_10U_o_expo_and_3_nl)
      , (~ mux_1966_itm)});
  assign or_5069_cse = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_30!=5'b00000);
  assign and_1176_m1c = cvt_16_FpMantRNE_17U_11U_else_and_4_tmp & cvt_unequal_tmp_20
      & or_5189_cse;
  assign nl_cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_9_nl = (~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_31)
      + 5'b1;
  assign cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_9_nl = nl_cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_9_nl[4:0];
  assign FpIntToFloat_17U_5U_10U_o_expo_or_nl = ((~ cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_8_tmp_4)
      & and_1176_m1c) | ((~ cvt_16_FpMantRNE_17U_11U_else_and_4_tmp) & cvt_unequal_tmp_20
      & or_5189_cse);
  assign FpIntToFloat_17U_5U_10U_o_expo_and_1_nl = cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_8_tmp_4
      & and_1176_m1c;
  assign FpIntToFloat_17U_5U_10U_o_expo_mux1h_31_itm = MUX1HOT_v_5_3_2((~ libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_31),
      (cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_9_nl), ({1'b0 , FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_9_3_0_1}),
      {(FpIntToFloat_17U_5U_10U_o_expo_or_nl) , (FpIntToFloat_17U_5U_10U_o_expo_and_1_nl)
      , (~ mux_1966_itm)});
  assign or_5086_cse = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_31!=5'b00000);
  assign and_271_nl = main_stage_v_3 & mux_tmp_986;
  assign mux_1267_nl = MUX_s_1_2_2((and_271_nl), and_tmp_94, or_5189_cse);
  assign cfg_proc_precision_and_40_cse = core_wen & (~ and_dcpl_93) & (mux_1267_nl);
  assign and_295_nl = main_stage_v_3 & or_1159_cse;
  assign mux_1268_nl = MUX_s_1_2_2((and_295_nl), and_2237_cse, or_5189_cse);
  assign cfg_proc_precision_and_43_cse = core_wen & (~ and_dcpl_93) & (mux_1268_nl);
  assign FpFloatToInt_16U_5U_10U_and_nl = (~ (chn_idata_data_sva_2_47_31_1[0])) &
      FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_m1c & and_dcpl_408;
  assign FpFloatToInt_16U_5U_10U_and_32_nl = (chn_idata_data_sva_2_47_31_1[0]) &
      FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_m1c & and_dcpl_408;
  assign FpFloatToInt_16U_5U_10U_and_1_nl = cvt_1_FpFloatToInt_16U_5U_10U_if_acc_itm_11_1
      & (~ IsNaN_5U_10U_land_1_lpi_1_dfm_mx0w0) & and_dcpl_408;
  assign FpFloatToInt_16U_5U_10U_o_int_and_15_nl = IsNaN_5U_10U_land_1_lpi_1_dfm_mx0w0
      & and_dcpl_408;
  assign and_908_nl = or_4862_cse & (~ (cfg_out_precision_1_sva_st_113[0])) & and_dcpl_420;
  assign FpFloatToInt_16U_5U_10U_o_int_mux1h_nl = MUX1HOT_v_15_6_2((FpFloatToInt_16U_5U_10U_internal_int_24_1_1_sva[14:0]),
      (FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_1_sva[15:1]), (FpFloatToInt_16U_5U_10U_if_qr_1_lpi_1_dfm_mx0[15:1]),
      15'b100000000000000, IntSaturation_17U_16U_o_15_1_1_lpi_1_dfm_5, IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_2,
      {(FpFloatToInt_16U_5U_10U_and_nl) , (FpFloatToInt_16U_5U_10U_and_32_nl) , (FpFloatToInt_16U_5U_10U_and_1_nl)
      , (FpFloatToInt_16U_5U_10U_o_int_and_15_nl) , and_dcpl_425 , (and_908_nl)});
  assign nl_cvt_1_FpMantRNE_17U_11U_else_acc_nl = (FpIntToFloat_17U_5U_10U_else_int_mant_1_sva[15:6])
      + conv_u2u_1_10(FpMantRNE_17U_11U_else_carry_1_sva);
  assign cvt_1_FpMantRNE_17U_11U_else_acc_nl = nl_cvt_1_FpMantRNE_17U_11U_else_acc_nl[9:0];
  assign FpIntToFloat_17U_5U_10U_if_not_176_nl = ~ IsNaN_5U_10U_IsNaN_5U_10U_nand_1_itm_2;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_1_nl = MUX_v_10_2_2(10'b0000000000,
      (cvt_1_FpMantRNE_17U_11U_else_acc_nl), (FpIntToFloat_17U_5U_10U_if_not_176_nl));
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_14_nl = MUX_v_10_2_2((FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_1_nl),
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_1_lpi_1_dfm_8, and_dcpl_408);
  assign and_1179_nl = or_5189_cse & cfg_mode_eql_1_sva_5;
  assign mux_2010_nl = MUX_s_1_2_2((cfg_out_precision_1_sva_st_113[1]), or_300_cse,
      cfg_proc_precision_1_sva_st_65[1]);
  assign mux_2011_nl = MUX_s_1_2_2((mux_2010_nl), (cfg_out_precision_1_sva_st_113[1]),
      cfg_proc_precision_1_sva_st_65[0]);
  assign or_3597_nl = cfg_mode_eql_1_sva_5 | (mux_2011_nl);
  assign mux_2012_nl = MUX_s_1_2_2(or_1176_cse, cfg_mode_eql_1_sva_6, cvt_unequal_tmp_21);
  assign or_3600_nl = (cfg_out_precision_1_sva_6[1]) | cfg_mode_eql_1_sva_6;
  assign mux_2013_nl = MUX_s_1_2_2(cfg_mode_eql_1_sva_6, (or_3600_nl), cvt_unequal_tmp_21);
  assign mux_2014_nl = MUX_s_1_2_2((mux_2013_nl), (mux_2012_nl), nor_1672_cse);
  assign mux_2015_nl = MUX_s_1_2_2((mux_2014_nl), (or_3597_nl), or_5189_cse);
  assign mux_2017_nl = MUX_s_1_2_2(or_1198_cse, or_4709_cse, nor_50_cse);
  assign or_3606_nl = cfg_mode_eql_1_sva_5 | (mux_2017_nl);
  assign or_3607_nl = nor_1672_cse | (cfg_out_precision_1_sva_6!=2'b10) | cfg_mode_eql_1_sva_6;
  assign or_3609_nl = nor_1629_cse | cfg_mode_eql_1_sva_6;
  assign mux_2018_nl = MUX_s_1_2_2(cfg_mode_eql_1_sva_6, (or_3609_nl), nor_1672_cse);
  assign mux_2019_nl = MUX_s_1_2_2((mux_2018_nl), (or_3607_nl), cvt_unequal_tmp_21);
  assign mux_2020_nl = MUX_s_1_2_2((mux_2019_nl), (or_3606_nl), or_5189_cse);
  assign chn_idata_data_mux1h_65_rgt = MUX1HOT_v_16_3_2(chn_idata_data_sva_2_15_0_1,
      ({1'b0 , (FpFloatToInt_16U_5U_10U_o_int_mux1h_nl)}), ({6'b0 , (FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_mux_14_nl)}),
      {(and_1179_nl) , (~ (mux_2015_nl)) , (~ (mux_2020_nl))});
  assign or_3817_cse = (~ mux_tmp_455) | and_1021_cse;
  assign or_3774_cse = or_dcpl_163 | and_1021_cse;
  assign or_3623_cse = nor_8_cse | (cfg_out_precision_1_sva_st_154[0]);
  assign FpIntToFloat_17U_5U_10U_is_inf_FpIntToFloat_17U_5U_10U_is_inf_or_10_cse
      = (or_3696_cse & or_4862_cse & or_4714_cse & or_400_cse_1 & or_5189_cse & main_stage_v_2
      & (cfg_out_precision_1_sva_st_149==2'b10)) | and_1249_cse;
  assign mux_1342_nl = MUX_s_1_2_2(mux_tmp_1341, (~ mux_tmp_1332), reg_cfg_proc_precision_1_sva_st_40_cse[1]);
  assign mux_1343_nl = MUX_s_1_2_2((mux_1342_nl), mux_tmp_1341, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign mux_1344_nl = MUX_s_1_2_2(mux_tmp_1332, (~ (mux_1343_nl)), cfg_out_precision_1_sva_st_154[1]);
  assign mux_1345_nl = MUX_s_1_2_2((mux_1344_nl), mux_tmp_1332, or_3623_cse);
  assign FpIntToFloat_17U_5U_10U_is_inf_and_23_cse = core_wen & FpIntToFloat_17U_5U_10U_is_inf_FpIntToFloat_17U_5U_10U_is_inf_or_10_cse
      & (~ (mux_1345_nl));
  assign and_1213_rgt = and_tmp_12 & and_dcpl_363 & or_5189_cse;
  assign nand_190_cse = ~((cfg_out_precision_1_sva_st_149[1]) & main_stage_v_2);
  assign nor_1314_nl = ~(nor_50_cse | nor_2219_cse | nor_151_cse | (cfg_out_precision_1_sva_st_149[0])
      | nand_190_cse);
  assign mux_1436_cse = MUX_s_1_2_2(main_stage_v_2, (nor_1314_nl), or_1587_cse);
  assign mux_1437_cse = MUX_s_1_2_2(mux_1436_cse, main_stage_v_1, or_5189_cse);
  assign mux_1438_nl = MUX_s_1_2_2(mux_tmp_1435, (~ mux_1437_cse), cfg_out_precision_1_sva_st_154[1]);
  assign mux_1439_nl = MUX_s_1_2_2((mux_1438_nl), mux_tmp_1435, or_4559_cse);
  assign mux_1441_nl = MUX_s_1_2_2((mux_1439_nl), mux_tmp_1435, nor_2150_cse);
  assign mux_1442_nl = MUX_s_1_2_2((mux_1441_nl), mux_tmp_1435, nor_8_cse);
  assign FpIntToFloat_17U_5U_10U_is_inf_and_26_cse = core_wen & FpIntToFloat_17U_5U_10U_is_inf_FpIntToFloat_17U_5U_10U_is_inf_or_10_cse
      & (~ (mux_1442_nl));
  assign nor_1309_cse = ~((~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | (~ cvt_unequal_tmp_19) | cfg_mode_eql_1_sva_4);
  assign nor_1310_cse = ~((~ cvt_unequal_tmp_20) | (cfg_out_precision_1_sva_st_113!=2'b10)
      | cfg_mode_eql_1_sva_5 | (~ main_stage_v_2));
  assign mux_1458_nl = MUX_s_1_2_2(nor_1310_cse, nor_1309_cse, or_5189_cse);
  assign FpIntToFloat_17U_5U_10U_if_and_16_cse = core_wen & (~ and_dcpl_93) & (mux_1458_nl);
  assign or_2289_cse = (~ cvt_unequal_tmp_19) | cfg_mode_eql_1_sva_4 | (cfg_out_precision_1_sva_st_154!=2'b10);
  assign nor_1306_nl = ~((cfg_proc_precision_1_sva_st_89[1]) | (~ mux_tmp_658));
  assign mux_1463_cse = MUX_s_1_2_2((nor_1306_nl), mux_tmp_658, cfg_proc_precision_1_sva_st_89[0]);
  assign nor_2130_nl = ~(nor_50_cse | (cfg_out_precision_1_sva_st_149[0]) | (~((cfg_out_precision_1_sva_st_149[1])
      & mux_1463_cse)));
  assign mux_1464_cse = MUX_s_1_2_2(main_stage_v_2, (nor_2130_nl), or_1587_cse);
  assign and_1247_rgt = or_3696_cse & or_5189_cse;
  assign nor_1305_nl = ~((reg_cfg_proc_precision_1_sva_st_40_cse[1]) | (~ mux_1466_cse));
  assign mux_1460_cse = MUX_s_1_2_2((nor_1305_nl), mux_1466_cse, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign FpIntToFloat_17U_5U_10U_if_FpIntToFloat_17U_5U_10U_if_or_11_cse = and_1249_cse
      | and_1247_rgt;
  assign nor_2114_nl = ~(nor_8_cse | (cfg_out_precision_1_sva_st_154[0]) | (~((cfg_out_precision_1_sva_st_154[1])
      & mux_1460_cse)));
  assign mux_1461_nl = MUX_s_1_2_2(main_stage_v_1, (nor_2114_nl), or_2289_cse);
  assign mux_1465_nl = MUX_s_1_2_2(mux_1464_cse, (mux_1461_nl), or_5189_cse);
  assign FpIntToFloat_17U_5U_10U_if_and_18_cse = core_wen & FpIntToFloat_17U_5U_10U_if_FpIntToFloat_17U_5U_10U_if_or_11_cse
      & (mux_1465_nl);
  assign and_1250_rgt = or_tmp_2960 & or_5189_cse;
  assign nor_1301_nl = ~((reg_cfg_proc_precision_1_sva_st_40_cse[1]) | (~ main_stage_v_1));
  assign mux_1466_cse = MUX_s_1_2_2((nor_1301_nl), main_stage_v_1, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign and_1249_cse = and_tmp_12 & and_dcpl_228 & or_5189_cse;
  assign nor_2127_nl = ~(nor_50_cse | (cfg_out_precision_1_sva_st_149[0]) | (~((cfg_out_precision_1_sva_st_149[1])
      & mux_786_cse_1)));
  assign mux_1494_cse = MUX_s_1_2_2(main_stage_v_2, (nor_2127_nl), or_1587_cse);
  assign nor_1287_nl = ~((reg_cfg_proc_precision_1_sva_st_40_cse[1]) | (~ mux_1460_cse));
  assign mux_1489_cse = MUX_s_1_2_2((nor_1287_nl), mux_1460_cse, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign nor_2110_nl = ~(nor_8_cse | (cfg_out_precision_1_sva_st_154[0]) | (~((cfg_out_precision_1_sva_st_154[1])
      & mux_1489_cse)));
  assign mux_1490_nl = MUX_s_1_2_2(main_stage_v_1, (nor_2110_nl), or_2289_cse);
  assign mux_1495_nl = MUX_s_1_2_2(mux_1494_cse, (mux_1490_nl), or_5189_cse);
  assign FpIntToFloat_17U_5U_10U_if_and_22_cse = core_wen & FpIntToFloat_17U_5U_10U_if_FpIntToFloat_17U_5U_10U_if_or_11_cse
      & (mux_1495_nl);
  assign nand_171_cse = ~((cfg_out_precision_1_sva_st_154[1]) & main_stage_v_1);
  assign nor_1271_nl = ~(nor_8_cse | nor_2150_cse | (cfg_out_precision_1_sva_st_154[0])
      | nand_171_cse);
  assign mux_1519_nl = MUX_s_1_2_2(main_stage_v_1, (nor_1271_nl), or_2289_cse);
  assign mux_1521_cse = MUX_s_1_2_2(mux_1436_cse, (mux_1519_nl), or_5189_cse);
  assign FpIntToFloat_17U_5U_10U_if_and_27_cse = core_wen & FpIntToFloat_17U_5U_10U_if_FpIntToFloat_17U_5U_10U_if_or_11_cse
      & mux_1521_cse;
  assign or_3696_cse = or_dcpl_15 | (cfg_out_precision_1_sva_st_154!=2'b10);
  assign mux_124_nl = MUX_s_1_2_2(and_tmp_19, and_2186_cse, or_5189_cse);
  assign IntShiftRightSat_49U_6U_17U_o_and_107_cse = cvt_else_and_cse & (~ or_dcpl_16)
      & (~ (mux_124_nl));
  assign mux_130_nl = MUX_s_1_2_2(mux_tmp_129, and_2186_cse, or_5189_cse);
  assign IntShiftRightSat_49U_6U_17U_o_and_108_cse = cvt_else_and_cse & (~ or_dcpl_32)
      & (~ (mux_130_nl));
  assign mux_133_cse = MUX_s_1_2_2(and_1386_cse, and_2186_cse, or_5189_cse);
  assign IntShiftRightSat_49U_6U_17U_o_and_109_cse = cvt_else_and_cse & (~ or_dcpl_16)
      & (~ mux_133_cse);
  assign IntShiftRightSat_49U_6U_17U_o_and_111_cse = cvt_else_and_cse & (~ or_dcpl_32)
      & (~ mux_133_cse);
  assign mux_118_nl = MUX_s_1_2_2(and_tmp_16, and_2186_cse, or_5189_cse);
  assign IntShiftRightSat_49U_6U_17U_o_and_112_cse = cvt_else_and_cse & (~ or_dcpl_16)
      & (~ (mux_118_nl));
  assign mux_149_nl = MUX_s_1_2_2(and_tmp_33, and_2186_cse, or_5189_cse);
  assign IntShiftRightSat_49U_6U_17U_o_and_114_cse = cvt_else_and_cse & (~ or_dcpl_32)
      & (~ (mux_149_nl));
  assign mux_152_nl = MUX_s_1_2_2(mux_tmp_151, and_2186_cse, or_5189_cse);
  assign IntShiftRightSat_49U_6U_17U_o_and_115_cse = cvt_else_and_cse & (~ or_dcpl_32)
      & (~ (mux_152_nl));
  assign nand_164_cse = ~(cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_nand_itm_2);
  assign nand_162_cse = ~(cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_nand_1_itm_2);
  assign nand_160_cse = ~(cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_nand_2_itm_2);
  assign nand_158_cse = ~(cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_nand_3_itm_2);
  assign nand_156_cse = ~(cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_nand_4_itm_2);
  assign nand_153_cse = ~(cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_nand_5_itm_2);
  assign nand_151_cse = ~(cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_nand_6_itm_2);
  assign nand_149_cse = ~(cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_nand_7_itm_2);
  assign nand_147_cse = ~(cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_nand_8_itm_2);
  assign nand_145_cse = ~(cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_nand_9_itm_2);
  assign nand_143_cse = ~(cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_nand_10_itm_2);
  assign nand_141_cse = ~(cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_nand_11_itm_2);
  assign nand_139_cse = ~(cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_nand_12_itm_2);
  assign nand_137_cse = ~(cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_nand_13_itm_2);
  assign nand_135_cse = ~(cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_nand_14_itm_2);
  assign nand_133_cse = ~(cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_4_svs_st_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_nand_15_itm_2);
  assign and_1321_rgt = or_dcpl_320 & or_5189_cse;
  assign and_1325_rgt = or_dcpl_322 & or_5189_cse;
  assign and_1329_rgt = or_dcpl_324 & or_5189_cse;
  assign and_1333_rgt = or_dcpl_326 & or_5189_cse;
  assign and_1337_rgt = or_dcpl_328 & or_5189_cse;
  assign and_1341_rgt = or_dcpl_330 & or_5189_cse;
  assign and_1345_rgt = or_dcpl_332 & or_5189_cse;
  assign and_1349_rgt = or_dcpl_334 & or_5189_cse;
  assign and_1353_rgt = or_dcpl_336 & or_5189_cse;
  assign and_1357_rgt = or_dcpl_338 & or_5189_cse;
  assign and_1361_rgt = or_dcpl_340 & or_5189_cse;
  assign and_1365_rgt = or_dcpl_342 & or_5189_cse;
  assign and_1369_rgt = or_dcpl_344 & or_5189_cse;
  assign and_1373_rgt = or_dcpl_346 & or_5189_cse;
  assign and_1377_rgt = or_dcpl_348 & or_5189_cse;
  assign and_1381_rgt = or_dcpl_350 & or_5189_cse;
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_rgt = ~(cvt_16_IntSaturation_17U_16U_else_if_acc_4_itm_2_1
      | cvt_16_IntSaturation_17U_16U_if_acc_4_itm_2_1 | and_dcpl_93);
  assign IntSaturation_17U_16U_and_31_rgt = cvt_16_IntSaturation_17U_16U_else_if_acc_4_itm_2_1
      & (~ cvt_16_IntSaturation_17U_16U_if_acc_4_itm_2_1) & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_and_31_rgt = cvt_16_IntSaturation_17U_16U_if_acc_4_itm_2_1
      & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_1_rgt = ~(cvt_15_IntSaturation_17U_16U_else_if_acc_3_itm_2_1
      | cvt_15_IntSaturation_17U_16U_if_acc_3_itm_2_1 | and_dcpl_93);
  assign IntSaturation_17U_16U_and_29_rgt = cvt_15_IntSaturation_17U_16U_else_if_acc_3_itm_2_1
      & (~ cvt_15_IntSaturation_17U_16U_if_acc_3_itm_2_1) & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_and_29_rgt = cvt_15_IntSaturation_17U_16U_if_acc_3_itm_2_1
      & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_2_rgt = ~(cvt_14_IntSaturation_17U_16U_else_if_acc_3_itm_2_1
      | cvt_14_IntSaturation_17U_16U_if_acc_3_itm_2_1 | and_dcpl_93);
  assign IntSaturation_17U_16U_and_27_rgt = cvt_14_IntSaturation_17U_16U_else_if_acc_3_itm_2_1
      & (~ cvt_14_IntSaturation_17U_16U_if_acc_3_itm_2_1) & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_and_27_rgt = cvt_14_IntSaturation_17U_16U_if_acc_3_itm_2_1
      & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_3_rgt = ~(cvt_13_IntSaturation_17U_16U_else_if_acc_2_itm_2_1
      | cvt_13_IntSaturation_17U_16U_if_acc_2_itm_2_1 | and_dcpl_93);
  assign IntSaturation_17U_16U_and_25_rgt = cvt_13_IntSaturation_17U_16U_else_if_acc_2_itm_2_1
      & (~ cvt_13_IntSaturation_17U_16U_if_acc_2_itm_2_1) & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_and_25_rgt = cvt_13_IntSaturation_17U_16U_if_acc_2_itm_2_1
      & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_4_rgt = ~(cvt_12_IntSaturation_17U_16U_else_if_acc_3_itm_2_1
      | cvt_12_IntSaturation_17U_16U_if_acc_3_itm_2_1 | and_dcpl_93);
  assign IntSaturation_17U_16U_and_23_rgt = cvt_12_IntSaturation_17U_16U_else_if_acc_3_itm_2_1
      & (~ cvt_12_IntSaturation_17U_16U_if_acc_3_itm_2_1) & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_and_23_rgt = cvt_12_IntSaturation_17U_16U_if_acc_3_itm_2_1
      & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_5_rgt = ~(cvt_11_IntSaturation_17U_16U_else_if_acc_2_itm_2_1
      | cvt_11_IntSaturation_17U_16U_if_acc_2_itm_2_1 | and_dcpl_93);
  assign IntSaturation_17U_16U_and_21_rgt = cvt_11_IntSaturation_17U_16U_else_if_acc_2_itm_2_1
      & (~ cvt_11_IntSaturation_17U_16U_if_acc_2_itm_2_1) & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_and_21_rgt = cvt_11_IntSaturation_17U_16U_if_acc_2_itm_2_1
      & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_6_rgt = ~(cvt_10_IntSaturation_17U_16U_else_if_acc_2_itm_2_1
      | cvt_10_IntSaturation_17U_16U_if_acc_2_itm_2_1 | and_dcpl_93);
  assign IntSaturation_17U_16U_and_19_rgt = cvt_10_IntSaturation_17U_16U_else_if_acc_2_itm_2_1
      & (~ cvt_10_IntSaturation_17U_16U_if_acc_2_itm_2_1) & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_and_19_rgt = cvt_10_IntSaturation_17U_16U_if_acc_2_itm_2_1
      & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_7_rgt = ~(cvt_9_IntSaturation_17U_16U_else_if_acc_1_itm_2_1
      | cvt_9_IntSaturation_17U_16U_if_acc_1_itm_2_1 | and_dcpl_93);
  assign IntSaturation_17U_16U_and_17_rgt = cvt_9_IntSaturation_17U_16U_else_if_acc_1_itm_2_1
      & (~ cvt_9_IntSaturation_17U_16U_if_acc_1_itm_2_1) & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_and_17_rgt = cvt_9_IntSaturation_17U_16U_if_acc_1_itm_2_1
      & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_8_rgt = ~(cvt_8_IntSaturation_17U_16U_else_if_acc_3_itm_2_1
      | cvt_8_IntSaturation_17U_16U_if_acc_3_itm_2_1 | and_dcpl_93);
  assign IntSaturation_17U_16U_and_15_rgt = cvt_8_IntSaturation_17U_16U_else_if_acc_3_itm_2_1
      & (~ cvt_8_IntSaturation_17U_16U_if_acc_3_itm_2_1) & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_and_15_rgt = cvt_8_IntSaturation_17U_16U_if_acc_3_itm_2_1
      & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_9_rgt = ~(cvt_7_IntSaturation_17U_16U_else_if_acc_2_itm_2_1
      | cvt_7_IntSaturation_17U_16U_if_acc_2_itm_2_1 | and_dcpl_93);
  assign IntSaturation_17U_16U_and_13_rgt = cvt_7_IntSaturation_17U_16U_else_if_acc_2_itm_2_1
      & (~ cvt_7_IntSaturation_17U_16U_if_acc_2_itm_2_1) & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_and_13_rgt = cvt_7_IntSaturation_17U_16U_if_acc_2_itm_2_1
      & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_10_rgt = ~(cvt_6_IntSaturation_17U_16U_else_if_acc_2_itm_2_1
      | cvt_6_IntSaturation_17U_16U_if_acc_2_itm_2_1 | and_dcpl_93);
  assign IntSaturation_17U_16U_and_11_rgt = cvt_6_IntSaturation_17U_16U_else_if_acc_2_itm_2_1
      & (~ cvt_6_IntSaturation_17U_16U_if_acc_2_itm_2_1) & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_and_11_rgt = cvt_6_IntSaturation_17U_16U_if_acc_2_itm_2_1
      & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_11_rgt = ~(cvt_5_IntSaturation_17U_16U_else_if_acc_1_itm_2_1
      | cvt_5_IntSaturation_17U_16U_if_acc_1_itm_2_1 | and_dcpl_93);
  assign IntSaturation_17U_16U_and_9_rgt = cvt_5_IntSaturation_17U_16U_else_if_acc_1_itm_2_1
      & (~ cvt_5_IntSaturation_17U_16U_if_acc_1_itm_2_1) & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_and_9_rgt = cvt_5_IntSaturation_17U_16U_if_acc_1_itm_2_1
      & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_12_rgt = ~(cvt_4_IntSaturation_17U_16U_else_if_acc_2_itm_2_1
      | cvt_4_IntSaturation_17U_16U_if_acc_2_itm_2_1 | and_dcpl_93);
  assign IntSaturation_17U_16U_and_7_rgt = cvt_4_IntSaturation_17U_16U_else_if_acc_2_itm_2_1
      & (~ cvt_4_IntSaturation_17U_16U_if_acc_2_itm_2_1) & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_and_7_rgt = cvt_4_IntSaturation_17U_16U_if_acc_2_itm_2_1
      & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_13_rgt = ~(cvt_3_IntSaturation_17U_16U_else_if_acc_1_itm_2_1
      | cvt_3_IntSaturation_17U_16U_if_acc_1_itm_2_1 | and_dcpl_93);
  assign IntSaturation_17U_16U_and_5_rgt = cvt_3_IntSaturation_17U_16U_else_if_acc_1_itm_2_1
      & (~ cvt_3_IntSaturation_17U_16U_if_acc_1_itm_2_1) & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_and_5_rgt = cvt_3_IntSaturation_17U_16U_if_acc_1_itm_2_1
      & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_14_rgt = ~(cvt_2_IntSaturation_17U_16U_else_if_acc_1_itm_2_1
      | cvt_2_IntSaturation_17U_16U_if_acc_1_itm_2_1 | and_dcpl_93);
  assign IntSaturation_17U_16U_and_3_rgt = cvt_2_IntSaturation_17U_16U_else_if_acc_1_itm_2_1
      & (~ cvt_2_IntSaturation_17U_16U_if_acc_1_itm_2_1) & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_and_3_rgt = cvt_2_IntSaturation_17U_16U_if_acc_1_itm_2_1
      & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_15_rgt = ~(cvt_1_IntSaturation_17U_16U_else_if_acc_itm_2_1
      | cvt_1_IntSaturation_17U_16U_if_acc_itm_2_1 | and_dcpl_93);
  assign IntSaturation_17U_16U_and_1_rgt = cvt_1_IntSaturation_17U_16U_else_if_acc_itm_2_1
      & (~ cvt_1_IntSaturation_17U_16U_if_acc_itm_2_1) & (~ and_dcpl_93);
  assign IntSaturation_17U_16U_o_and_1_rgt = cvt_1_IntSaturation_17U_16U_if_acc_itm_2_1
      & (~ and_dcpl_93);
  assign nor_1195_nl = ~((~ main_stage_v_1) | (~ cvt_unequal_tmp_19) | cfg_mode_eql_1_sva_4);
  assign mux_1626_nl = MUX_s_1_2_2(nor_1556_cse, (nor_1195_nl), or_5189_cse);
  assign IntSaturation_17U_16U_and_33_cse = core_wen & (~ and_dcpl_93) & (mux_1626_nl);
  assign nor_1185_cse = ~((cfg_out_precision_1_sva_st_154!=2'b01) | (~ main_stage_v_1));
  assign nor_1186_cse = ~((cfg_out_precision_1_sva_st_149!=2'b01) | (~ main_stage_v_2));
  assign mux_1653_nl = MUX_s_1_2_2(mux_1489_cse, nor_1185_cse, cfg_proc_precision_1_sva_st_64[1]);
  assign mux_1654_cse = MUX_s_1_2_2((mux_1653_nl), mux_1489_cse, cfg_proc_precision_1_sva_st_64[0]);
  assign and_1386_cse = main_stage_v_1 & and_tmp_12;
  assign and_1385_rgt = and_tmp_12 & and_dcpl_114;
  assign IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_19_cse
      = (or_dcpl_16 & or_4862_cse & or_4714_cse & and_dcpl_401) | and_1385_rgt;
  assign or_479_nl = main_stage_v_2 | (~ and_1386_cse);
  assign mux_272_cse = MUX_s_1_2_2((or_479_nl), or_5379_cse, or_5189_cse);
  assign IntShiftRightSat_49U_6U_17U_oelse_and_cse = cvt_else_and_cse & IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_19_cse
      & mux_272_cse;
  assign or_547_nl = main_stage_v_2 | (~ and_tmp_16);
  assign mux_320_cse = MUX_s_1_2_2((or_547_nl), or_5379_cse, or_5189_cse);
  assign IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_18_cse
      = (or_dcpl_16 & or_4862_cse & or_4714_cse & or_400_cse_1 & and_dcpl_401) |
      and_1385_rgt;
  assign or_626_nl = main_stage_v_2 | (~ and_tmp_19);
  assign mux_377_nl = MUX_s_1_2_2((or_626_nl), or_5379_cse, or_5189_cse);
  assign IntShiftRightSat_49U_6U_17U_oelse_and_18_cse = cvt_else_and_cse & IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_18_cse
      & (mux_377_nl);
  assign IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_15_cse
      = (or_dcpl_32 & or_4862_cse & or_4714_cse & or_400_cse_1 & and_dcpl_401) |
      and_1385_rgt;
  assign IntShiftRightSat_49U_6U_17U_oelse_and_22_cse = cvt_else_and_cse & IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_18_cse
      & mux_272_cse;
  assign IntShiftRightSat_49U_6U_17U_oelse_and_25_cse = cvt_else_and_cse & ((or_dcpl_16
      & or_4862_cse & or_4714_cse & or_5189_cse & and_dcpl_626) | and_1385_rgt) &
      mux_320_cse;
  assign IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_8_cse
      = (or_dcpl_32 & or_4862_cse & or_4714_cse & or_5189_cse & and_dcpl_626) | and_1385_rgt;
  assign or_5379_cse = (~ and_2186_cse) | main_stage_v_1;
  assign and_1467_rgt = and_tmp_11 & or_5189_cse;
  assign or_186_cse = (reg_cfg_proc_precision_1_sva_st_40_cse!=2'b10) | and_dcpl_3;
  assign and_1021_cse = (cfg_proc_precision_1_sva_st_101==2'b10);
  assign mux_1283_nl = MUX_s_1_2_2(mux_tmp_1282, (~ mux_tmp_1276), reg_cfg_proc_precision_1_sva_st_40_cse[1]);
  assign mux_1284_nl = MUX_s_1_2_2((mux_1283_nl), mux_tmp_1282, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign mux_1285_nl = MUX_s_1_2_2(mux_tmp_1276, (~ (mux_1284_nl)), cfg_out_precision_1_sva_st_154[1]);
  assign mux_1286_nl = MUX_s_1_2_2((mux_1285_nl), mux_tmp_1276, or_3623_cse);
  assign FpIntToFloat_17U_5U_10U_is_inf_and_28_cse = core_wen & FpIntToFloat_17U_5U_10U_is_inf_FpIntToFloat_17U_5U_10U_is_inf_or_10_cse
      & (~ (mux_1286_nl));
  assign FpIntToFloat_17U_5U_10U_if_nor_10_cse = ~(or_dcpl_15 | (~ main_stage_v_1)
      | (cfg_out_precision_1_sva_st_154!=2'b10));
  assign or_217_nl = (cfg_out_precision_1_sva_st_154!=2'b10) | (~ and_tmp_16);
  assign mux_119_nl = MUX_s_1_2_2((or_217_nl), or_tmp_213, or_5189_cse);
  assign FpIntToFloat_17U_5U_10U_if_and_31_cse = cvt_else_and_cse & FpIntToFloat_17U_5U_10U_if_nor_10_cse
      & (mux_119_nl);
  assign or_226_nl = (cfg_out_precision_1_sva_st_154!=2'b10) | (~ and_tmp_19);
  assign mux_125_nl = MUX_s_1_2_2((or_226_nl), or_tmp_213, or_5189_cse);
  assign FpIntToFloat_17U_5U_10U_if_and_33_cse = cvt_else_and_cse & FpIntToFloat_17U_5U_10U_if_nor_10_cse
      & (mux_125_nl);
  assign FpIntToFloat_17U_5U_10U_if_nor_6_cse = ~(or_dcpl_15 | or_dcpl_30 | (cfg_out_precision_1_sva_st_154!=2'b10));
  assign or_243_nl = (cfg_out_precision_1_sva_st_154!=2'b10) | (~ and_1386_cse);
  assign mux_134_cse = MUX_s_1_2_2((or_243_nl), or_tmp_213, or_5189_cse);
  assign FpIntToFloat_17U_5U_10U_if_and_36_cse = cvt_else_and_cse & FpIntToFloat_17U_5U_10U_if_nor_10_cse
      & mux_134_cse;
  assign cvt_cvt_nand_cse = ~((cfg_proc_precision_rsci_d==2'b10));
  assign or_2943_nl = (and_dcpl_71 & or_5189_cse & (fsm_output[1])) | (and_dcpl_71
      & and_dcpl_73);
  assign cvt_16_NV_NVDLA_SDP_CORE_c_core_nvdla_float_h_ln670_assert_iExpoWidth_ge_oExpoWidth_4_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, or_2943_nl);
  assign and_550_cse = and_2186_cse & or_5189_cse & (fsm_output[1]);
  assign cvt_2_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln346_assert_oWidth_ge_aWidth_p_bWidth_1_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, and_550_cse);
  assign or_2944_nl = (and_dcpl_77 & and_dcpl_75 & (fsm_output[1])) | (and_dcpl_77
      & and_dcpl_80);
  assign cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, or_2944_nl);
  assign or_2945_nl = (and_dcpl_83 & and_dcpl_75 & (fsm_output[1])) | (and_dcpl_83
      & and_dcpl_80);
  assign cvt_1_NV_NVDLA_SDP_CORE_c_core_nvdla_int_h_ln402_assert_oWidth_le_iWidth_1_sig_mx0w1
      = MUX1HOT_s_1_1_2(1'b1, or_2945_nl);
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_2_sva_mx0w0
      = (~ (chn_in_rsci_d_mxwt[26:24])) + 3'b1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_2_sva_mx0w0
      = nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_2_sva_mx0w0[2:0];
  assign nl_cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_nl = ({1'b1 , (~ (chn_in_rsci_d_mxwt[30:23]))})
      + 9'b1110001;
  assign cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_nl = nl_cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_nl[8:0];
  assign cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_itm_8_1 = readslicef_9_1_8((cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_nl));
  assign nl_cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_nl = conv_u2u_7_8(chn_in_rsci_d_mxwt[30:24])
      + 8'b11001101;
  assign cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_nl = nl_cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_nl[7:0];
  assign cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1 = readslicef_8_1_7((cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_nl));
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_3_sva_mx0w0
      = (~ (chn_in_rsci_d_mxwt[58:56])) + 3'b1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_3_sva_mx0w0
      = nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_3_sva_mx0w0[2:0];
  assign nl_cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl = ({1'b1 , (~
      (chn_in_rsci_d_mxwt[62:55]))}) + 9'b1110001;
  assign cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl = nl_cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8:0];
  assign cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1 = readslicef_9_1_8((cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl));
  assign nl_cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl = conv_u2u_7_8(chn_in_rsci_d_mxwt[62:56])
      + 8'b11001101;
  assign cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl = nl_cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7:0];
  assign cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1 = readslicef_8_1_7((cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl));
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_4_sva_mx0w0
      = (~ (chn_in_rsci_d_mxwt[90:88])) + 3'b1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_4_sva_mx0w0
      = nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_4_sva_mx0w0[2:0];
  assign nl_cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl = ({1'b1 , (~
      (chn_in_rsci_d_mxwt[94:87]))}) + 9'b1110001;
  assign cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl = nl_cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8:0];
  assign cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1 = readslicef_9_1_8((cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl));
  assign nl_cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl = conv_u2u_7_8(chn_in_rsci_d_mxwt[94:88])
      + 8'b11001101;
  assign cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl = nl_cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7:0];
  assign cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1 = readslicef_8_1_7((cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl));
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_5_sva_mx0w0
      = (~ (chn_in_rsci_d_mxwt[122:120])) + 3'b1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_5_sva_mx0w0
      = nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_5_sva_mx0w0[2:0];
  assign nl_cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl = ({1'b1 , (~
      (chn_in_rsci_d_mxwt[126:119]))}) + 9'b1110001;
  assign cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl = nl_cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8:0];
  assign cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1 = readslicef_9_1_8((cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl));
  assign nl_cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl = conv_u2u_7_8(chn_in_rsci_d_mxwt[126:120])
      + 8'b11001101;
  assign cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl = nl_cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7:0];
  assign cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 = readslicef_8_1_7((cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl));
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_6_sva_mx0w0
      = (~ (chn_in_rsci_d_mxwt[154:152])) + 3'b1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_6_sva_mx0w0
      = nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_6_sva_mx0w0[2:0];
  assign nl_cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl = ({1'b1 , (~
      (chn_in_rsci_d_mxwt[158:151]))}) + 9'b1110001;
  assign cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl = nl_cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8:0];
  assign cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1 = readslicef_9_1_8((cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl));
  assign nl_cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl = conv_u2u_7_8(chn_in_rsci_d_mxwt[158:152])
      + 8'b11001101;
  assign cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl = nl_cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7:0];
  assign cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1 = readslicef_8_1_7((cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl));
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_7_sva_mx0w0
      = (~ (chn_in_rsci_d_mxwt[186:184])) + 3'b1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_7_sva_mx0w0
      = nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_7_sva_mx0w0[2:0];
  assign nl_cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl = ({1'b1 , (~
      (chn_in_rsci_d_mxwt[190:183]))}) + 9'b1110001;
  assign cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl = nl_cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8:0];
  assign cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1 = readslicef_9_1_8((cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl));
  assign nl_cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl = conv_u2u_7_8(chn_in_rsci_d_mxwt[190:184])
      + 8'b11001101;
  assign cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl = nl_cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7:0];
  assign cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 = readslicef_8_1_7((cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl));
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_8_sva_mx0w0
      = (~ (chn_in_rsci_d_mxwt[218:216])) + 3'b1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_8_sva_mx0w0
      = nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_8_sva_mx0w0[2:0];
  assign nl_cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl = ({1'b1 , (~
      (chn_in_rsci_d_mxwt[222:215]))}) + 9'b1110001;
  assign cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl = nl_cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8:0];
  assign cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1 = readslicef_9_1_8((cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl));
  assign nl_cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl = conv_u2u_7_8(chn_in_rsci_d_mxwt[222:216])
      + 8'b11001101;
  assign cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl = nl_cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7:0];
  assign cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 = readslicef_8_1_7((cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl));
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_9_sva_mx0w0
      = (~ (chn_in_rsci_d_mxwt[250:248])) + 3'b1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_9_sva_mx0w0
      = nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_9_sva_mx0w0[2:0];
  assign nl_cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl = ({1'b1 , (~
      (chn_in_rsci_d_mxwt[254:247]))}) + 9'b1110001;
  assign cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl = nl_cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8:0];
  assign cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1 = readslicef_9_1_8((cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl));
  assign nl_cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl = conv_u2u_7_8(chn_in_rsci_d_mxwt[254:248])
      + 8'b11001101;
  assign cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl = nl_cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7:0];
  assign cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 = readslicef_8_1_7((cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl));
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_10_sva_mx0w0
      = (~ (chn_in_rsci_d_mxwt[282:280])) + 3'b1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_10_sva_mx0w0
      = nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_10_sva_mx0w0[2:0];
  assign nl_cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl = ({1'b1 , (~
      (chn_in_rsci_d_mxwt[286:279]))}) + 9'b1110001;
  assign cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl = nl_cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl[8:0];
  assign cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1 = readslicef_9_1_8((cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_nl));
  assign nl_cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl = conv_u2u_7_8(chn_in_rsci_d_mxwt[286:280])
      + 8'b11001101;
  assign cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl = nl_cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl[7:0];
  assign cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1 = readslicef_8_1_7((cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_nl));
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_11_sva_mx0w0
      = (~ (chn_in_rsci_d_mxwt[314:312])) + 3'b1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_11_sva_mx0w0
      = nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_11_sva_mx0w0[2:0];
  assign nl_cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl = ({1'b1 , (~
      (chn_in_rsci_d_mxwt[318:311]))}) + 9'b1110001;
  assign cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl = nl_cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8:0];
  assign cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1 = readslicef_9_1_8((cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl));
  assign nl_cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl = conv_u2u_7_8(chn_in_rsci_d_mxwt[318:312])
      + 8'b11001101;
  assign cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl = nl_cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7:0];
  assign cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 = readslicef_8_1_7((cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl));
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_12_sva_mx0w0
      = (~ (chn_in_rsci_d_mxwt[346:344])) + 3'b1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_12_sva_mx0w0
      = nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_12_sva_mx0w0[2:0];
  assign nl_cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl = ({1'b1 , (~
      (chn_in_rsci_d_mxwt[350:343]))}) + 9'b1110001;
  assign cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl = nl_cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8:0];
  assign cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1 = readslicef_9_1_8((cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl));
  assign nl_cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl = conv_u2u_7_8(chn_in_rsci_d_mxwt[350:344])
      + 8'b11001101;
  assign cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl = nl_cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7:0];
  assign cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 = readslicef_8_1_7((cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl));
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_13_sva_mx0w0
      = (~ (chn_in_rsci_d_mxwt[378:376])) + 3'b1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_13_sva_mx0w0
      = nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_13_sva_mx0w0[2:0];
  assign nl_cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl = ({1'b1 , (~
      (chn_in_rsci_d_mxwt[382:375]))}) + 9'b1110001;
  assign cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl = nl_cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8:0];
  assign cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1 = readslicef_9_1_8((cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl));
  assign nl_cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl = conv_u2u_7_8(chn_in_rsci_d_mxwt[382:376])
      + 8'b11001101;
  assign cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl = nl_cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7:0];
  assign cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 = readslicef_8_1_7((cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl));
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_14_sva_mx0w0
      = (~ (chn_in_rsci_d_mxwt[410:408])) + 3'b1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_14_sva_mx0w0
      = nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_14_sva_mx0w0[2:0];
  assign nl_cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl = ({1'b1 , (~
      (chn_in_rsci_d_mxwt[414:407]))}) + 9'b1110001;
  assign cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl = nl_cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl[8:0];
  assign cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1 = readslicef_9_1_8((cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_nl));
  assign nl_cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl = conv_u2u_7_8(chn_in_rsci_d_mxwt[414:408])
      + 8'b11001101;
  assign cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl = nl_cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl[7:0];
  assign cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 = readslicef_8_1_7((cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_nl));
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_15_sva_mx0w0
      = (~ (chn_in_rsci_d_mxwt[442:440])) + 3'b1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_15_sva_mx0w0
      = nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_15_sva_mx0w0[2:0];
  assign nl_cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl = ({1'b1 , (~
      (chn_in_rsci_d_mxwt[446:439]))}) + 9'b1110001;
  assign cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl = nl_cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8:0];
  assign cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1 = readslicef_9_1_8((cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl));
  assign nl_cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl = conv_u2u_7_8(chn_in_rsci_d_mxwt[446:440])
      + 8'b11001101;
  assign cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl = nl_cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7:0];
  assign cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 = readslicef_8_1_7((cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl));
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_16_sva_mx0w0
      = (~ (chn_in_rsci_d_mxwt[474:472])) + 3'b1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_16_sva_mx0w0
      = nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_16_sva_mx0w0[2:0];
  assign nl_cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl = ({1'b1 , (~
      (chn_in_rsci_d_mxwt[478:471]))}) + 9'b1110001;
  assign cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl = nl_cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl[8:0];
  assign cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1 = readslicef_9_1_8((cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_nl));
  assign nl_cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl = conv_u2u_7_8(chn_in_rsci_d_mxwt[478:472])
      + 8'b11001101;
  assign cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl = nl_cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl[7:0];
  assign cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 = readslicef_8_1_7((cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_nl));
  assign nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_mx0w0
      = (~ (chn_in_rsci_d_mxwt[506:504])) + 3'b1;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_mx0w0
      = nl_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_mx0w0[2:0];
  assign nl_cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_nl = ({1'b1 , (~
      (chn_in_rsci_d_mxwt[510:503]))}) + 9'b1110001;
  assign cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_nl = nl_cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_nl[8:0];
  assign cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_itm_8_1 = readslicef_9_1_8((cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_nl));
  assign nl_cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_nl = conv_u2u_7_8(chn_in_rsci_d_mxwt[510:504])
      + 8'b11001101;
  assign cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_nl = nl_cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_nl[7:0];
  assign cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_itm_7_1 = readslicef_8_1_7((cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_nl));
  assign nl_cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_nl = conv_u2s_8_9(chn_in_rsci_d_mxwt[510:503])
      + 9'b101110001;
  assign cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_nl = nl_cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_nl[8:0];
  assign cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_itm_8_1 = readslicef_9_1_8((cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_nl));
  assign nl_cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl = conv_u2s_8_9(chn_in_rsci_d_mxwt[478:471])
      + 9'b101110001;
  assign cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl = nl_cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8:0];
  assign cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1 = readslicef_9_1_8((cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl));
  assign nl_cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl = conv_u2s_8_9(chn_in_rsci_d_mxwt[446:439])
      + 9'b101110001;
  assign cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl = nl_cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8:0];
  assign cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1 = readslicef_9_1_8((cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl));
  assign nl_cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl = conv_u2s_8_9(chn_in_rsci_d_mxwt[414:407])
      + 9'b101110001;
  assign cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl = nl_cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8:0];
  assign cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1 = readslicef_9_1_8((cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl));
  assign nl_cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl = conv_u2s_8_9(chn_in_rsci_d_mxwt[382:375])
      + 9'b101110001;
  assign cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl = nl_cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8:0];
  assign cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1 = readslicef_9_1_8((cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl));
  assign nl_cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl = conv_u2s_8_9(chn_in_rsci_d_mxwt[350:343])
      + 9'b101110001;
  assign cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl = nl_cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8:0];
  assign cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1 = readslicef_9_1_8((cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl));
  assign nl_cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl = conv_u2s_8_9(chn_in_rsci_d_mxwt[318:311])
      + 9'b101110001;
  assign cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl = nl_cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8:0];
  assign cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1 = readslicef_9_1_8((cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl));
  assign nl_cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl = conv_u2s_8_9(chn_in_rsci_d_mxwt[286:279])
      + 9'b101110001;
  assign cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl = nl_cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8:0];
  assign cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1 = readslicef_9_1_8((cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl));
  assign nl_cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl = conv_u2s_8_9(chn_in_rsci_d_mxwt[254:247])
      + 9'b101110001;
  assign cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl = nl_cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl[8:0];
  assign cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1 = readslicef_9_1_8((cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_nl));
  assign nl_cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl = conv_u2s_8_9(chn_in_rsci_d_mxwt[222:215])
      + 9'b101110001;
  assign cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl = nl_cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8:0];
  assign cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1 = readslicef_9_1_8((cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl));
  assign nl_cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl = conv_u2s_8_9(chn_in_rsci_d_mxwt[190:183])
      + 9'b101110001;
  assign cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl = nl_cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8:0];
  assign cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1 = readslicef_9_1_8((cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl));
  assign nl_cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl = conv_u2s_8_9(chn_in_rsci_d_mxwt[158:151])
      + 9'b101110001;
  assign cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl = nl_cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8:0];
  assign cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1 = readslicef_9_1_8((cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl));
  assign nl_cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl = conv_u2s_8_9(chn_in_rsci_d_mxwt[126:119])
      + 9'b101110001;
  assign cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl = nl_cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl[8:0];
  assign cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1 = readslicef_9_1_8((cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_nl));
  assign nl_cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl = conv_u2s_8_9(chn_in_rsci_d_mxwt[94:87])
      + 9'b101110001;
  assign cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl = nl_cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8:0];
  assign cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1 = readslicef_9_1_8((cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl));
  assign nl_cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl = conv_u2s_8_9(chn_in_rsci_d_mxwt[62:55])
      + 9'b101110001;
  assign cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl = nl_cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl[8:0];
  assign cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1 = readslicef_9_1_8((cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_nl));
  assign nl_cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_nl = conv_u2s_8_9(chn_in_rsci_d_mxwt[30:23])
      + 9'b101110001;
  assign cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_nl = nl_cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_nl[8:0];
  assign cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_itm_8_1 = readslicef_9_1_8((cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_nl));
  assign nl_cvt_1_FpMantRNE_24U_11U_else_acc_nl = (chn_idata_data_sva_1_27_0_1[22:13])
      + conv_u2u_1_10(FpMantRNE_24U_11U_else_carry_1_sva_2);
  assign cvt_1_FpMantRNE_24U_11U_else_acc_nl = nl_cvt_1_FpMantRNE_24U_11U_else_acc_nl[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_1_nl = MUX_v_10_2_2((FpMantDecShiftRight_23U_8U_10U_o_mant_sum_1_sva[9:0]),
      (cvt_1_FpMantRNE_24U_11U_else_acc_nl), cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_nl = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_1_nl),
      10'b1111111111, nand_164_cse));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_mx0w1
      = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_nl), 10'b1111111111,
      FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_1_lpi_1_dfm));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_47_nl = (~ cvt_1_FpMantRNE_24U_11U_else_and_svs_2)
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_1_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_48_nl = cvt_1_FpMantRNE_24U_11U_else_and_svs_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_1_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_nl =
      MUX1HOT_v_4_4_2(({3'b0 , (FpMantDecShiftRight_23U_8U_10U_o_mant_sum_1_sva[10])}),
      (chn_idata_data_sva_1_27_0_1[26:23]), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_sva_9[3:0]),
      4'b1110, {FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_ssc
      , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_47_nl) , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_48_nl)
      , nand_164_cse});
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_32_nl = ~ FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_1_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_nl
      = MUX_v_4_2_2(4'b0000, (FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_nl),
      (FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_32_nl));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_7_3_0_mx0w0 = MUX_v_4_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_nl),
      4'b1111, IsNaN_8U_23U_land_1_lpi_1_dfm_3);
  assign nl_cvt_2_FpMantRNE_24U_11U_else_acc_1_nl = (chn_idata_data_sva_1_59_31_1[23:14])
      + conv_u2u_1_10(FpMantRNE_24U_11U_else_carry_2_sva_2);
  assign cvt_2_FpMantRNE_24U_11U_else_acc_1_nl = nl_cvt_2_FpMantRNE_24U_11U_else_acc_1_nl[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_13_nl = MUX_v_10_2_2((FpMantDecShiftRight_23U_8U_10U_o_mant_sum_2_sva[9:0]),
      (cvt_2_FpMantRNE_24U_11U_else_acc_1_nl), cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_1_nl = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_13_nl),
      10'b1111111111, nand_162_cse));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_1_mx0w1
      = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_1_nl), 10'b1111111111,
      FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_2_lpi_1_dfm));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_49_nl = (~ cvt_2_FpMantRNE_24U_11U_else_and_1_svs_2)
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_3_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_50_nl = cvt_2_FpMantRNE_24U_11U_else_and_1_svs_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_3_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_1_nl
      = MUX1HOT_v_4_4_2(({3'b0 , (FpMantDecShiftRight_23U_8U_10U_o_mant_sum_2_sva[10])}),
      (chn_idata_data_sva_1_59_31_1[27:24]), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_sva_9[3:0]),
      4'b1110, {FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_1_ssc
      , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_49_nl) , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_50_nl)
      , nand_162_cse});
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_33_nl = ~ FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_2_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_2_nl
      = MUX_v_4_2_2(4'b0000, (FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_1_nl),
      (FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_33_nl));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_7_3_0_mx0w0 = MUX_v_4_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_2_nl),
      4'b1111, IsNaN_8U_23U_land_2_lpi_1_dfm_3);
  assign nl_cvt_3_FpMantRNE_24U_11U_else_acc_1_nl = (chn_idata_data_sva_1_91_63_1[23:14])
      + conv_u2u_1_10(FpMantRNE_24U_11U_else_carry_3_sva_2);
  assign cvt_3_FpMantRNE_24U_11U_else_acc_1_nl = nl_cvt_3_FpMantRNE_24U_11U_else_acc_1_nl[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_25_nl = MUX_v_10_2_2((FpMantDecShiftRight_23U_8U_10U_o_mant_sum_3_sva[9:0]),
      (cvt_3_FpMantRNE_24U_11U_else_acc_1_nl), cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_2_nl = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_25_nl),
      10'b1111111111, nand_160_cse));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_2_mx0w1
      = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_2_nl), 10'b1111111111,
      FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_3_lpi_1_dfm));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_51_nl = (~ cvt_3_FpMantRNE_24U_11U_else_and_1_svs_2)
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_5_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_52_nl = cvt_3_FpMantRNE_24U_11U_else_and_1_svs_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_5_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_2_nl
      = MUX1HOT_v_4_4_2(({3'b0 , (FpMantDecShiftRight_23U_8U_10U_o_mant_sum_3_sva[10])}),
      (chn_idata_data_sva_1_91_63_1[27:24]), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_sva_9[3:0]),
      4'b1110, {FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_2_ssc
      , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_51_nl) , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_52_nl)
      , nand_160_cse});
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_34_nl = ~ FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_3_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_4_nl
      = MUX_v_4_2_2(4'b0000, (FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_2_nl),
      (FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_34_nl));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_7_3_0_mx0w0 = MUX_v_4_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_4_nl),
      4'b1111, IsNaN_8U_23U_land_3_lpi_1_dfm_3);
  assign nl_cvt_4_FpMantRNE_24U_11U_else_acc_2_nl = (chn_idata_data_sva_1_123_95_1[23:14])
      + conv_u2u_1_10(FpMantRNE_24U_11U_else_carry_4_sva_2);
  assign cvt_4_FpMantRNE_24U_11U_else_acc_2_nl = nl_cvt_4_FpMantRNE_24U_11U_else_acc_2_nl[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_37_nl = MUX_v_10_2_2((FpMantDecShiftRight_23U_8U_10U_o_mant_sum_4_sva[9:0]),
      (cvt_4_FpMantRNE_24U_11U_else_acc_2_nl), cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_3_nl = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_37_nl),
      10'b1111111111, nand_158_cse));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_3_mx0w1
      = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_3_nl), 10'b1111111111,
      FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_4_lpi_1_dfm));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_53_nl = (~ cvt_4_FpMantRNE_24U_11U_else_and_2_svs_2)
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_7_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_54_nl = cvt_4_FpMantRNE_24U_11U_else_and_2_svs_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_7_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_3_nl
      = MUX1HOT_v_4_4_2(({3'b0 , (FpMantDecShiftRight_23U_8U_10U_o_mant_sum_4_sva[10])}),
      (chn_idata_data_sva_1_123_95_1[27:24]), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_sva_9[3:0]),
      4'b1110, {FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_3_ssc
      , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_53_nl) , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_54_nl)
      , nand_158_cse});
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_35_nl = ~ FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_4_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_6_nl
      = MUX_v_4_2_2(4'b0000, (FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_3_nl),
      (FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_35_nl));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_7_3_0_mx0w0 = MUX_v_4_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_6_nl),
      4'b1111, IsNaN_8U_23U_land_4_lpi_1_dfm_3);
  assign nl_cvt_5_FpMantRNE_24U_11U_else_acc_1_nl = (chn_idata_data_sva_1_155_127_1[23:14])
      + conv_u2u_1_10(FpMantRNE_24U_11U_else_carry_5_sva_2);
  assign cvt_5_FpMantRNE_24U_11U_else_acc_1_nl = nl_cvt_5_FpMantRNE_24U_11U_else_acc_1_nl[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_49_nl = MUX_v_10_2_2((FpMantDecShiftRight_23U_8U_10U_o_mant_sum_5_sva[9:0]),
      (cvt_5_FpMantRNE_24U_11U_else_acc_1_nl), cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_4_nl = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_49_nl),
      10'b1111111111, nand_156_cse));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_4_mx0w1
      = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_4_nl), 10'b1111111111,
      FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_5_lpi_1_dfm));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_55_nl = (~ cvt_5_FpMantRNE_24U_11U_else_and_1_svs_2)
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_9_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_56_nl = cvt_5_FpMantRNE_24U_11U_else_and_1_svs_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_9_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_4_nl
      = MUX1HOT_v_4_4_2(({3'b0 , (FpMantDecShiftRight_23U_8U_10U_o_mant_sum_5_sva[10])}),
      (chn_idata_data_sva_1_155_127_1[27:24]), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_sva_9[3:0]),
      4'b1110, {FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_4_ssc
      , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_55_nl) , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_56_nl)
      , nand_156_cse});
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_36_nl = ~ FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_5_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_8_nl
      = MUX_v_4_2_2(4'b0000, (FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_4_nl),
      (FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_36_nl));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_7_3_0_mx0w0 = MUX_v_4_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_8_nl),
      4'b1111, nor_1099_cse);
  assign nl_cvt_6_FpMantRNE_24U_11U_else_acc_2_nl = (chn_idata_data_sva_1_187_159_1[23:14])
      + conv_u2u_1_10(FpMantRNE_24U_11U_else_carry_6_sva_2);
  assign cvt_6_FpMantRNE_24U_11U_else_acc_2_nl = nl_cvt_6_FpMantRNE_24U_11U_else_acc_2_nl[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_61_nl = MUX_v_10_2_2((FpMantDecShiftRight_23U_8U_10U_o_mant_sum_6_sva[9:0]),
      (cvt_6_FpMantRNE_24U_11U_else_acc_2_nl), cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_5_nl = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_61_nl),
      10'b1111111111, nand_153_cse));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_5_mx0w1
      = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_5_nl), 10'b1111111111,
      FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_6_lpi_1_dfm));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_57_nl = (~ cvt_6_FpMantRNE_24U_11U_else_and_2_svs_2)
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_11_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_58_nl = cvt_6_FpMantRNE_24U_11U_else_and_2_svs_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_11_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_5_nl
      = MUX1HOT_v_4_4_2(({3'b0 , (FpMantDecShiftRight_23U_8U_10U_o_mant_sum_6_sva[10])}),
      (chn_idata_data_sva_1_187_159_1[27:24]), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_sva_9[3:0]),
      4'b1110, {FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_5_ssc
      , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_57_nl) , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_58_nl)
      , nand_153_cse});
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_37_nl = ~ FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_6_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_10_nl
      = MUX_v_4_2_2(4'b0000, (FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_5_nl),
      (FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_37_nl));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_7_3_0_mx0w0 = MUX_v_4_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_10_nl),
      4'b1111, IsNaN_8U_23U_land_6_lpi_1_dfm_3);
  assign nl_cvt_7_FpMantRNE_24U_11U_else_acc_2_nl = (chn_idata_data_sva_1_219_191_1[23:14])
      + conv_u2u_1_10(FpMantRNE_24U_11U_else_carry_7_sva_2);
  assign cvt_7_FpMantRNE_24U_11U_else_acc_2_nl = nl_cvt_7_FpMantRNE_24U_11U_else_acc_2_nl[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_73_nl = MUX_v_10_2_2((FpMantDecShiftRight_23U_8U_10U_o_mant_sum_7_sva[9:0]),
      (cvt_7_FpMantRNE_24U_11U_else_acc_2_nl), cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_6_nl = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_73_nl),
      10'b1111111111, nand_151_cse));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_6_mx0w1
      = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_6_nl), 10'b1111111111,
      FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_7_lpi_1_dfm));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_59_nl = (~ cvt_7_FpMantRNE_24U_11U_else_and_2_svs_2)
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_13_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_60_nl = cvt_7_FpMantRNE_24U_11U_else_and_2_svs_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_13_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_6_nl
      = MUX1HOT_v_4_4_2(({3'b0 , (FpMantDecShiftRight_23U_8U_10U_o_mant_sum_7_sva[10])}),
      (chn_idata_data_sva_1_219_191_1[27:24]), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_sva_9[3:0]),
      4'b1110, {FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_6_ssc
      , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_59_nl) , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_60_nl)
      , nand_151_cse});
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_38_nl = ~ FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_7_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_12_nl
      = MUX_v_4_2_2(4'b0000, (FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_6_nl),
      (FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_38_nl));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_7_3_0_mx0w0 = MUX_v_4_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_12_nl),
      4'b1111, IsNaN_8U_23U_land_7_lpi_1_dfm_3);
  assign nl_cvt_8_FpMantRNE_24U_11U_else_acc_3_nl = (chn_idata_data_sva_1_251_223_1[23:14])
      + conv_u2u_1_10(FpMantRNE_24U_11U_else_carry_8_sva_2);
  assign cvt_8_FpMantRNE_24U_11U_else_acc_3_nl = nl_cvt_8_FpMantRNE_24U_11U_else_acc_3_nl[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_85_nl = MUX_v_10_2_2((FpMantDecShiftRight_23U_8U_10U_o_mant_sum_8_sva[9:0]),
      (cvt_8_FpMantRNE_24U_11U_else_acc_3_nl), cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_7_nl = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_85_nl),
      10'b1111111111, nand_149_cse));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_7_mx0w1
      = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_7_nl), 10'b1111111111,
      FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_8_lpi_1_dfm));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_61_nl = (~ cvt_8_FpMantRNE_24U_11U_else_and_3_svs_2)
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_15_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_62_nl = cvt_8_FpMantRNE_24U_11U_else_and_3_svs_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_15_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_7_nl
      = MUX1HOT_v_4_4_2(({3'b0 , (FpMantDecShiftRight_23U_8U_10U_o_mant_sum_8_sva[10])}),
      (chn_idata_data_sva_1_251_223_1[27:24]), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_sva_9[3:0]),
      4'b1110, {FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_7_ssc
      , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_61_nl) , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_62_nl)
      , nand_149_cse});
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_39_nl = ~ FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_8_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_14_nl
      = MUX_v_4_2_2(4'b0000, (FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_7_nl),
      (FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_39_nl));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_7_3_0_mx0w0 = MUX_v_4_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_14_nl),
      4'b1111, IsNaN_8U_23U_land_8_lpi_1_dfm_3);
  assign nl_cvt_9_FpMantRNE_24U_11U_else_acc_1_nl = (chn_idata_data_sva_1_283_255_1[23:14])
      + conv_u2u_1_10(FpMantRNE_24U_11U_else_carry_9_sva_2);
  assign cvt_9_FpMantRNE_24U_11U_else_acc_1_nl = nl_cvt_9_FpMantRNE_24U_11U_else_acc_1_nl[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_97_nl = MUX_v_10_2_2((FpMantDecShiftRight_23U_8U_10U_o_mant_sum_9_sva[9:0]),
      (cvt_9_FpMantRNE_24U_11U_else_acc_1_nl), cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_8_nl = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_97_nl),
      10'b1111111111, nand_147_cse));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_8_mx0w1
      = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_8_nl), 10'b1111111111,
      FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_9_lpi_1_dfm));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_63_nl = (~ cvt_9_FpMantRNE_24U_11U_else_and_1_svs_2)
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_17_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_64_nl = cvt_9_FpMantRNE_24U_11U_else_and_1_svs_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_17_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_8_nl
      = MUX1HOT_v_4_4_2(({3'b0 , (FpMantDecShiftRight_23U_8U_10U_o_mant_sum_9_sva[10])}),
      (chn_idata_data_sva_1_283_255_1[27:24]), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_sva_9[3:0]),
      4'b1110, {FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_8_ssc
      , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_63_nl) , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_64_nl)
      , nand_147_cse});
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_40_nl = ~ FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_9_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_16_nl
      = MUX_v_4_2_2(4'b0000, (FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_8_nl),
      (FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_40_nl));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_7_3_0_mx0w0 = MUX_v_4_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_16_nl),
      4'b1111, IsNaN_8U_23U_land_9_lpi_1_dfm_3);
  assign nl_cvt_10_FpMantRNE_24U_11U_else_acc_2_nl = (chn_idata_data_sva_1_315_287_1[23:14])
      + conv_u2u_1_10(FpMantRNE_24U_11U_else_carry_10_sva_2);
  assign cvt_10_FpMantRNE_24U_11U_else_acc_2_nl = nl_cvt_10_FpMantRNE_24U_11U_else_acc_2_nl[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_109_nl = MUX_v_10_2_2((FpMantDecShiftRight_23U_8U_10U_o_mant_sum_10_sva[9:0]),
      (cvt_10_FpMantRNE_24U_11U_else_acc_2_nl), cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_9_nl = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_109_nl),
      10'b1111111111, nand_145_cse));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_9_mx0w1
      = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_9_nl), 10'b1111111111,
      FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_10_lpi_1_dfm));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_65_nl = (~ cvt_10_FpMantRNE_24U_11U_else_and_2_svs_2)
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_19_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_66_nl = cvt_10_FpMantRNE_24U_11U_else_and_2_svs_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_19_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_9_nl
      = MUX1HOT_v_4_4_2(({3'b0 , (FpMantDecShiftRight_23U_8U_10U_o_mant_sum_10_sva[10])}),
      (chn_idata_data_sva_1_315_287_1[27:24]), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_sva_9[3:0]),
      4'b1110, {FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_9_ssc
      , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_65_nl) , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_66_nl)
      , nand_145_cse});
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_41_nl = ~ FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_10_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_18_nl
      = MUX_v_4_2_2(4'b0000, (FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_9_nl),
      (FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_41_nl));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_7_3_0_mx0w0 = MUX_v_4_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_18_nl),
      4'b1111, IsNaN_8U_23U_land_10_lpi_1_dfm_3);
  assign nl_cvt_11_FpMantRNE_24U_11U_else_acc_2_nl = (chn_idata_data_sva_1_347_319_1[23:14])
      + conv_u2u_1_10(FpMantRNE_24U_11U_else_carry_11_sva_2);
  assign cvt_11_FpMantRNE_24U_11U_else_acc_2_nl = nl_cvt_11_FpMantRNE_24U_11U_else_acc_2_nl[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_121_nl = MUX_v_10_2_2((FpMantDecShiftRight_23U_8U_10U_o_mant_sum_11_sva[9:0]),
      (cvt_11_FpMantRNE_24U_11U_else_acc_2_nl), cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_10_nl = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_121_nl),
      10'b1111111111, nand_143_cse));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_10_mx0w1
      = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_10_nl), 10'b1111111111,
      FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_11_lpi_1_dfm));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_67_nl = (~ cvt_11_FpMantRNE_24U_11U_else_and_2_svs_2)
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_21_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_68_nl = cvt_11_FpMantRNE_24U_11U_else_and_2_svs_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_21_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_10_nl
      = MUX1HOT_v_4_4_2(({3'b0 , (FpMantDecShiftRight_23U_8U_10U_o_mant_sum_11_sva[10])}),
      (chn_idata_data_sva_1_347_319_1[27:24]), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_sva_9[3:0]),
      4'b1110, {FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_10_ssc
      , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_67_nl) , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_68_nl)
      , nand_143_cse});
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_42_nl = ~ FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_11_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_20_nl
      = MUX_v_4_2_2(4'b0000, (FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_10_nl),
      (FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_42_nl));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_7_3_0_mx0w0 = MUX_v_4_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_20_nl),
      4'b1111, IsNaN_8U_23U_land_11_lpi_1_dfm_3);
  assign nl_cvt_12_FpMantRNE_24U_11U_else_acc_3_nl = (chn_idata_data_sva_1_379_351_1[23:14])
      + conv_u2u_1_10(FpMantRNE_24U_11U_else_carry_12_sva_2);
  assign cvt_12_FpMantRNE_24U_11U_else_acc_3_nl = nl_cvt_12_FpMantRNE_24U_11U_else_acc_3_nl[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_133_nl = MUX_v_10_2_2((FpMantDecShiftRight_23U_8U_10U_o_mant_sum_12_sva[9:0]),
      (cvt_12_FpMantRNE_24U_11U_else_acc_3_nl), cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_11_nl = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_133_nl),
      10'b1111111111, nand_141_cse));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_11_mx0w1
      = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_11_nl), 10'b1111111111,
      FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_12_lpi_1_dfm));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_69_nl = (~ cvt_12_FpMantRNE_24U_11U_else_and_3_svs_2)
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_23_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_70_nl = cvt_12_FpMantRNE_24U_11U_else_and_3_svs_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_23_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_11_nl
      = MUX1HOT_v_4_4_2(({3'b0 , (FpMantDecShiftRight_23U_8U_10U_o_mant_sum_12_sva[10])}),
      (chn_idata_data_sva_1_379_351_1[27:24]), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_sva_9[3:0]),
      4'b1110, {FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_11_ssc
      , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_69_nl) , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_70_nl)
      , nand_141_cse});
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_43_nl = ~ FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_12_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_22_nl
      = MUX_v_4_2_2(4'b0000, (FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_11_nl),
      (FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_43_nl));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_7_3_0_mx0w0 = MUX_v_4_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_22_nl),
      4'b1111, IsNaN_8U_23U_land_12_lpi_1_dfm_3);
  assign nl_cvt_13_FpMantRNE_24U_11U_else_acc_2_nl = (chn_idata_data_sva_1_411_383_1[23:14])
      + conv_u2u_1_10(FpMantRNE_24U_11U_else_carry_13_sva_2);
  assign cvt_13_FpMantRNE_24U_11U_else_acc_2_nl = nl_cvt_13_FpMantRNE_24U_11U_else_acc_2_nl[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_145_nl = MUX_v_10_2_2((FpMantDecShiftRight_23U_8U_10U_o_mant_sum_13_sva[9:0]),
      (cvt_13_FpMantRNE_24U_11U_else_acc_2_nl), cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_12_nl = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_145_nl),
      10'b1111111111, nand_139_cse));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_12_mx0w1
      = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_12_nl), 10'b1111111111,
      FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_13_lpi_1_dfm));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_71_nl = (~ cvt_13_FpMantRNE_24U_11U_else_and_2_svs_2)
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_25_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_72_nl = cvt_13_FpMantRNE_24U_11U_else_and_2_svs_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_25_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_12_nl
      = MUX1HOT_v_4_4_2(({3'b0 , (FpMantDecShiftRight_23U_8U_10U_o_mant_sum_13_sva[10])}),
      (chn_idata_data_sva_1_411_383_1[27:24]), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_sva_9[3:0]),
      4'b1110, {FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_12_ssc
      , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_71_nl) , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_72_nl)
      , nand_139_cse});
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_44_nl = ~ FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_13_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_24_nl
      = MUX_v_4_2_2(4'b0000, (FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_12_nl),
      (FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_44_nl));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_7_3_0_mx0w0 = MUX_v_4_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_24_nl),
      4'b1111, IsNaN_8U_23U_land_13_lpi_1_dfm_3);
  assign nl_cvt_14_FpMantRNE_24U_11U_else_acc_3_nl = (chn_idata_data_sva_1_443_415_1[23:14])
      + conv_u2u_1_10(FpMantRNE_24U_11U_else_carry_14_sva_2);
  assign cvt_14_FpMantRNE_24U_11U_else_acc_3_nl = nl_cvt_14_FpMantRNE_24U_11U_else_acc_3_nl[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_157_nl = MUX_v_10_2_2((FpMantDecShiftRight_23U_8U_10U_o_mant_sum_14_sva[9:0]),
      (cvt_14_FpMantRNE_24U_11U_else_acc_3_nl), cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_13_nl = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_157_nl),
      10'b1111111111, nand_137_cse));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_13_mx0w1
      = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_13_nl), 10'b1111111111,
      FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_14_lpi_1_dfm));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_73_nl = (~ cvt_14_FpMantRNE_24U_11U_else_and_3_svs_2)
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_27_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_74_nl = cvt_14_FpMantRNE_24U_11U_else_and_3_svs_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_27_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_13_nl
      = MUX1HOT_v_4_4_2(({3'b0 , (FpMantDecShiftRight_23U_8U_10U_o_mant_sum_14_sva[10])}),
      (chn_idata_data_sva_1_443_415_1[27:24]), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_sva_9[3:0]),
      4'b1110, {FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_13_ssc
      , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_73_nl) , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_74_nl)
      , nand_137_cse});
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_45_nl = ~ FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_14_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_26_nl
      = MUX_v_4_2_2(4'b0000, (FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_13_nl),
      (FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_45_nl));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_7_3_0_mx0w0 = MUX_v_4_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_26_nl),
      4'b1111, IsNaN_8U_23U_land_14_lpi_1_dfm_3);
  assign nl_cvt_15_FpMantRNE_24U_11U_else_acc_3_nl = (chn_idata_data_sva_1_475_447_1[23:14])
      + conv_u2u_1_10(FpMantRNE_24U_11U_else_carry_15_sva_2);
  assign cvt_15_FpMantRNE_24U_11U_else_acc_3_nl = nl_cvt_15_FpMantRNE_24U_11U_else_acc_3_nl[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_169_nl = MUX_v_10_2_2((FpMantDecShiftRight_23U_8U_10U_o_mant_sum_15_sva[9:0]),
      (cvt_15_FpMantRNE_24U_11U_else_acc_3_nl), cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_14_nl = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_169_nl),
      10'b1111111111, nand_135_cse));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_14_mx0w1
      = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_14_nl), 10'b1111111111,
      FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_15_lpi_1_dfm));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_75_nl = (~ cvt_15_FpMantRNE_24U_11U_else_and_3_svs_2)
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_29_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_76_nl = cvt_15_FpMantRNE_24U_11U_else_and_3_svs_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_29_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_14_nl
      = MUX1HOT_v_4_4_2(({3'b0 , (FpMantDecShiftRight_23U_8U_10U_o_mant_sum_15_sva[10])}),
      (chn_idata_data_sva_1_475_447_1[27:24]), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_sva_9[3:0]),
      4'b1110, {FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_14_ssc
      , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_75_nl) , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_76_nl)
      , nand_135_cse});
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_46_nl = ~ FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_15_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_28_nl
      = MUX_v_4_2_2(4'b0000, (FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_14_nl),
      (FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_46_nl));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_7_3_0_mx0w0 = MUX_v_4_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_28_nl),
      4'b1111, IsNaN_8U_23U_land_15_lpi_1_dfm_3);
  assign nl_cvt_16_FpMantRNE_24U_11U_else_acc_4_nl = (chn_idata_data_sva_1_507_479_1[23:14])
      + conv_u2u_1_10(FpMantRNE_24U_11U_else_carry_sva_2);
  assign cvt_16_FpMantRNE_24U_11U_else_acc_4_nl = nl_cvt_16_FpMantRNE_24U_11U_else_acc_4_nl[9:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_181_nl = MUX_v_10_2_2((FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva[9:0]),
      (cvt_16_FpMantRNE_24U_11U_else_acc_4_nl), cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_15_nl = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_mux_181_nl),
      10'b1111111111, nand_133_cse));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_15_mx0w1
      = ~(MUX_v_10_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_15_nl), 10'b1111111111,
      FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_lpi_1_dfm));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_77_nl = (~ cvt_16_FpMantRNE_24U_11U_else_and_4_svs_2)
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_31_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_78_nl = cvt_16_FpMantRNE_24U_11U_else_and_4_svs_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_and_31_m1c;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_15_nl
      = MUX1HOT_v_4_4_2(({3'b0 , (FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva[10])}),
      (chn_idata_data_sva_1_507_479_1[27:24]), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_sva_9[3:0]),
      4'b1110, {FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_15_ssc
      , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_77_nl) , (FpWidthDec_8U_23U_5U_10U_1U_1U_and_78_nl)
      , nand_133_cse});
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_47_nl = ~ FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_lpi_1_dfm;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_30_nl
      = MUX_v_4_2_2(4'b0000, (FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_mux1h_15_nl),
      (FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_not_47_nl));
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_7_3_0_mx0w0 = MUX_v_4_2_2((FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_and_30_nl),
      4'b1111, IsNaN_8U_23U_land_lpi_1_dfm_3);
  assign cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_nor_4_cse = ~((cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_acc_tmp[16])
      | cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_and_1_tmp);
  assign IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0 = ~(cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_nor_4_cse
      | cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_nor_tmp);
  assign cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_nor_2_nl = ~(MUX_v_15_2_2((cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_acc_tmp[15:1]),
      15'b111111111111111, cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_nor_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_mx0w0 = ~(MUX_v_15_2_2((cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_nor_2_nl),
      15'b111111111111111, cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_and_1_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_0_1_sva_mx0w0 = ~((~((cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_acc_tmp[0])
      | cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_nor_tmp)) | cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_and_1_tmp);
  assign cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_tmp = ~(IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0
      | (IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_mx0w0!=15'b000000000000000) | IntShiftRightSat_49U_6U_17U_o_0_1_sva_mx0w0);
  assign cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse = ~((cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[16])
      | cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp);
  assign IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0 = ~(cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse
      | cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp);
  assign cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_nor_7_nl = ~(MUX_v_15_2_2((cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[15:1]),
      15'b111111111111111, cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_mx0w0 = ~(MUX_v_15_2_2((cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_nor_7_nl),
      15'b111111111111111, cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_0_2_sva_mx0w0 = ~((~((cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[0])
      | cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp)) | cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp);
  assign cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp = ~(IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0
      | (IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_mx0w0!=15'b000000000000000) | IntShiftRightSat_49U_6U_17U_o_0_2_sva_mx0w0);
  assign cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp
      = IntShiftRightSat_49U_6U_17U_i_2_sva_mx0w0 != conv_s2s_17_49({IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0
      , IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_mx0w0 , IntShiftRightSat_49U_6U_17U_o_0_2_sva_mx0w0});
  assign cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse = ~((cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[16])
      | cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp);
  assign IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0 = ~(cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse
      | cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp);
  assign cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_nor_7_nl = ~(MUX_v_15_2_2((cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[15:1]),
      15'b111111111111111, cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_mx0w0 = ~(MUX_v_15_2_2((cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_nor_7_nl),
      15'b111111111111111, cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_0_3_sva_mx0w0 = ~((~((cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[0])
      | cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp)) | cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp);
  assign cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp = ~(IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0
      | (IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_mx0w0!=15'b000000000000000) | IntShiftRightSat_49U_6U_17U_o_0_3_sva_mx0w0);
  assign cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse = ~((cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[16])
      | cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp);
  assign IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0 = ~(cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse
      | cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp);
  assign cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl = ~(MUX_v_15_2_2((cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[15:1]),
      15'b111111111111111, cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_mx0w0 = ~(MUX_v_15_2_2((cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl),
      15'b111111111111111, cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_0_4_sva_mx0w0 = ~((~((cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[0])
      | cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp)) | cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp);
  assign cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp
      = IntShiftRightSat_49U_6U_17U_i_4_sva_mx0w1 != conv_s2s_17_49({IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0
      , IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_mx0w0 , IntShiftRightSat_49U_6U_17U_o_0_4_sva_mx0w0});
  assign cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp
      = IntShiftRightSat_49U_6U_17U_i_3_sva_mx0w0 != conv_s2s_17_49({IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0
      , IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_mx0w0 , IntShiftRightSat_49U_6U_17U_o_0_3_sva_mx0w0});
  assign cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse = ~((cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[16])
      | cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp);
  assign IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0 = ~(cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse
      | cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp);
  assign cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_nor_7_nl = ~(MUX_v_15_2_2((cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[15:1]),
      15'b111111111111111, cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_mx0w0 = ~(MUX_v_15_2_2((cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_nor_7_nl),
      15'b111111111111111, cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_0_5_sva_mx0w0 = ~((~((cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[0])
      | cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp)) | cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp);
  assign cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp = ~(IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0
      | (IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_mx0w0!=15'b000000000000000) | IntShiftRightSat_49U_6U_17U_o_0_5_sva_mx0w0);
  assign cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse = ~((cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[16])
      | cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp);
  assign IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0 = ~(cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse
      | cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp);
  assign cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl = ~(MUX_v_15_2_2((cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[15:1]),
      15'b111111111111111, cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_mx0w0 = ~(MUX_v_15_2_2((cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl),
      15'b111111111111111, cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_0_6_sva_mx0w0 = ~((~((cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[0])
      | cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp)) | cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp);
  assign cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp
      = IntShiftRightSat_49U_6U_17U_i_6_sva_mx0w1 != conv_s2s_17_49({IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0
      , IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_mx0w0 , IntShiftRightSat_49U_6U_17U_o_0_6_sva_mx0w0});
  assign cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse = ~((cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[16])
      | cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp);
  assign IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0 = ~(cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse
      | cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp);
  assign cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl = ~(MUX_v_15_2_2((cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[15:1]),
      15'b111111111111111, cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_mx0w0 = ~(MUX_v_15_2_2((cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl),
      15'b111111111111111, cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_0_7_sva_mx0w0 = ~((~((cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[0])
      | cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp)) | cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp);
  assign cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse = ~((cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[16])
      | cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp);
  assign IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0 = ~(cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse
      | cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp);
  assign cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_nor_17_nl = ~(MUX_v_15_2_2((cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[15:1]),
      15'b111111111111111, cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_mx0w0 = ~(MUX_v_15_2_2((cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_nor_17_nl),
      15'b111111111111111, cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_0_8_sva_mx0w0 = ~((~((cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[0])
      | cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp)) | cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp);
  assign cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp
      = IntShiftRightSat_49U_6U_17U_i_8_sva_mx0w1 != conv_s2s_17_49({IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0
      , IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_mx0w0 , IntShiftRightSat_49U_6U_17U_o_0_8_sva_mx0w0});
  assign cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp
      = IntShiftRightSat_49U_6U_17U_i_7_sva_mx0w1 != conv_s2s_17_49({IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0
      , IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_mx0w0 , IntShiftRightSat_49U_6U_17U_o_0_7_sva_mx0w0});
  assign cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp
      = IntShiftRightSat_49U_6U_17U_i_5_sva_mx0w0 != conv_s2s_17_49({IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0
      , IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_mx0w0 , IntShiftRightSat_49U_6U_17U_o_0_5_sva_mx0w0});
  assign cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse = ~((cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[16])
      | cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp);
  assign IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0 = ~(cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse
      | cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp);
  assign cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_nor_7_nl = ~(MUX_v_15_2_2((cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[15:1]),
      15'b111111111111111, cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_mx0w0 = ~(MUX_v_15_2_2((cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_nor_7_nl),
      15'b111111111111111, cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_0_9_sva_mx0w0 = ~((~((cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[0])
      | cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp)) | cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp);
  assign cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp = ~(IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0
      | (IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_mx0w0!=15'b000000000000000) | IntShiftRightSat_49U_6U_17U_o_0_9_sva_mx0w0);
  assign cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse = ~((cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[16])
      | cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp);
  assign IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0 = ~(cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse
      | cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp);
  assign cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl = ~(MUX_v_15_2_2((cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[15:1]),
      15'b111111111111111, cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_mx0w0 = ~(MUX_v_15_2_2((cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl),
      15'b111111111111111, cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_0_10_sva_mx0w0 = ~((~((cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[0])
      | cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp)) | cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp);
  assign cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse = ~((cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[16])
      | cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp);
  assign IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0 = ~(cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse
      | cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp);
  assign cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl = ~(MUX_v_15_2_2((cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[15:1]),
      15'b111111111111111, cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_mx0w0 = ~(MUX_v_15_2_2((cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl),
      15'b111111111111111, cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_0_11_sva_mx0w0 = ~((~((cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[0])
      | cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp)) | cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp);
  assign cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse = ~((cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[16])
      | cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp);
  assign IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0 = ~(cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse
      | cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp);
  assign cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_nor_17_nl = ~(MUX_v_15_2_2((cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[15:1]),
      15'b111111111111111, cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_mx0w0 = ~(MUX_v_15_2_2((cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_nor_17_nl),
      15'b111111111111111, cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_0_12_sva_mx0w0 = ~((~((cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[0])
      | cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp)) | cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp);
  assign cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse = ~((cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[16])
      | cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp);
  assign IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0 = ~(cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse
      | cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp);
  assign cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl = ~(MUX_v_15_2_2((cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[15:1]),
      15'b111111111111111, cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_mx0w0 = ~(MUX_v_15_2_2((cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_nor_12_nl),
      15'b111111111111111, cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_0_13_sva_mx0w0 = ~((~((cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[0])
      | cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp)) | cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp);
  assign cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse = ~((cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[16])
      | cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp);
  assign IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0 = ~(cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse
      | cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp);
  assign cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_nor_17_nl = ~(MUX_v_15_2_2((cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[15:1]),
      15'b111111111111111, cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_mx0w0 = ~(MUX_v_15_2_2((cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_nor_17_nl),
      15'b111111111111111, cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_0_14_sva_mx0w0 = ~((~((cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[0])
      | cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp)) | cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp);
  assign cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse = ~((cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[16])
      | cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp);
  assign IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0 = ~(cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse
      | cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp);
  assign cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_nor_17_nl = ~(MUX_v_15_2_2((cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[15:1]),
      15'b111111111111111, cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_mx0w0 = ~(MUX_v_15_2_2((cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_nor_17_nl),
      15'b111111111111111, cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_0_15_sva_mx0w0 = ~((~((cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[0])
      | cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp)) | cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp);
  assign cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_nor_24_cse = ~((cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_acc_4_tmp[16])
      | cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_and_9_tmp);
  assign IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0 = ~(cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_nor_24_cse
      | cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_nor_20_tmp);
  assign cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_nor_22_nl = ~(MUX_v_15_2_2((cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_acc_4_tmp[15:1]),
      15'b111111111111111, cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_nor_20_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_15_1_sva_mx0w0 = ~(MUX_v_15_2_2((cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_nor_22_nl),
      15'b111111111111111, cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_and_9_tmp));
  assign IntShiftRightSat_49U_6U_17U_o_0_sva_mx0w0 = ~((~((cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_acc_4_tmp[0])
      | cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_nor_20_tmp)) | cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_and_9_tmp);
  assign cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp
      = IntShiftRightSat_49U_6U_17U_i_9_sva_mx0w0 != conv_s2s_17_49({IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0
      , IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_mx0w0 , IntShiftRightSat_49U_6U_17U_o_0_9_sva_mx0w0});
  assign cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_tmp
      = IntShiftRightSat_49U_6U_17U_i_1_sva_mx0w0 != conv_s2s_17_49({IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0
      , IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_mx0w0 , IntShiftRightSat_49U_6U_17U_o_0_1_sva_mx0w0});
  assign FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_mx0w0 = ~((~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_1_sva[0])
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_1_sva)) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_1_sva);
  assign cvt_1_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_nl
      = (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_1_sva[25]) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_1_sva))
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_1_sva;
  assign nl_cvt_1_FpFloatToInt_16U_5U_10U_if_acc_nl = ({1'b1 , (cvt_1_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_nl)
      , (~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_1_sva[23:14]))}) + 12'b1;
  assign cvt_1_FpFloatToInt_16U_5U_10U_if_acc_nl = nl_cvt_1_FpFloatToInt_16U_5U_10U_if_acc_nl[11:0];
  assign cvt_1_FpFloatToInt_16U_5U_10U_if_acc_itm_11_1 = readslicef_12_1_11((cvt_1_FpFloatToInt_16U_5U_10U_if_acc_nl));
  assign IsNaN_5U_10U_land_1_lpi_1_dfm_mx0w0 = ~(IsNaN_5U_10U_nor_itm_2 | IsNaN_5U_10U_IsNaN_5U_10U_nand_itm_2);
  assign FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_mx0w0 = ~((~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_2_sva[0])
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_2_sva)) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_2_sva);
  assign cvt_2_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_1_nl
      = (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_2_sva[25]) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_2_sva))
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_2_sva;
  assign nl_cvt_2_FpFloatToInt_16U_5U_10U_if_acc_1_nl = ({1'b1 , (cvt_2_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_1_nl)
      , (~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_2_sva[23:14]))}) + 12'b1;
  assign cvt_2_FpFloatToInt_16U_5U_10U_if_acc_1_nl = nl_cvt_2_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11:0];
  assign cvt_2_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1 = readslicef_12_1_11((cvt_2_FpFloatToInt_16U_5U_10U_if_acc_1_nl));
  assign IsNaN_5U_10U_land_2_lpi_1_dfm_mx0w0 = ~(IsNaN_5U_10U_nor_1_itm_2 | IsNaN_5U_10U_IsNaN_5U_10U_nand_1_itm_2);
  assign FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_mx0w0 = ~((~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_3_sva[0])
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_3_sva)) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_3_sva);
  assign nl_cvt_3_IntSaturation_17U_8U_if_acc_1_nl = conv_s2u_10_11({(~ IntShiftRightSat_49U_6U_17U_o_16_3_sva_3)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_2[14:6]))}) + 11'b1;
  assign cvt_3_IntSaturation_17U_8U_if_acc_1_nl = nl_cvt_3_IntSaturation_17U_8U_if_acc_1_nl[10:0];
  assign cvt_3_IntSaturation_17U_8U_if_acc_1_itm_10_1 = readslicef_11_1_10((cvt_3_IntSaturation_17U_8U_if_acc_1_nl));
  assign cvt_3_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_1_nl
      = (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_3_sva[25]) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_3_sva))
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_3_sva;
  assign nl_cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_nl = ({1'b1 , (cvt_3_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_1_nl)
      , (~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_3_sva[23:14]))}) + 12'b1;
  assign cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_nl = nl_cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11:0];
  assign cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1 = readslicef_12_1_11((cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_nl));
  assign FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_mx0w0 = ~((~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_4_sva[0])
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_4_sva)) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_4_sva);
  assign cvt_4_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl
      = (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_4_sva[25]) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_4_sva))
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_4_sva;
  assign nl_cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_nl = ({1'b1 , (cvt_4_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl)
      , (~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_4_sva[23:14]))}) + 12'b1;
  assign cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_nl = nl_cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11:0];
  assign cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1 = readslicef_12_1_11((cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_nl));
  assign FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_mx0w0 = ~((~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_5_sva[0])
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_5_sva)) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_5_sva);
  assign nl_cvt_5_IntSaturation_17U_8U_if_acc_1_nl = conv_s2u_10_11({(~ IntShiftRightSat_49U_6U_17U_o_16_5_sva_3)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_2[14:6]))}) + 11'b1;
  assign cvt_5_IntSaturation_17U_8U_if_acc_1_nl = nl_cvt_5_IntSaturation_17U_8U_if_acc_1_nl[10:0];
  assign cvt_5_IntSaturation_17U_8U_if_acc_1_itm_10_1 = readslicef_11_1_10((cvt_5_IntSaturation_17U_8U_if_acc_1_nl));
  assign cvt_5_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_1_nl
      = (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_5_sva[25]) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_5_sva))
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_5_sva;
  assign nl_cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_nl = ({1'b1 , (cvt_5_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_1_nl)
      , (~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_5_sva[23:14]))}) + 12'b1;
  assign cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_nl = nl_cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11:0];
  assign cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1 = readslicef_12_1_11((cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_nl));
  assign FpFloatToInt_16U_5U_10U_internal_int_0_sva_mx0w0 = ~((~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_sva[0])
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_sva)) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_sva);
  assign cvt_16_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_4_nl
      = (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_sva[25]) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_sva))
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_sva;
  assign nl_cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_nl = ({1'b1 , (cvt_16_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_4_nl)
      , (~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_sva[23:14]))}) + 12'b1;
  assign cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_nl = nl_cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_nl[11:0];
  assign cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_itm_11_1 = readslicef_12_1_11((cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_nl));
  assign FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_mx0w0 = ~((~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_6_sva[0])
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_6_sva)) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_6_sva);
  assign cvt_6_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl
      = (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_6_sva[25]) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_6_sva))
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_6_sva;
  assign nl_cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_nl = ({1'b1 , (cvt_6_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl)
      , (~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_6_sva[23:14]))}) + 12'b1;
  assign cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_nl = nl_cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11:0];
  assign cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1 = readslicef_12_1_11((cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_nl));
  assign FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_mx0w0 = ~((~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_15_sva[0])
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_15_sva)) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_15_sva);
  assign nl_cvt_1_IntSaturation_17U_8U_if_acc_nl = conv_s2u_10_11({(~ IntShiftRightSat_49U_6U_17U_o_16_1_sva_3)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_2[14:6]))}) + 11'b1;
  assign cvt_1_IntSaturation_17U_8U_if_acc_nl = nl_cvt_1_IntSaturation_17U_8U_if_acc_nl[10:0];
  assign cvt_1_IntSaturation_17U_8U_if_acc_itm_10_1 = readslicef_11_1_10((cvt_1_IntSaturation_17U_8U_if_acc_nl));
  assign cvt_15_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_3_nl
      = (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_15_sva[25]) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_15_sva))
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_15_sva;
  assign nl_cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_nl = ({1'b1 , (cvt_15_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_3_nl)
      , (~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_15_sva[23:14]))}) + 12'b1;
  assign cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_nl = nl_cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11:0];
  assign cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1 = readslicef_12_1_11((cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_nl));
  assign IsNaN_5U_10U_land_15_lpi_1_dfm_mx0w0 = ~(IsNaN_5U_10U_nor_14_itm_2 | IsNaN_5U_10U_IsNaN_5U_10U_nand_14_itm_2);
  assign FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_mx0w0 = ~((~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_7_sva[0])
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_7_sva)) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_7_sva);
  assign cvt_7_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl
      = (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_7_sva[25]) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_7_sva))
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_7_sva;
  assign nl_cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_nl = ({1'b1 , (cvt_7_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl)
      , (~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_7_sva[23:14]))}) + 12'b1;
  assign cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_nl = nl_cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11:0];
  assign cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1 = readslicef_12_1_11((cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_nl));
  assign FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_mx0w0 = ~((~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_14_sva[0])
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_14_sva)) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_14_sva);
  assign cvt_14_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_3_nl
      = (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_14_sva[25]) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_14_sva))
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_14_sva;
  assign nl_cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_nl = ({1'b1 , (cvt_14_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_3_nl)
      , (~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_14_sva[23:14]))}) + 12'b1;
  assign cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_nl = nl_cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11:0];
  assign cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1 = readslicef_12_1_11((cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_nl));
  assign FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_mx0w0 = ~((~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_8_sva[0])
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_8_sva)) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_8_sva);
  assign cvt_8_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_3_nl
      = (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_8_sva[25]) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_8_sva))
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_8_sva;
  assign nl_cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_nl = ({1'b1 , (cvt_8_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_3_nl)
      , (~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_8_sva[23:14]))}) + 12'b1;
  assign cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_nl = nl_cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11:0];
  assign cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1 = readslicef_12_1_11((cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_nl));
  assign FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_mx0w0 = ~((~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_13_sva[0])
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_13_sva)) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_13_sva);
  assign cvt_13_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl
      = (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_13_sva[25]) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_13_sva))
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_13_sva;
  assign nl_cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_nl = ({1'b1 , (cvt_13_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl)
      , (~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_13_sva[23:14]))}) + 12'b1;
  assign cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_nl = nl_cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11:0];
  assign cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1 = readslicef_12_1_11((cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_nl));
  assign FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_mx0w0 = ~((~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_9_sva[0])
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_9_sva)) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_9_sva);
  assign nl_cvt_9_IntSaturation_17U_8U_if_acc_1_nl = conv_s2u_10_11({(~ IntShiftRightSat_49U_6U_17U_o_16_9_sva_3)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_2[14:6]))}) + 11'b1;
  assign cvt_9_IntSaturation_17U_8U_if_acc_1_nl = nl_cvt_9_IntSaturation_17U_8U_if_acc_1_nl[10:0];
  assign cvt_9_IntSaturation_17U_8U_if_acc_1_itm_10_1 = readslicef_11_1_10((cvt_9_IntSaturation_17U_8U_if_acc_1_nl));
  assign cvt_9_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_1_nl
      = (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_9_sva[25]) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_9_sva))
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_9_sva;
  assign nl_cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_nl = ({1'b1 , (cvt_9_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_1_nl)
      , (~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_9_sva[23:14]))}) + 12'b1;
  assign cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_nl = nl_cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_nl[11:0];
  assign cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1 = readslicef_12_1_11((cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_nl));
  assign FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_mx0w0 = ~((~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_12_sva[0])
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_12_sva)) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_12_sva);
  assign cvt_12_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_3_nl
      = (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_12_sva[25]) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_12_sva))
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_12_sva;
  assign nl_cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_nl = ({1'b1 , (cvt_12_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_3_nl)
      , (~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_12_sva[23:14]))}) + 12'b1;
  assign cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_nl = nl_cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_nl[11:0];
  assign cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1 = readslicef_12_1_11((cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_nl));
  assign FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_mx0w0 = ~((~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_10_sva[0])
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_10_sva)) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_10_sva);
  assign cvt_10_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl
      = (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_10_sva[25]) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_10_sva))
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_10_sva;
  assign nl_cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_nl = ({1'b1 , (cvt_10_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl)
      , (~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_10_sva[23:14]))}) + 12'b1;
  assign cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_nl = nl_cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11:0];
  assign cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1 = readslicef_12_1_11((cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_nl));
  assign FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_mx0w0 = ~((~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_11_sva[0])
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_11_sva)) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_11_sva);
  assign cvt_11_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl
      = (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_11_sva[25]) | IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_11_sva))
      | IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_11_sva;
  assign nl_cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_nl = ({1'b1 , (cvt_11_FpFloatToInt_16U_5U_10U_IntSignedShiftRight_12U_6U_26U_obits_fixed_or_2_nl)
      , (~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_11_sva[23:14]))}) + 12'b1;
  assign cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_nl = nl_cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_nl[11:0];
  assign cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1 = readslicef_12_1_11((cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_nl));
  assign cvt_else_nor_dfs_1_mx1 = MUX_s_1_2_2(cvt_else_nor_dfs, cvt_else_nor_dfs_2,
      or_dcpl_178);
  assign cvt_else_equal_tmp_4_mx1 = MUX_s_1_2_2(cvt_else_equal_tmp_1, cvt_else_equal_tmp_5,
      or_dcpl_178);
  assign cvt_else_equal_tmp_3_mx0 = MUX_s_1_2_2(cvt_else_equal_tmp, FpIntToFloat_17U_5U_10U_is_inf_2_lpi_1_dfm_6,
      or_dcpl_178);
  assign cvt_else_nor_dfs_3_mx1 = MUX_s_1_2_2(cvt_else_nor_dfs, cvt_else_nor_dfs_10,
      or_dcpl_181);
  assign cvt_else_equal_tmp_10_mx0 = MUX_s_1_2_2(cvt_else_equal_tmp_1, FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_7,
      or_dcpl_181);
  assign cvt_else_equal_tmp_9_mx1 = MUX_s_1_2_2(cvt_else_equal_tmp, cvt_else_equal_tmp_9,
      or_dcpl_181);
  assign cvt_else_nor_dfs_5_mx1 = MUX_s_1_2_2(cvt_else_nor_dfs, cvt_else_nor_dfs_10,
      or_dcpl_184);
  assign cvt_else_equal_tmp_16_mx1 = MUX_s_1_2_2(cvt_else_equal_tmp_1, cvt_else_equal_tmp_16,
      or_dcpl_184);
  assign cvt_else_equal_tmp_15_mx0 = MUX_s_1_2_2(cvt_else_equal_tmp, FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_7,
      or_dcpl_184);
  assign cvt_else_nor_dfs_7_mx1 = MUX_s_1_2_2(cvt_else_nor_dfs, cvt_else_nor_dfs_11,
      or_dcpl_188);
  assign cvt_else_equal_tmp_22_mx1 = MUX_s_1_2_2(cvt_else_equal_tmp_1, cvt_else_equal_tmp_34,
      or_dcpl_188);
  assign cvt_else_equal_tmp_21_mx1 = MUX_s_1_2_2(cvt_else_equal_tmp, cvt_else_equal_tmp_33,
      or_dcpl_188);
  assign cvt_else_nor_dfs_6_mx1 = MUX_s_1_2_2(cvt_else_nor_dfs_10, cvt_else_nor_dfs,
      mux_tmp_1899);
  assign cvt_else_equal_tmp_19_mx0 = MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_8,
      cvt_else_equal_tmp_1, mux_tmp_1899);
  assign cvt_else_equal_tmp_18_mx0 = MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_7,
      cvt_else_equal_tmp, mux_tmp_1899);
  assign cvt_else_nor_dfs_9_mx1 = MUX_s_1_2_2(cvt_else_nor_dfs, reg_cvt_else_nor_dfs_9_cse,
      or_dcpl_195);
  assign cvt_else_equal_tmp_28_mx1 = MUX_s_1_2_2(cvt_else_equal_tmp_1, cvt_else_equal_tmp_28,
      or_dcpl_195);
  assign cvt_else_equal_tmp_27_mx0 = MUX_s_1_2_2(cvt_else_equal_tmp, FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_7,
      or_dcpl_195);
  assign cvt_else_nor_dfs_11_mx1 = MUX_s_1_2_2(cvt_else_nor_dfs, cvt_else_nor_dfs_11,
      or_dcpl_197);
  assign cvt_else_equal_tmp_34_mx1 = MUX_s_1_2_2(cvt_else_equal_tmp_1, cvt_else_equal_tmp_34,
      or_dcpl_197);
  assign cvt_else_equal_tmp_33_mx1 = MUX_s_1_2_2(cvt_else_equal_tmp, cvt_else_equal_tmp_33,
      or_dcpl_197);
  assign cvt_else_nor_dfs_10_mx1 = MUX_s_1_2_2(cvt_else_nor_dfs_10, cvt_else_nor_dfs,
      mux_tmp_987);
  assign cvt_else_equal_tmp_31_mx0 = MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_8,
      cvt_else_equal_tmp_1, mux_tmp_987);
  assign cvt_else_equal_tmp_30_mx0 = MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_7,
      cvt_else_equal_tmp, mux_tmp_987);
  assign cvt_else_nor_dfs_13_mx1 = MUX_s_1_2_2(cvt_else_nor_dfs, cvt_else_nor_dfs_15,
      or_dcpl_197);
  assign cvt_else_equal_tmp_40_mx1 = MUX_s_1_2_2(cvt_else_equal_tmp_1, cvt_else_equal_tmp_46,
      or_dcpl_197);
  assign cvt_else_equal_tmp_39_mx1 = MUX_s_1_2_2(cvt_else_equal_tmp, cvt_else_equal_tmp_45,
      or_dcpl_197);
  assign cvt_else_nor_dfs_15_mx1 = MUX_s_1_2_2(cvt_else_nor_dfs, cvt_else_nor_dfs_15,
      or_dcpl_210);
  assign cvt_else_equal_tmp_46_mx1 = MUX_s_1_2_2(cvt_else_equal_tmp_1, cvt_else_equal_tmp_46,
      or_dcpl_210);
  assign cvt_else_equal_tmp_45_mx1 = MUX_s_1_2_2(cvt_else_equal_tmp, cvt_else_equal_tmp_45,
      or_dcpl_210);
  assign cvt_else_nor_dfs_14_mx1 = MUX_s_1_2_2(cvt_else_nor_dfs_15, cvt_else_nor_dfs,
      and_tmp_248);
  assign cvt_else_equal_tmp_43_mx0 = MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_9,
      cvt_else_equal_tmp_1, and_tmp_248);
  assign cvt_else_equal_tmp_42_mx0 = MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_8,
      cvt_else_equal_tmp, and_tmp_248);
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_13_nl = (IntShiftRightSat_49U_6U_17U_o_0_14_sva_4
      & (~ cvt_14_IntSaturation_17U_8U_else_if_acc_3_itm_10)) | cvt_14_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_3_svs_1;
  assign cvt_else_mux_56_nl = MUX_s_1_2_2(cvt_else_nor_dfs, cvt_else_nor_dfs_15,
      and_1059_cse);
  assign cvt_else_mux_62_nl = MUX_s_1_2_2(cvt_else_equal_tmp, cvt_else_equal_tmp_45,
      and_1059_cse);
  assign cvt_else_mux_59_nl = MUX_s_1_2_2(cvt_else_equal_tmp_1, cvt_else_equal_tmp_46,
      and_1059_cse);
  assign chn_odata_data_13_0_lpi_1_dfm_1_mx0w0 = MUX1HOT_s_1_3_2((FpIntToFloat_17U_5U_10U_o_mant_14_lpi_1_dfm_1[0]),
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm_4, (IntSaturation_17U_8U_IntSaturation_17U_8U_or_13_nl),
      {(cvt_else_mux_56_nl) , (cvt_else_mux_62_nl) , (cvt_else_mux_59_nl)});
  assign cvt_else_equal_tmp_37_mx0 = MUX_s_1_2_2(cvt_else_equal_tmp_1, FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_8,
      or_dcpl_195);
  assign cvt_else_equal_tmp_36_mx0 = MUX_s_1_2_2(cvt_else_equal_tmp, FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_7,
      or_dcpl_195);
  assign nl_cvt_4_FpMantRNE_17U_11U_else_acc_2_nl = (cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[15:6])
      + conv_u2u_1_10(FpMantRNE_17U_11U_else_carry_4_sva);
  assign cvt_4_FpMantRNE_17U_11U_else_acc_2_nl = nl_cvt_4_FpMantRNE_17U_11U_else_acc_2_nl[9:0];
  assign FpIntToFloat_17U_5U_10U_if_not_185_nl = ~ cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_10_itm_mx0w0 = MUX_v_10_2_2(10'b0000000000,
      (cvt_4_FpMantRNE_17U_11U_else_acc_2_nl), (FpIntToFloat_17U_5U_10U_if_not_185_nl));
  assign or_3872_nl = and_dcpl_954 | FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_3;
  assign FpMantRNE_17U_11U_else_mux_7_nl = MUX_s_1_2_2(cvt_4_FpMantRNE_17U_11U_else_and_2_tmp,
      cvt_4_FpMantRNE_17U_11U_else_and_2_svs, or_3872_nl);
  assign FpIntToFloat_17U_5U_10U_else_mux_10_nl = MUX_s_1_2_2(or_1659_cse_1, FpIntToFloat_17U_5U_10U_else_unequal_tmp_3,
      FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_3);
  assign FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_2_mx1w0 = ~(((~((~ cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4)
      & (FpMantRNE_17U_11U_else_mux_7_nl))) & (FpIntToFloat_17U_5U_10U_else_mux_10_nl))
      | cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2);
  assign nl_cvt_5_FpMantRNE_17U_11U_else_acc_1_nl = (cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[15:6])
      + conv_u2u_1_10(FpMantRNE_17U_11U_else_carry_5_sva);
  assign cvt_5_FpMantRNE_17U_11U_else_acc_1_nl = nl_cvt_5_FpMantRNE_17U_11U_else_acc_1_nl[9:0];
  assign FpIntToFloat_17U_5U_10U_if_not_188_nl = ~ cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_13_itm_mx0w0 = MUX_v_10_2_2(10'b0000000000,
      (cvt_5_FpMantRNE_17U_11U_else_acc_1_nl), (FpIntToFloat_17U_5U_10U_if_not_188_nl));
  assign nl_cvt_6_FpMantRNE_17U_11U_else_acc_2_nl = (cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[15:6])
      + conv_u2u_1_10(FpMantRNE_17U_11U_else_carry_6_sva);
  assign cvt_6_FpMantRNE_17U_11U_else_acc_2_nl = nl_cvt_6_FpMantRNE_17U_11U_else_acc_2_nl[9:0];
  assign FpIntToFloat_17U_5U_10U_if_not_191_nl = ~ cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_16_itm_mx0w0 = MUX_v_10_2_2(10'b0000000000,
      (cvt_6_FpMantRNE_17U_11U_else_acc_2_nl), (FpIntToFloat_17U_5U_10U_if_not_191_nl));
  assign or_3891_nl = and_dcpl_962 | FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_3;
  assign FpMantRNE_17U_11U_else_mux_11_nl = MUX_s_1_2_2(cvt_6_FpMantRNE_17U_11U_else_and_2_tmp,
      cvt_6_FpMantRNE_17U_11U_else_and_2_svs, or_3891_nl);
  assign FpIntToFloat_17U_5U_10U_else_mux_16_nl = MUX_s_1_2_2(or_1720_cse_1, FpIntToFloat_17U_5U_10U_else_unequal_tmp_5,
      FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_3);
  assign FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_2_mx1w0 = ~(((~((~ cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4)
      & (FpMantRNE_17U_11U_else_mux_11_nl))) & (FpIntToFloat_17U_5U_10U_else_mux_16_nl))
      | cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2);
  assign nl_cvt_7_FpMantRNE_17U_11U_else_acc_2_nl = (cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[15:6])
      + conv_u2u_1_10(FpMantRNE_17U_11U_else_carry_7_sva);
  assign cvt_7_FpMantRNE_17U_11U_else_acc_2_nl = nl_cvt_7_FpMantRNE_17U_11U_else_acc_2_nl[9:0];
  assign FpIntToFloat_17U_5U_10U_if_not_194_nl = ~ cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_19_itm_mx0w0 = MUX_v_10_2_2(10'b0000000000,
      (cvt_7_FpMantRNE_17U_11U_else_acc_2_nl), (FpIntToFloat_17U_5U_10U_if_not_194_nl));
  assign or_3900_nl = and_dcpl_966 | FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_3;
  assign FpMantRNE_17U_11U_else_mux_13_nl = MUX_s_1_2_2(cvt_7_FpMantRNE_17U_11U_else_and_2_tmp,
      cvt_7_FpMantRNE_17U_11U_else_and_2_svs, or_3900_nl);
  assign FpIntToFloat_17U_5U_10U_else_mux_19_nl = MUX_s_1_2_2(or_1752_cse_1, FpIntToFloat_17U_5U_10U_else_unequal_tmp_6,
      FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_3);
  assign FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_2_mx1w0 = ~(((~((~ cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4)
      & (FpMantRNE_17U_11U_else_mux_13_nl))) & (FpIntToFloat_17U_5U_10U_else_mux_19_nl))
      | cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2);
  assign nl_cvt_8_FpMantRNE_17U_11U_else_acc_3_nl = (cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[15:6])
      + conv_u2u_1_10(FpMantRNE_17U_11U_else_carry_8_sva);
  assign cvt_8_FpMantRNE_17U_11U_else_acc_3_nl = nl_cvt_8_FpMantRNE_17U_11U_else_acc_3_nl[9:0];
  assign FpIntToFloat_17U_5U_10U_if_not_197_nl = ~ cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_22_itm_mx0w0 = MUX_v_10_2_2(10'b0000000000,
      (cvt_8_FpMantRNE_17U_11U_else_acc_3_nl), (FpIntToFloat_17U_5U_10U_if_not_197_nl));
  assign or_3911_nl = and_dcpl_970 | FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_3;
  assign FpMantRNE_17U_11U_else_mux_15_nl = MUX_s_1_2_2(cvt_8_FpMantRNE_17U_11U_else_and_3_tmp,
      cvt_8_FpMantRNE_17U_11U_else_and_3_svs, or_3911_nl);
  assign FpIntToFloat_17U_5U_10U_else_mux_22_nl = MUX_s_1_2_2(or_1789_cse_1, FpIntToFloat_17U_5U_10U_else_unequal_tmp_7,
      FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_3);
  assign FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_2_mx1w0 = ~(((~((~ cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4)
      & (FpMantRNE_17U_11U_else_mux_15_nl))) & (FpIntToFloat_17U_5U_10U_else_mux_22_nl))
      | cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2);
  assign nl_cvt_10_FpMantRNE_17U_11U_else_acc_2_nl = (cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[15:6])
      + conv_u2u_1_10(FpMantRNE_17U_11U_else_carry_10_sva);
  assign cvt_10_FpMantRNE_17U_11U_else_acc_2_nl = nl_cvt_10_FpMantRNE_17U_11U_else_acc_2_nl[9:0];
  assign FpIntToFloat_17U_5U_10U_if_not_203_nl = ~ cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_28_itm_mx0w0 = MUX_v_10_2_2(10'b0000000000,
      (cvt_10_FpMantRNE_17U_11U_else_acc_2_nl), (FpIntToFloat_17U_5U_10U_if_not_203_nl));
  assign or_3932_nl = and_dcpl_978 | FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_3;
  assign FpMantRNE_17U_11U_else_mux_19_nl = MUX_s_1_2_2(cvt_10_FpMantRNE_17U_11U_else_and_2_tmp,
      cvt_10_FpMantRNE_17U_11U_else_and_2_svs, or_3932_nl);
  assign FpIntToFloat_17U_5U_10U_else_mux_28_nl = MUX_s_1_2_2(or_1851_cse_1, FpIntToFloat_17U_5U_10U_else_unequal_tmp_9,
      FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_3);
  assign FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_2_mx0w0 = ~(((~((~ cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4)
      & (FpMantRNE_17U_11U_else_mux_19_nl))) & (FpIntToFloat_17U_5U_10U_else_mux_28_nl))
      | cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2);
  assign nl_cvt_11_FpMantRNE_17U_11U_else_acc_2_nl = (cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[15:6])
      + conv_u2u_1_10(FpMantRNE_17U_11U_else_carry_11_sva);
  assign cvt_11_FpMantRNE_17U_11U_else_acc_2_nl = nl_cvt_11_FpMantRNE_17U_11U_else_acc_2_nl[9:0];
  assign FpIntToFloat_17U_5U_10U_if_not_206_nl = ~ cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_31_itm_mx0w0 = MUX_v_10_2_2(10'b0000000000,
      (cvt_11_FpMantRNE_17U_11U_else_acc_2_nl), (FpIntToFloat_17U_5U_10U_if_not_206_nl));
  assign or_3942_nl = and_dcpl_982 | FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_3;
  assign FpMantRNE_17U_11U_else_mux_21_nl = MUX_s_1_2_2(cvt_11_FpMantRNE_17U_11U_else_and_2_tmp,
      cvt_11_FpMantRNE_17U_11U_else_and_2_svs, or_3942_nl);
  assign FpIntToFloat_17U_5U_10U_else_mux_31_nl = MUX_s_1_2_2(or_1892_cse_1, FpIntToFloat_17U_5U_10U_else_unequal_tmp_10,
      FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_3);
  assign FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_2_mx1w0 = ~(((~((~ cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4)
      & (FpMantRNE_17U_11U_else_mux_21_nl))) & (FpIntToFloat_17U_5U_10U_else_mux_31_nl))
      | cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2);
  assign nl_cvt_12_FpMantRNE_17U_11U_else_acc_3_nl = (cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[15:6])
      + conv_u2u_1_10(FpMantRNE_17U_11U_else_carry_12_sva);
  assign cvt_12_FpMantRNE_17U_11U_else_acc_3_nl = nl_cvt_12_FpMantRNE_17U_11U_else_acc_3_nl[9:0];
  assign FpIntToFloat_17U_5U_10U_if_not_209_nl = ~ cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_34_itm_mx0w0 = MUX_v_10_2_2(10'b0000000000,
      (cvt_12_FpMantRNE_17U_11U_else_acc_3_nl), (FpIntToFloat_17U_5U_10U_if_not_209_nl));
  assign or_3953_nl = and_dcpl_987 | FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_3;
  assign FpMantRNE_17U_11U_else_mux_23_nl = MUX_s_1_2_2(cvt_12_FpMantRNE_17U_11U_else_and_3_tmp,
      cvt_12_FpMantRNE_17U_11U_else_and_3_svs, or_3953_nl);
  assign FpIntToFloat_17U_5U_10U_else_mux_34_nl = MUX_s_1_2_2(or_1925_cse_1, FpIntToFloat_17U_5U_10U_else_unequal_tmp_11,
      FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_3);
  assign FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_2_mx1w0 = ~(((~((~ cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4)
      & (FpMantRNE_17U_11U_else_mux_23_nl))) & (FpIntToFloat_17U_5U_10U_else_mux_34_nl))
      | cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2);
  assign nl_cvt_13_FpMantRNE_17U_11U_else_acc_2_nl = (cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[15:6])
      + conv_u2u_1_10(FpMantRNE_17U_11U_else_carry_13_sva);
  assign cvt_13_FpMantRNE_17U_11U_else_acc_2_nl = nl_cvt_13_FpMantRNE_17U_11U_else_acc_2_nl[9:0];
  assign FpIntToFloat_17U_5U_10U_if_not_212_nl = ~ cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_37_itm_mx0w0 = MUX_v_10_2_2(10'b0000000000,
      (cvt_13_FpMantRNE_17U_11U_else_acc_2_nl), (FpIntToFloat_17U_5U_10U_if_not_212_nl));
  assign or_3965_nl = and_dcpl_991 | FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_3;
  assign FpMantRNE_17U_11U_else_mux_25_nl = MUX_s_1_2_2(cvt_13_FpMantRNE_17U_11U_else_and_2_tmp,
      cvt_13_FpMantRNE_17U_11U_else_and_2_svs, or_3965_nl);
  assign FpIntToFloat_17U_5U_10U_else_mux_37_nl = MUX_s_1_2_2(or_5038_cse, FpIntToFloat_17U_5U_10U_else_unequal_tmp_12,
      FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_3);
  assign FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_2_mx0w0 = ~(((~((~ cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4)
      & (FpMantRNE_17U_11U_else_mux_25_nl))) & (FpIntToFloat_17U_5U_10U_else_mux_37_nl))
      | cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2);
  assign nl_cvt_14_FpMantRNE_17U_11U_else_acc_3_nl = (cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[15:6])
      + conv_u2u_1_10(FpMantRNE_17U_11U_else_carry_14_sva);
  assign cvt_14_FpMantRNE_17U_11U_else_acc_3_nl = nl_cvt_14_FpMantRNE_17U_11U_else_acc_3_nl[9:0];
  assign FpIntToFloat_17U_5U_10U_if_not_215_nl = ~ cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_40_itm_mx0w0 = MUX_v_10_2_2(10'b0000000000,
      (cvt_14_FpMantRNE_17U_11U_else_acc_3_nl), (FpIntToFloat_17U_5U_10U_if_not_215_nl));
  assign or_3977_nl = and_dcpl_995 | FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2;
  assign FpMantRNE_17U_11U_else_mux_27_nl = MUX_s_1_2_2(cvt_14_FpMantRNE_17U_11U_else_and_3_tmp,
      cvt_14_FpMantRNE_17U_11U_else_and_3_svs, or_3977_nl);
  assign FpIntToFloat_17U_5U_10U_else_mux_40_nl = MUX_s_1_2_2(or_5053_cse, FpIntToFloat_17U_5U_10U_else_unequal_tmp_13,
      FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2);
  assign FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2_mx0w0 = ~(((~((~ cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4)
      & (FpMantRNE_17U_11U_else_mux_27_nl))) & (FpIntToFloat_17U_5U_10U_else_mux_40_nl))
      | cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2);
  assign nl_cvt_15_FpMantRNE_17U_11U_else_acc_3_nl = (cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[15:6])
      + conv_u2u_1_10(FpMantRNE_17U_11U_else_carry_15_sva);
  assign cvt_15_FpMantRNE_17U_11U_else_acc_3_nl = nl_cvt_15_FpMantRNE_17U_11U_else_acc_3_nl[9:0];
  assign FpIntToFloat_17U_5U_10U_if_not_218_nl = ~ cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_43_itm_mx0w0 = MUX_v_10_2_2(10'b0000000000,
      (cvt_15_FpMantRNE_17U_11U_else_acc_3_nl), (FpIntToFloat_17U_5U_10U_if_not_218_nl));
  assign or_3989_nl = and_dcpl_999 | FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_3;
  assign FpMantRNE_17U_11U_else_mux_29_nl = MUX_s_1_2_2(cvt_15_FpMantRNE_17U_11U_else_and_3_tmp,
      cvt_15_FpMantRNE_17U_11U_else_and_3_svs, or_3989_nl);
  assign FpIntToFloat_17U_5U_10U_else_mux_43_nl = MUX_s_1_2_2(or_5069_cse, FpIntToFloat_17U_5U_10U_else_unequal_tmp_14,
      FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_3);
  assign FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_2_mx0w0 = ~(((~((~ cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4)
      & (FpMantRNE_17U_11U_else_mux_29_nl))) & (FpIntToFloat_17U_5U_10U_else_mux_43_nl))
      | cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2);
  assign nl_cvt_16_FpMantRNE_17U_11U_else_acc_4_nl = (cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_tmp[15:6])
      + conv_u2u_1_10(FpMantRNE_17U_11U_else_carry_sva);
  assign cvt_16_FpMantRNE_17U_11U_else_acc_4_nl = nl_cvt_16_FpMantRNE_17U_11U_else_acc_4_nl[9:0];
  assign FpIntToFloat_17U_5U_10U_if_not_221_nl = ~ cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_svs_2;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_46_itm_mx0w0 = MUX_v_10_2_2(10'b0000000000,
      (cvt_16_FpMantRNE_17U_11U_else_acc_4_nl), (FpIntToFloat_17U_5U_10U_if_not_221_nl));
  assign or_3999_nl = and_dcpl_1003 | FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_3;
  assign FpMantRNE_17U_11U_else_mux_31_nl = MUX_s_1_2_2(cvt_16_FpMantRNE_17U_11U_else_and_4_tmp,
      cvt_16_FpMantRNE_17U_11U_else_and_4_svs, or_3999_nl);
  assign FpIntToFloat_17U_5U_10U_else_mux_46_nl = MUX_s_1_2_2(or_5086_cse, FpIntToFloat_17U_5U_10U_else_unequal_tmp_15,
      FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_3);
  assign FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_2_mx0w0 = ~(((~((~ cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_8_tmp_4)
      & (FpMantRNE_17U_11U_else_mux_31_nl))) & (FpIntToFloat_17U_5U_10U_else_mux_46_nl))
      | cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_svs_2);
  assign cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp = ~(IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0
      | (IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_mx0w0!=15'b000000000000000) | IntShiftRightSat_49U_6U_17U_o_0_8_sva_mx0w0);
  assign cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp = ~(IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0
      | (IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_mx0w0!=15'b000000000000000) |
      IntShiftRightSat_49U_6U_17U_o_0_12_sva_mx0w0);
  assign cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp = ~(IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0
      | (IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_mx0w0!=15'b000000000000000) |
      IntShiftRightSat_49U_6U_17U_o_0_14_sva_mx0w0);
  assign cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp = ~(IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0
      | (IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_mx0w0!=15'b000000000000000) |
      IntShiftRightSat_49U_6U_17U_o_0_15_sva_mx0w0);
  assign cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_tmp = ~(IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0
      | (IntShiftRightSat_49U_6U_17U_o_15_1_sva_mx0w0!=15'b000000000000000) | IntShiftRightSat_49U_6U_17U_o_0_sva_mx0w0);
  assign cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp = ~(IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0
      | (IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_mx0w0!=15'b000000000000000) | IntShiftRightSat_49U_6U_17U_o_0_4_sva_mx0w0);
  assign cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp = ~(IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0
      | (IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_mx0w0!=15'b000000000000000) | IntShiftRightSat_49U_6U_17U_o_0_6_sva_mx0w0);
  assign cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp = ~(IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0
      | (IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_mx0w0!=15'b000000000000000) | IntShiftRightSat_49U_6U_17U_o_0_7_sva_mx0w0);
  assign cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp = ~(IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0
      | (IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_mx0w0!=15'b000000000000000) |
      IntShiftRightSat_49U_6U_17U_o_0_10_sva_mx0w0);
  assign cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp = ~(IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0
      | (IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_mx0w0!=15'b000000000000000) |
      IntShiftRightSat_49U_6U_17U_o_0_11_sva_mx0w0);
  assign cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp = ~(IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0
      | (IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_mx0w0!=15'b000000000000000) |
      IntShiftRightSat_49U_6U_17U_o_0_13_sva_mx0w0);
  assign FpMantRNE_24U_11U_else_carry_1_sva_mx0w0 = (chn_in_rsci_d_mxwt[12]) & ((chn_in_rsci_d_mxwt[0])
      | (chn_in_rsci_d_mxwt[1]) | (chn_in_rsci_d_mxwt[2]) | (chn_in_rsci_d_mxwt[3])
      | (chn_in_rsci_d_mxwt[4]) | (chn_in_rsci_d_mxwt[5]) | (chn_in_rsci_d_mxwt[6])
      | (chn_in_rsci_d_mxwt[7]) | (chn_in_rsci_d_mxwt[8]) | (chn_in_rsci_d_mxwt[9])
      | (chn_in_rsci_d_mxwt[10]) | (chn_in_rsci_d_mxwt[11]) | (chn_in_rsci_d_mxwt[13]));
  assign FpMantRNE_24U_11U_else_carry_2_sva_mx0w0 = (chn_in_rsci_d_mxwt[44]) & ((chn_in_rsci_d_mxwt[32])
      | (chn_in_rsci_d_mxwt[33]) | (chn_in_rsci_d_mxwt[34]) | (chn_in_rsci_d_mxwt[35])
      | (chn_in_rsci_d_mxwt[36]) | (chn_in_rsci_d_mxwt[37]) | (chn_in_rsci_d_mxwt[38])
      | (chn_in_rsci_d_mxwt[39]) | (chn_in_rsci_d_mxwt[40]) | (chn_in_rsci_d_mxwt[41])
      | (chn_in_rsci_d_mxwt[42]) | (chn_in_rsci_d_mxwt[43]) | (chn_in_rsci_d_mxwt[45]));
  assign FpMantRNE_24U_11U_else_carry_3_sva_mx0w0 = (chn_in_rsci_d_mxwt[76]) & ((chn_in_rsci_d_mxwt[64])
      | (chn_in_rsci_d_mxwt[65]) | (chn_in_rsci_d_mxwt[66]) | (chn_in_rsci_d_mxwt[67])
      | (chn_in_rsci_d_mxwt[68]) | (chn_in_rsci_d_mxwt[69]) | (chn_in_rsci_d_mxwt[70])
      | (chn_in_rsci_d_mxwt[71]) | (chn_in_rsci_d_mxwt[72]) | (chn_in_rsci_d_mxwt[73])
      | (chn_in_rsci_d_mxwt[74]) | (chn_in_rsci_d_mxwt[75]) | (chn_in_rsci_d_mxwt[77]));
  assign FpMantRNE_24U_11U_else_carry_4_sva_mx0w0 = (chn_in_rsci_d_mxwt[108]) & ((chn_in_rsci_d_mxwt[96])
      | (chn_in_rsci_d_mxwt[97]) | (chn_in_rsci_d_mxwt[98]) | (chn_in_rsci_d_mxwt[99])
      | (chn_in_rsci_d_mxwt[100]) | (chn_in_rsci_d_mxwt[101]) | (chn_in_rsci_d_mxwt[102])
      | (chn_in_rsci_d_mxwt[103]) | (chn_in_rsci_d_mxwt[104]) | (chn_in_rsci_d_mxwt[105])
      | (chn_in_rsci_d_mxwt[106]) | (chn_in_rsci_d_mxwt[107]) | (chn_in_rsci_d_mxwt[109]));
  assign FpMantRNE_24U_11U_else_carry_5_sva_mx0w0 = (chn_in_rsci_d_mxwt[140]) & ((chn_in_rsci_d_mxwt[128])
      | (chn_in_rsci_d_mxwt[129]) | (chn_in_rsci_d_mxwt[130]) | (chn_in_rsci_d_mxwt[131])
      | (chn_in_rsci_d_mxwt[132]) | (chn_in_rsci_d_mxwt[133]) | (chn_in_rsci_d_mxwt[134])
      | (chn_in_rsci_d_mxwt[135]) | (chn_in_rsci_d_mxwt[136]) | (chn_in_rsci_d_mxwt[137])
      | (chn_in_rsci_d_mxwt[138]) | (chn_in_rsci_d_mxwt[139]) | (chn_in_rsci_d_mxwt[141]));
  assign FpMantRNE_24U_11U_else_carry_6_sva_mx0w0 = (chn_in_rsci_d_mxwt[172]) & ((chn_in_rsci_d_mxwt[160])
      | (chn_in_rsci_d_mxwt[161]) | (chn_in_rsci_d_mxwt[162]) | (chn_in_rsci_d_mxwt[163])
      | (chn_in_rsci_d_mxwt[164]) | (chn_in_rsci_d_mxwt[165]) | (chn_in_rsci_d_mxwt[166])
      | (chn_in_rsci_d_mxwt[167]) | (chn_in_rsci_d_mxwt[168]) | (chn_in_rsci_d_mxwt[169])
      | (chn_in_rsci_d_mxwt[170]) | (chn_in_rsci_d_mxwt[171]) | (chn_in_rsci_d_mxwt[173]));
  assign FpMantRNE_24U_11U_else_carry_7_sva_mx0w0 = (chn_in_rsci_d_mxwt[204]) & ((chn_in_rsci_d_mxwt[192])
      | (chn_in_rsci_d_mxwt[193]) | (chn_in_rsci_d_mxwt[194]) | (chn_in_rsci_d_mxwt[195])
      | (chn_in_rsci_d_mxwt[196]) | (chn_in_rsci_d_mxwt[197]) | (chn_in_rsci_d_mxwt[198])
      | (chn_in_rsci_d_mxwt[199]) | (chn_in_rsci_d_mxwt[200]) | (chn_in_rsci_d_mxwt[201])
      | (chn_in_rsci_d_mxwt[202]) | (chn_in_rsci_d_mxwt[203]) | (chn_in_rsci_d_mxwt[205]));
  assign FpMantRNE_24U_11U_else_carry_8_sva_mx0w0 = (chn_in_rsci_d_mxwt[236]) & ((chn_in_rsci_d_mxwt[224])
      | (chn_in_rsci_d_mxwt[225]) | (chn_in_rsci_d_mxwt[226]) | (chn_in_rsci_d_mxwt[227])
      | (chn_in_rsci_d_mxwt[228]) | (chn_in_rsci_d_mxwt[229]) | (chn_in_rsci_d_mxwt[230])
      | (chn_in_rsci_d_mxwt[231]) | (chn_in_rsci_d_mxwt[232]) | (chn_in_rsci_d_mxwt[233])
      | (chn_in_rsci_d_mxwt[234]) | (chn_in_rsci_d_mxwt[235]) | (chn_in_rsci_d_mxwt[237]));
  assign FpMantRNE_24U_11U_else_carry_9_sva_mx0w0 = (chn_in_rsci_d_mxwt[268]) & ((chn_in_rsci_d_mxwt[256])
      | (chn_in_rsci_d_mxwt[257]) | (chn_in_rsci_d_mxwt[258]) | (chn_in_rsci_d_mxwt[259])
      | (chn_in_rsci_d_mxwt[260]) | (chn_in_rsci_d_mxwt[261]) | (chn_in_rsci_d_mxwt[262])
      | (chn_in_rsci_d_mxwt[263]) | (chn_in_rsci_d_mxwt[264]) | (chn_in_rsci_d_mxwt[265])
      | (chn_in_rsci_d_mxwt[266]) | (chn_in_rsci_d_mxwt[267]) | (chn_in_rsci_d_mxwt[269]));
  assign FpMantRNE_24U_11U_else_carry_10_sva_mx0w0 = (chn_in_rsci_d_mxwt[300]) &
      ((chn_in_rsci_d_mxwt[288]) | (chn_in_rsci_d_mxwt[289]) | (chn_in_rsci_d_mxwt[290])
      | (chn_in_rsci_d_mxwt[291]) | (chn_in_rsci_d_mxwt[292]) | (chn_in_rsci_d_mxwt[293])
      | (chn_in_rsci_d_mxwt[294]) | (chn_in_rsci_d_mxwt[295]) | (chn_in_rsci_d_mxwt[296])
      | (chn_in_rsci_d_mxwt[297]) | (chn_in_rsci_d_mxwt[298]) | (chn_in_rsci_d_mxwt[299])
      | (chn_in_rsci_d_mxwt[301]));
  assign FpMantRNE_24U_11U_else_carry_11_sva_mx0w0 = (chn_in_rsci_d_mxwt[332]) &
      ((chn_in_rsci_d_mxwt[320]) | (chn_in_rsci_d_mxwt[321]) | (chn_in_rsci_d_mxwt[322])
      | (chn_in_rsci_d_mxwt[323]) | (chn_in_rsci_d_mxwt[324]) | (chn_in_rsci_d_mxwt[325])
      | (chn_in_rsci_d_mxwt[326]) | (chn_in_rsci_d_mxwt[327]) | (chn_in_rsci_d_mxwt[328])
      | (chn_in_rsci_d_mxwt[329]) | (chn_in_rsci_d_mxwt[330]) | (chn_in_rsci_d_mxwt[331])
      | (chn_in_rsci_d_mxwt[333]));
  assign FpMantRNE_24U_11U_else_carry_12_sva_mx0w0 = (chn_in_rsci_d_mxwt[364]) &
      ((chn_in_rsci_d_mxwt[352]) | (chn_in_rsci_d_mxwt[353]) | (chn_in_rsci_d_mxwt[354])
      | (chn_in_rsci_d_mxwt[355]) | (chn_in_rsci_d_mxwt[356]) | (chn_in_rsci_d_mxwt[357])
      | (chn_in_rsci_d_mxwt[358]) | (chn_in_rsci_d_mxwt[359]) | (chn_in_rsci_d_mxwt[360])
      | (chn_in_rsci_d_mxwt[361]) | (chn_in_rsci_d_mxwt[362]) | (chn_in_rsci_d_mxwt[363])
      | (chn_in_rsci_d_mxwt[365]));
  assign FpMantRNE_24U_11U_else_carry_13_sva_mx0w0 = (chn_in_rsci_d_mxwt[396]) &
      ((chn_in_rsci_d_mxwt[384]) | (chn_in_rsci_d_mxwt[385]) | (chn_in_rsci_d_mxwt[386])
      | (chn_in_rsci_d_mxwt[387]) | (chn_in_rsci_d_mxwt[388]) | (chn_in_rsci_d_mxwt[389])
      | (chn_in_rsci_d_mxwt[390]) | (chn_in_rsci_d_mxwt[391]) | (chn_in_rsci_d_mxwt[392])
      | (chn_in_rsci_d_mxwt[393]) | (chn_in_rsci_d_mxwt[394]) | (chn_in_rsci_d_mxwt[395])
      | (chn_in_rsci_d_mxwt[397]));
  assign FpMantRNE_24U_11U_else_carry_14_sva_mx0w0 = (chn_in_rsci_d_mxwt[428]) &
      ((chn_in_rsci_d_mxwt[416]) | (chn_in_rsci_d_mxwt[417]) | (chn_in_rsci_d_mxwt[418])
      | (chn_in_rsci_d_mxwt[419]) | (chn_in_rsci_d_mxwt[420]) | (chn_in_rsci_d_mxwt[421])
      | (chn_in_rsci_d_mxwt[422]) | (chn_in_rsci_d_mxwt[423]) | (chn_in_rsci_d_mxwt[424])
      | (chn_in_rsci_d_mxwt[425]) | (chn_in_rsci_d_mxwt[426]) | (chn_in_rsci_d_mxwt[427])
      | (chn_in_rsci_d_mxwt[429]));
  assign FpMantRNE_24U_11U_else_carry_15_sva_mx0w0 = (chn_in_rsci_d_mxwt[460]) &
      ((chn_in_rsci_d_mxwt[448]) | (chn_in_rsci_d_mxwt[449]) | (chn_in_rsci_d_mxwt[450])
      | (chn_in_rsci_d_mxwt[451]) | (chn_in_rsci_d_mxwt[452]) | (chn_in_rsci_d_mxwt[453])
      | (chn_in_rsci_d_mxwt[454]) | (chn_in_rsci_d_mxwt[455]) | (chn_in_rsci_d_mxwt[456])
      | (chn_in_rsci_d_mxwt[457]) | (chn_in_rsci_d_mxwt[458]) | (chn_in_rsci_d_mxwt[459])
      | (chn_in_rsci_d_mxwt[461]));
  assign FpMantRNE_24U_11U_else_carry_sva_mx0w0 = (chn_in_rsci_d_mxwt[492]) & ((chn_in_rsci_d_mxwt[480])
      | (chn_in_rsci_d_mxwt[481]) | (chn_in_rsci_d_mxwt[482]) | (chn_in_rsci_d_mxwt[483])
      | (chn_in_rsci_d_mxwt[484]) | (chn_in_rsci_d_mxwt[485]) | (chn_in_rsci_d_mxwt[486])
      | (chn_in_rsci_d_mxwt[487]) | (chn_in_rsci_d_mxwt[488]) | (chn_in_rsci_d_mxwt[489])
      | (chn_in_rsci_d_mxwt[490]) | (chn_in_rsci_d_mxwt[491]) | (chn_in_rsci_d_mxwt[493]));
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_15_tmp = ~((~((chn_in_rsci_d_mxwt[502:480]!=23'b00000000000000000000000)))
      | (chn_in_rsci_d_mxwt[510:503]!=8'b11111111));
  assign nl_cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_4_tmp = ({(~
      (chn_in_rsci_d_mxwt[507])) , (chn_in_rsci_d_mxwt[506:503])}) + 5'b1;
  assign cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_4_tmp = nl_cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_4_tmp[4:0];
  assign cvt_16_FpMantRNE_24U_11U_else_and_4_tmp = FpMantRNE_24U_11U_else_carry_sva_mx0w0
      & (chn_in_rsci_d_mxwt[502:493]==10'b1111111111);
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_14_tmp = ~((~((chn_in_rsci_d_mxwt[470:448]!=23'b00000000000000000000000)))
      | (chn_in_rsci_d_mxwt[478:471]!=8'b11111111));
  assign nl_cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp = ({(~
      (chn_in_rsci_d_mxwt[475])) , (chn_in_rsci_d_mxwt[474:471])}) + 5'b1;
  assign cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp = nl_cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp[4:0];
  assign cvt_15_FpMantRNE_24U_11U_else_and_3_tmp = FpMantRNE_24U_11U_else_carry_15_sva_mx0w0
      & (chn_in_rsci_d_mxwt[470:461]==10'b1111111111);
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_13_tmp = ~((~((chn_in_rsci_d_mxwt[438:416]!=23'b00000000000000000000000)))
      | (chn_in_rsci_d_mxwt[446:439]!=8'b11111111));
  assign nl_cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp = ({(~
      (chn_in_rsci_d_mxwt[443])) , (chn_in_rsci_d_mxwt[442:439])}) + 5'b1;
  assign cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp = nl_cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp[4:0];
  assign cvt_14_FpMantRNE_24U_11U_else_and_3_tmp = FpMantRNE_24U_11U_else_carry_14_sva_mx0w0
      & (chn_in_rsci_d_mxwt[438:429]==10'b1111111111);
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_12_tmp = ~((~((chn_in_rsci_d_mxwt[406:384]!=23'b00000000000000000000000)))
      | (chn_in_rsci_d_mxwt[414:407]!=8'b11111111));
  assign nl_cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp = ({(~
      (chn_in_rsci_d_mxwt[411])) , (chn_in_rsci_d_mxwt[410:407])}) + 5'b1;
  assign cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp = nl_cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp[4:0];
  assign cvt_13_FpMantRNE_24U_11U_else_and_2_tmp = FpMantRNE_24U_11U_else_carry_13_sva_mx0w0
      & (chn_in_rsci_d_mxwt[406:397]==10'b1111111111);
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_11_tmp = ~((~((chn_in_rsci_d_mxwt[374:352]!=23'b00000000000000000000000)))
      | (chn_in_rsci_d_mxwt[382:375]!=8'b11111111));
  assign nl_cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp = ({(~
      (chn_in_rsci_d_mxwt[379])) , (chn_in_rsci_d_mxwt[378:375])}) + 5'b1;
  assign cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp = nl_cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp[4:0];
  assign cvt_12_FpMantRNE_24U_11U_else_and_3_tmp = FpMantRNE_24U_11U_else_carry_12_sva_mx0w0
      & (chn_in_rsci_d_mxwt[374:365]==10'b1111111111);
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_10_tmp = ~((~((chn_in_rsci_d_mxwt[342:320]!=23'b00000000000000000000000)))
      | (chn_in_rsci_d_mxwt[350:343]!=8'b11111111));
  assign nl_cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp = ({(~
      (chn_in_rsci_d_mxwt[347])) , (chn_in_rsci_d_mxwt[346:343])}) + 5'b1;
  assign cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp = nl_cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp[4:0];
  assign cvt_11_FpMantRNE_24U_11U_else_and_2_tmp = FpMantRNE_24U_11U_else_carry_11_sva_mx0w0
      & (chn_in_rsci_d_mxwt[342:333]==10'b1111111111);
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_9_tmp = ~((~((chn_in_rsci_d_mxwt[310:288]!=23'b00000000000000000000000)))
      | (chn_in_rsci_d_mxwt[318:311]!=8'b11111111));
  assign nl_cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp = ({(~
      (chn_in_rsci_d_mxwt[315])) , (chn_in_rsci_d_mxwt[314:311])}) + 5'b1;
  assign cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp = nl_cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp[4:0];
  assign cvt_10_FpMantRNE_24U_11U_else_and_2_tmp = FpMantRNE_24U_11U_else_carry_10_sva_mx0w0
      & (chn_in_rsci_d_mxwt[310:301]==10'b1111111111);
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_8_tmp = ~((~((chn_in_rsci_d_mxwt[278:256]!=23'b00000000000000000000000)))
      | (chn_in_rsci_d_mxwt[286:279]!=8'b11111111));
  assign nl_cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp = ({(~
      (chn_in_rsci_d_mxwt[283])) , (chn_in_rsci_d_mxwt[282:279])}) + 5'b1;
  assign cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp = nl_cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp[4:0];
  assign cvt_9_FpMantRNE_24U_11U_else_and_1_tmp = FpMantRNE_24U_11U_else_carry_9_sva_mx0w0
      & (chn_in_rsci_d_mxwt[278:269]==10'b1111111111);
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_7_tmp = ~((~((chn_in_rsci_d_mxwt[246:224]!=23'b00000000000000000000000)))
      | (chn_in_rsci_d_mxwt[254:247]!=8'b11111111));
  assign nl_cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp = ({(~
      (chn_in_rsci_d_mxwt[251])) , (chn_in_rsci_d_mxwt[250:247])}) + 5'b1;
  assign cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp = nl_cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp[4:0];
  assign cvt_8_FpMantRNE_24U_11U_else_and_3_tmp = FpMantRNE_24U_11U_else_carry_8_sva_mx0w0
      & (chn_in_rsci_d_mxwt[246:237]==10'b1111111111);
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_6_tmp = ~((~((chn_in_rsci_d_mxwt[214:192]!=23'b00000000000000000000000)))
      | (chn_in_rsci_d_mxwt[222:215]!=8'b11111111));
  assign nl_cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp = ({(~
      (chn_in_rsci_d_mxwt[219])) , (chn_in_rsci_d_mxwt[218:215])}) + 5'b1;
  assign cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp = nl_cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp[4:0];
  assign cvt_7_FpMantRNE_24U_11U_else_and_2_tmp = FpMantRNE_24U_11U_else_carry_7_sva_mx0w0
      & (chn_in_rsci_d_mxwt[214:205]==10'b1111111111);
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_5_tmp = ~((~((chn_in_rsci_d_mxwt[182:160]!=23'b00000000000000000000000)))
      | (chn_in_rsci_d_mxwt[190:183]!=8'b11111111));
  assign nl_cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp = ({(~
      (chn_in_rsci_d_mxwt[187])) , (chn_in_rsci_d_mxwt[186:183])}) + 5'b1;
  assign cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp = nl_cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp[4:0];
  assign cvt_6_FpMantRNE_24U_11U_else_and_2_tmp = FpMantRNE_24U_11U_else_carry_6_sva_mx0w0
      & (chn_in_rsci_d_mxwt[182:173]==10'b1111111111);
  assign nl_cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp = ({(~
      (chn_in_rsci_d_mxwt[155])) , (chn_in_rsci_d_mxwt[154:151])}) + 5'b1;
  assign cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp = nl_cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp[4:0];
  assign cvt_5_FpMantRNE_24U_11U_else_and_1_tmp = FpMantRNE_24U_11U_else_carry_5_sva_mx0w0
      & (chn_in_rsci_d_mxwt[150:141]==10'b1111111111);
  assign IsNaN_8U_23U_nor_4_tmp = ~((chn_in_rsci_d_mxwt[150:128]!=23'b00000000000000000000000));
  assign IsNaN_8U_23U_IsNaN_8U_23U_nand_4_tmp = ~((chn_in_rsci_d_mxwt[158:151]==8'b11111111));
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_3_tmp = ~((~((chn_in_rsci_d_mxwt[118:96]!=23'b00000000000000000000000)))
      | (chn_in_rsci_d_mxwt[126:119]!=8'b11111111));
  assign nl_cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp = ({(~
      (chn_in_rsci_d_mxwt[123])) , (chn_in_rsci_d_mxwt[122:119])}) + 5'b1;
  assign cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp = nl_cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp[4:0];
  assign cvt_4_FpMantRNE_24U_11U_else_and_2_tmp = FpMantRNE_24U_11U_else_carry_4_sva_mx0w0
      & (chn_in_rsci_d_mxwt[118:109]==10'b1111111111);
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_2_tmp = ~((~((chn_in_rsci_d_mxwt[86:64]!=23'b00000000000000000000000)))
      | (chn_in_rsci_d_mxwt[94:87]!=8'b11111111));
  assign nl_cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp = ({(~
      (chn_in_rsci_d_mxwt[91])) , (chn_in_rsci_d_mxwt[90:87])}) + 5'b1;
  assign cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp = nl_cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp[4:0];
  assign cvt_3_FpMantRNE_24U_11U_else_and_1_tmp = FpMantRNE_24U_11U_else_carry_3_sva_mx0w0
      & (chn_in_rsci_d_mxwt[86:77]==10'b1111111111);
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_1_tmp = ~((~((chn_in_rsci_d_mxwt[54:32]!=23'b00000000000000000000000)))
      | (chn_in_rsci_d_mxwt[62:55]!=8'b11111111));
  assign nl_cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp = ({(~
      (chn_in_rsci_d_mxwt[59])) , (chn_in_rsci_d_mxwt[58:55])}) + 5'b1;
  assign cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp = nl_cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp[4:0];
  assign cvt_2_FpMantRNE_24U_11U_else_and_1_tmp = FpMantRNE_24U_11U_else_carry_2_sva_mx0w0
      & (chn_in_rsci_d_mxwt[54:45]==10'b1111111111);
  assign IsNaN_8U_23U_IsNaN_8U_23U_nor_tmp = ~((~((chn_in_rsci_d_mxwt[22:0]!=23'b00000000000000000000000)))
      | (chn_in_rsci_d_mxwt[30:23]!=8'b11111111));
  assign nl_cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_tmp = ({(~
      (chn_in_rsci_d_mxwt[27])) , (chn_in_rsci_d_mxwt[26:23])}) + 5'b1;
  assign cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_tmp = nl_cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_tmp[4:0];
  assign cvt_1_FpMantRNE_24U_11U_else_and_tmp = FpMantRNE_24U_11U_else_carry_1_sva_mx0w0
      & (chn_in_rsci_d_mxwt[22:13]==10'b1111111111);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_32_nl = MUX_s_1_2_2((~
      (chn_idata_data_sva_1_27_0_1[27])), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_sva_9[4]),
      cvt_1_FpMantRNE_24U_11U_else_and_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_7_4_mx0w0 = (~((~(((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_32_nl)
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_ssc))
      | nand_164_cse)) | FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_1_lpi_1_dfm)) | IsNaN_8U_23U_land_1_lpi_1_dfm_3;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_33_nl = MUX_s_1_2_2((~
      (chn_idata_data_sva_1_59_31_1[28])), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_sva_9[4]),
      cvt_2_FpMantRNE_24U_11U_else_and_1_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_7_4_mx0w0 = (~((~(((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_33_nl)
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_1_ssc))
      | nand_162_cse)) | FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_2_lpi_1_dfm)) | IsNaN_8U_23U_land_2_lpi_1_dfm_3;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_34_nl = MUX_s_1_2_2((~
      (chn_idata_data_sva_1_91_63_1[28])), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_sva_9[4]),
      cvt_3_FpMantRNE_24U_11U_else_and_1_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_7_4_mx0w0 = (~((~(((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_34_nl)
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_2_ssc))
      | nand_160_cse)) | FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_3_lpi_1_dfm)) | IsNaN_8U_23U_land_3_lpi_1_dfm_3;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_35_nl = MUX_s_1_2_2((~
      (chn_idata_data_sva_1_123_95_1[28])), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_sva_9[4]),
      cvt_4_FpMantRNE_24U_11U_else_and_2_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_7_4_mx0w0 = (~((~(((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_35_nl)
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_3_ssc))
      | nand_158_cse)) | FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_4_lpi_1_dfm)) | IsNaN_8U_23U_land_4_lpi_1_dfm_3;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_36_nl = MUX_s_1_2_2((~
      (chn_idata_data_sva_1_155_127_1[28])), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_sva_9[4]),
      cvt_5_FpMantRNE_24U_11U_else_and_1_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_7_4_mx0w0 = (~((~(((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_36_nl)
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_4_ssc))
      | nand_156_cse)) | FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_5_lpi_1_dfm)) | nor_1099_cse;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_37_nl = MUX_s_1_2_2((~
      (chn_idata_data_sva_1_187_159_1[28])), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_sva_9[4]),
      cvt_6_FpMantRNE_24U_11U_else_and_2_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_7_4_mx0w0 = (~((~(((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_37_nl)
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_5_ssc))
      | nand_153_cse)) | FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_6_lpi_1_dfm)) | IsNaN_8U_23U_land_6_lpi_1_dfm_3;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_38_nl = MUX_s_1_2_2((~
      (chn_idata_data_sva_1_219_191_1[28])), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_sva_9[4]),
      cvt_7_FpMantRNE_24U_11U_else_and_2_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_7_4_mx0w0 = (~((~(((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_38_nl)
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_6_ssc))
      | nand_151_cse)) | FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_7_lpi_1_dfm)) | IsNaN_8U_23U_land_7_lpi_1_dfm_3;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_39_nl = MUX_s_1_2_2((~
      (chn_idata_data_sva_1_251_223_1[28])), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_sva_9[4]),
      cvt_8_FpMantRNE_24U_11U_else_and_3_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_7_4_mx0w0 = (~((~(((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_39_nl)
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_7_ssc))
      | nand_149_cse)) | FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_8_lpi_1_dfm)) | IsNaN_8U_23U_land_8_lpi_1_dfm_3;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_40_nl = MUX_s_1_2_2((~
      (chn_idata_data_sva_1_283_255_1[28])), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_sva_9[4]),
      cvt_9_FpMantRNE_24U_11U_else_and_1_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_7_4_mx0w0 = (~((~(((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_40_nl)
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_8_ssc))
      | nand_147_cse)) | FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_9_lpi_1_dfm)) | IsNaN_8U_23U_land_9_lpi_1_dfm_3;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_41_nl = MUX_s_1_2_2((~
      (chn_idata_data_sva_1_315_287_1[28])), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_sva_9[4]),
      cvt_10_FpMantRNE_24U_11U_else_and_2_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_7_4_mx0w0 = (~((~(((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_41_nl)
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_9_ssc))
      | nand_145_cse)) | FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_10_lpi_1_dfm)) |
      IsNaN_8U_23U_land_10_lpi_1_dfm_3;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_42_nl = MUX_s_1_2_2((~
      (chn_idata_data_sva_1_347_319_1[28])), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_sva_9[4]),
      cvt_11_FpMantRNE_24U_11U_else_and_2_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_7_4_mx0w0 = (~((~(((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_42_nl)
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_10_ssc))
      | nand_143_cse)) | FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_11_lpi_1_dfm)) |
      IsNaN_8U_23U_land_11_lpi_1_dfm_3;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_43_nl = MUX_s_1_2_2((~
      (chn_idata_data_sva_1_379_351_1[28])), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_sva_9[4]),
      cvt_12_FpMantRNE_24U_11U_else_and_3_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_7_4_mx0w0 = (~((~(((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_43_nl)
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_11_ssc))
      | nand_141_cse)) | FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_12_lpi_1_dfm)) |
      IsNaN_8U_23U_land_12_lpi_1_dfm_3;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_44_nl = MUX_s_1_2_2((~
      (chn_idata_data_sva_1_411_383_1[28])), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_sva_9[4]),
      cvt_13_FpMantRNE_24U_11U_else_and_2_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_7_4_mx0w0 = (~((~(((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_44_nl)
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_12_ssc))
      | nand_139_cse)) | FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_13_lpi_1_dfm)) |
      IsNaN_8U_23U_land_13_lpi_1_dfm_3;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_45_nl = MUX_s_1_2_2((~
      (chn_idata_data_sva_1_443_415_1[28])), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_sva_9[4]),
      cvt_14_FpMantRNE_24U_11U_else_and_3_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_7_4_mx0w0 = (~((~(((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_45_nl)
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_13_ssc))
      | nand_137_cse)) | FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_14_lpi_1_dfm)) |
      IsNaN_8U_23U_land_14_lpi_1_dfm_3;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_46_nl = MUX_s_1_2_2((~
      (chn_idata_data_sva_1_475_447_1[28])), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_sva_9[4]),
      cvt_15_FpMantRNE_24U_11U_else_and_3_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_7_4_mx0w0 = (~((~(((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_46_nl)
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_14_ssc))
      | nand_135_cse)) | FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_15_lpi_1_dfm)) |
      IsNaN_8U_23U_land_15_lpi_1_dfm_3;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_47_nl = MUX_s_1_2_2((~
      (chn_idata_data_sva_1_507_479_1[28])), (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_sva_9[4]),
      cvt_16_FpMantRNE_24U_11U_else_and_4_svs_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_7_4_mx0w0 = (~((~(((FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_mux_47_nl)
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_15_ssc))
      | nand_133_cse)) | FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_lpi_1_dfm)) | IsNaN_8U_23U_land_lpi_1_dfm_3;
  assign IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm_mx0w0 = (IntShiftRightSat_49U_6U_17U_o_0_14_sva_mx0w0
      & (~ cvt_14_IntSaturation_17U_16U_else_if_acc_3_itm_2_1)) | cvt_14_IntSaturation_17U_16U_if_acc_3_itm_2_1;
  assign cvt_16_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_4_tmp
      = IntShiftRightSat_49U_6U_17U_i_sva_mx0w1 != conv_s2s_17_49({IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0
      , IntShiftRightSat_49U_6U_17U_o_15_1_sva_mx0w0 , IntShiftRightSat_49U_6U_17U_o_0_sva_mx0w0});
  assign cvt_13_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp
      = IntShiftRightSat_49U_6U_17U_i_13_sva_mx0w1 != conv_s2s_17_49({IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0
      , IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_mx0w0 , IntShiftRightSat_49U_6U_17U_o_0_13_sva_mx0w0});
  assign cvt_14_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp
      = IntShiftRightSat_49U_6U_17U_i_14_sva_mx0w1 != conv_s2s_17_49({IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0
      , IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_mx0w0 , IntShiftRightSat_49U_6U_17U_o_0_14_sva_mx0w0});
  assign cvt_15_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp
      = IntShiftRightSat_49U_6U_17U_i_15_sva_mx0w1 != conv_s2s_17_49({IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0
      , IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_mx0w0 , IntShiftRightSat_49U_6U_17U_o_0_15_sva_mx0w0});
  assign cvt_12_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp
      = IntShiftRightSat_49U_6U_17U_i_12_sva_mx0w1 != conv_s2s_17_49({IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0
      , IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_mx0w0 , IntShiftRightSat_49U_6U_17U_o_0_12_sva_mx0w0});
  assign nl_cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_2_sva_2
      , IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_2_sva_2})
      + 18'b1;
  assign cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl = nl_cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_lor_3_lpi_1_dfm_mx1w0 = ~((IntShiftRightSat_49U_6U_17U_i_2_sva_2
      != conv_s2s_18_49(cvt_2_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl)) & IntShiftRightSat_49U_6U_17U_lor_3_lpi_1_dfm);
  assign nl_cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_4_sva_2
      , IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_4_sva_2})
      + 18'b1;
  assign cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl = nl_cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_lor_5_lpi_1_dfm_mx1w0 = ~((IntShiftRightSat_49U_6U_17U_i_4_sva_2
      != conv_s2s_18_49(cvt_4_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl)) & IntShiftRightSat_49U_6U_17U_lor_5_lpi_1_dfm);
  assign nl_cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_3_sva_3
      , IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_3_sva_3})
      + 18'b1;
  assign cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl = nl_cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_lor_4_lpi_1_dfm_mx1w0 = ~((IntShiftRightSat_49U_6U_17U_i_3_sva_2
      != conv_s2s_18_49(cvt_3_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl)) & IntShiftRightSat_49U_6U_17U_lor_4_lpi_1_dfm);
  assign nl_cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_6_sva_2
      , IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_6_sva_2})
      + 18'b1;
  assign cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl = nl_cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_lor_7_lpi_1_dfm_mx1w0 = ~((IntShiftRightSat_49U_6U_17U_i_6_sva_2
      != conv_s2s_18_49(cvt_6_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl)) & IntShiftRightSat_49U_6U_17U_lor_7_lpi_1_dfm);
  assign nl_cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_8_sva_2
      , IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_8_sva_2})
      + 18'b1;
  assign cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl = nl_cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_lor_9_lpi_1_dfm_mx1w0 = ~((IntShiftRightSat_49U_6U_17U_i_8_sva_2
      != conv_s2s_18_49(cvt_8_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl)) & IntShiftRightSat_49U_6U_17U_lor_9_lpi_1_dfm);
  assign nl_cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_7_sva_2
      , IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_7_sva_2})
      + 18'b1;
  assign cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl = nl_cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_lor_8_lpi_1_dfm_mx1w0 = ~((IntShiftRightSat_49U_6U_17U_i_7_sva_2
      != conv_s2s_18_49(cvt_7_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl)) & IntShiftRightSat_49U_6U_17U_lor_8_lpi_1_dfm);
  assign nl_cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_5_sva_3
      , IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_5_sva_3})
      + 18'b1;
  assign cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl = nl_cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_lor_6_lpi_1_dfm_mx1w0 = ~((IntShiftRightSat_49U_6U_17U_i_5_sva_2
      != conv_s2s_18_49(cvt_5_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl)) & IntShiftRightSat_49U_6U_17U_lor_6_lpi_1_dfm);
  assign nl_cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_10_sva_2
      , IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_10_sva_2})
      + 18'b1;
  assign cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl = nl_cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_lor_11_lpi_1_dfm_mx1w0 = ~((IntShiftRightSat_49U_6U_17U_i_10_sva_2
      != conv_s2s_18_49(cvt_10_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl)) & IntShiftRightSat_49U_6U_17U_lor_10_lpi_1_dfm);
  assign cvt_10_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp
      = IntShiftRightSat_49U_6U_17U_i_10_sva_mx0w1 != conv_s2s_17_49({IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0
      , IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_mx0w0 , IntShiftRightSat_49U_6U_17U_o_0_10_sva_mx0w0});
  assign nl_cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_12_sva_2
      , IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_12_sva_2})
      + 18'b1;
  assign cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl = nl_cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_lor_13_lpi_1_dfm_mx1w0 = ~((IntShiftRightSat_49U_6U_17U_i_12_sva_2
      != conv_s2s_18_49(cvt_12_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl)) & IntShiftRightSat_49U_6U_17U_lor_13_lpi_1_dfm);
  assign nl_cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_11_sva_2
      , IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_11_sva_2})
      + 18'b1;
  assign cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl = nl_cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_lor_12_lpi_1_dfm_mx1w0 = ~((IntShiftRightSat_49U_6U_17U_i_11_sva_2
      != conv_s2s_18_49(cvt_11_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl)) & IntShiftRightSat_49U_6U_17U_lor_12_lpi_1_dfm);
  assign cvt_11_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp
      = IntShiftRightSat_49U_6U_17U_i_11_sva_mx0w1 != conv_s2s_17_49({IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0
      , IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_mx0w0 , IntShiftRightSat_49U_6U_17U_o_0_11_sva_mx0w0});
  assign nl_cvt_14_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_14_sva_2
      , IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_14_sva_3})
      + 18'b1;
  assign cvt_14_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl = nl_cvt_14_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_lor_15_lpi_1_dfm_mx1w0 = ~((IntShiftRightSat_49U_6U_17U_i_14_sva_2
      != conv_s2s_18_49(cvt_14_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl)) & IntShiftRightSat_49U_6U_17U_lor_15_lpi_1_dfm);
  assign nl_cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_sva_2
      , IntShiftRightSat_49U_6U_17U_o_15_1_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_sva_2})
      + 18'b1;
  assign cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl = nl_cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_lor_lpi_1_dfm_mx1w0 = ~((IntShiftRightSat_49U_6U_17U_i_sva_2
      != conv_s2s_18_49(cvt_16_IntShiftRightSat_49U_6U_17U_oif_acc_4_nl)) & IntShiftRightSat_49U_6U_17U_lor_lpi_1_dfm);
  assign nl_cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_15_sva_2
      , IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_15_sva_2})
      + 18'b1;
  assign cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl = nl_cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_lor_16_lpi_1_dfm_mx1w0 = ~((IntShiftRightSat_49U_6U_17U_i_15_sva_2
      != conv_s2s_18_49(cvt_15_IntShiftRightSat_49U_6U_17U_oif_acc_3_nl)) & IntShiftRightSat_49U_6U_17U_lor_16_lpi_1_dfm);
  assign nl_cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_13_sva_2
      , IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_13_sva_2})
      + 18'b1;
  assign cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl = nl_cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_lor_14_lpi_1_dfm_mx1w0 = ~((IntShiftRightSat_49U_6U_17U_i_13_sva_2
      != conv_s2s_18_49(cvt_13_IntShiftRightSat_49U_6U_17U_oif_acc_2_nl)) & IntShiftRightSat_49U_6U_17U_lor_14_lpi_1_dfm);
  assign nl_cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_9_sva_3
      , IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_9_sva_3})
      + 18'b1;
  assign cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl = nl_cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_lor_10_lpi_1_dfm_mx1w0 = ~((IntShiftRightSat_49U_6U_17U_i_9_sva_2
      != conv_s2s_18_49(cvt_9_IntShiftRightSat_49U_6U_17U_oif_acc_1_nl)) & cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_2);
  assign nl_cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_1_sva_3
      , IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_1_sva_2})
      + 18'b1;
  assign cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl = nl_cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_lor_2_lpi_1_dfm_mx1w0 = ~((IntShiftRightSat_49U_6U_17U_i_1_sva_2
      != conv_s2s_18_49(cvt_1_IntShiftRightSat_49U_6U_17U_oif_acc_nl)) & cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_svs_2);
  assign cvt_1_FpMantRNE_17U_11U_else_and_tmp = FpMantRNE_17U_11U_else_carry_1_sva
      & (FpIntToFloat_17U_5U_10U_else_int_mant_1_sva[16:6]==11'b11111111111);
  assign cvt_2_FpMantRNE_17U_11U_else_and_1_tmp = FpMantRNE_17U_11U_else_carry_2_sva
      & (FpIntToFloat_17U_5U_10U_else_int_mant_2_sva[16:6]==11'b11111111111);
  assign cvt_3_FpMantRNE_17U_11U_else_and_1_tmp = FpMantRNE_17U_11U_else_carry_3_sva
      & (cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[16:6]==11'b11111111111);
  assign cvt_4_FpMantRNE_17U_11U_else_and_2_tmp = FpMantRNE_17U_11U_else_carry_4_sva
      & (cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:6]==11'b11111111111);
  assign cvt_5_FpMantRNE_17U_11U_else_and_1_tmp = FpMantRNE_17U_11U_else_carry_5_sva
      & (cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[16:6]==11'b11111111111);
  assign cvt_6_FpMantRNE_17U_11U_else_and_2_tmp = FpMantRNE_17U_11U_else_carry_6_sva
      & (cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:6]==11'b11111111111);
  assign cvt_7_FpMantRNE_17U_11U_else_and_2_tmp = FpMantRNE_17U_11U_else_carry_7_sva
      & (cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:6]==11'b11111111111);
  assign cvt_8_FpMantRNE_17U_11U_else_and_3_tmp = FpMantRNE_17U_11U_else_carry_8_sva
      & (cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[16:6]==11'b11111111111);
  assign cvt_9_FpMantRNE_17U_11U_else_and_1_tmp = FpMantRNE_17U_11U_else_carry_9_sva
      & (FpIntToFloat_17U_5U_10U_else_int_mant_9_sva[16:6]==11'b11111111111);
  assign cvt_10_FpMantRNE_17U_11U_else_and_2_tmp = FpMantRNE_17U_11U_else_carry_10_sva
      & (cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:6]==11'b11111111111);
  assign cvt_11_FpMantRNE_17U_11U_else_and_2_tmp = FpMantRNE_17U_11U_else_carry_11_sva
      & (cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:6]==11'b11111111111);
  assign cvt_12_FpMantRNE_17U_11U_else_and_3_tmp = FpMantRNE_17U_11U_else_carry_12_sva
      & (cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[16:6]==11'b11111111111);
  assign cvt_13_FpMantRNE_17U_11U_else_and_2_tmp = FpMantRNE_17U_11U_else_carry_13_sva
      & (cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:6]==11'b11111111111);
  assign cvt_14_FpMantRNE_17U_11U_else_and_3_tmp = FpMantRNE_17U_11U_else_carry_14_sva
      & (cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[16:6]==11'b11111111111);
  assign cvt_15_FpMantRNE_17U_11U_else_and_3_tmp = FpMantRNE_17U_11U_else_carry_15_sva
      & (cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[16:6]==11'b11111111111);
  assign cvt_16_FpMantRNE_17U_11U_else_and_4_tmp = FpMantRNE_17U_11U_else_carry_sva
      & (cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_tmp[16:6]==11'b11111111111);
  assign nl_cvt_1_IntSaturation_17U_16U_if_acc_nl = conv_s2u_2_3({(~ IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_mx0w0[14]))}) + 3'b1;
  assign cvt_1_IntSaturation_17U_16U_if_acc_nl = nl_cvt_1_IntSaturation_17U_16U_if_acc_nl[2:0];
  assign cvt_1_IntSaturation_17U_16U_if_acc_itm_2_1 = readslicef_3_1_2((cvt_1_IntSaturation_17U_16U_if_acc_nl));
  assign nl_cvt_2_IntSaturation_17U_16U_if_acc_1_nl = conv_s2u_2_3({(~ IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_mx0w0[14]))}) + 3'b1;
  assign cvt_2_IntSaturation_17U_16U_if_acc_1_nl = nl_cvt_2_IntSaturation_17U_16U_if_acc_1_nl[2:0];
  assign cvt_2_IntSaturation_17U_16U_if_acc_1_itm_2_1 = readslicef_3_1_2((cvt_2_IntSaturation_17U_16U_if_acc_1_nl));
  assign cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_and_2_nl = (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[62])
      & ((IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[0]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[1])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[2]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[3])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[4]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[5])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[6]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[7])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[8]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[9])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[10]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[11])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[12]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[13])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[14]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[15])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[16]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[17])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[18]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[19])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[20]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[21])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[22]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[23])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[24]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[25])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[26]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[27])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[28]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[29])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[30]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[31])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[32]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[33])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[34]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[35])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[36]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[37])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[38]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[39])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[40]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[41])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[42]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[43])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[44]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[45])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[46]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[47])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[48]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[49])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[50]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[51])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[52]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[53])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[54]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[55])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[56]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[57])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[58]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[59])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[60]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[61])
      | (~ (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[111])));
  assign nl_cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp = conv_s2s_49_50(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_2_sva[111:63])
      + conv_u2s_1_50(cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_and_2_nl);
  assign cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp = nl_cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[49:0];
  assign cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp = (cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[49])
      & (~((cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[48:16]==33'b111111111111111111111111111111111)));
  assign cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp = ~((cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[49])
      | (~((cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[48:16]!=33'b000000000000000000000000000000000))));
  assign nl_cvt_3_IntSaturation_17U_16U_if_acc_1_nl = conv_s2u_2_3({(~ IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_mx0w0[14]))}) + 3'b1;
  assign cvt_3_IntSaturation_17U_16U_if_acc_1_nl = nl_cvt_3_IntSaturation_17U_16U_if_acc_1_nl[2:0];
  assign cvt_3_IntSaturation_17U_16U_if_acc_1_itm_2_1 = readslicef_3_1_2((cvt_3_IntSaturation_17U_16U_if_acc_1_nl));
  assign nl_cvt_4_IntSaturation_17U_16U_if_acc_2_nl = conv_s2u_2_3({(~ IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_mx0w0[14]))}) + 3'b1;
  assign cvt_4_IntSaturation_17U_16U_if_acc_2_nl = nl_cvt_4_IntSaturation_17U_16U_if_acc_2_nl[2:0];
  assign cvt_4_IntSaturation_17U_16U_if_acc_2_itm_2_1 = readslicef_3_1_2((cvt_4_IntSaturation_17U_16U_if_acc_2_nl));
  assign cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl = (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[62])
      & ((IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[0]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[1])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[2]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[3])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[4]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[5])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[6]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[7])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[8]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[9])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[10]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[11])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[12]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[13])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[14]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[15])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[16]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[17])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[18]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[19])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[20]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[21])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[22]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[23])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[24]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[25])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[26]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[27])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[28]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[29])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[30]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[31])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[32]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[33])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[34]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[35])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[36]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[37])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[38]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[39])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[40]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[41])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[42]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[43])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[44]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[45])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[46]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[47])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[48]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[49])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[50]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[51])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[52]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[53])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[54]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[55])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[56]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[57])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[58]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[59])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[60]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[61])
      | (~ (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[111])));
  assign nl_cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp = conv_s2s_49_50(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_4_sva[111:63])
      + conv_u2s_1_50(cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl);
  assign cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp = nl_cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49:0];
  assign cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp = (cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49])
      & (~((cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[48:16]==33'b111111111111111111111111111111111)));
  assign cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp = ~((cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49])
      | (~((cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[48:16]!=33'b000000000000000000000000000000000))));
  assign cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_and_2_nl = (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[62])
      & ((IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[0]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[1])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[2]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[3])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[4]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[5])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[6]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[7])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[8]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[9])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[10]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[11])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[12]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[13])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[14]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[15])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[16]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[17])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[18]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[19])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[20]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[21])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[22]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[23])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[24]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[25])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[26]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[27])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[28]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[29])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[30]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[31])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[32]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[33])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[34]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[35])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[36]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[37])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[38]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[39])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[40]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[41])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[42]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[43])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[44]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[45])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[46]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[47])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[48]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[49])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[50]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[51])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[52]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[53])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[54]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[55])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[56]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[57])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[58]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[59])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[60]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[61])
      | (~ (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[111])));
  assign nl_cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp = conv_s2s_49_50(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_3_sva[111:63])
      + conv_u2s_1_50(cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_and_2_nl);
  assign cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp = nl_cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[49:0];
  assign cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp = (cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[49])
      & (~((cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[48:16]==33'b111111111111111111111111111111111)));
  assign cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp = ~((cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[49])
      | (~((cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[48:16]!=33'b000000000000000000000000000000000))));
  assign nl_cvt_5_IntSaturation_17U_16U_if_acc_1_nl = conv_s2u_2_3({(~ IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_mx0w0[14]))}) + 3'b1;
  assign cvt_5_IntSaturation_17U_16U_if_acc_1_nl = nl_cvt_5_IntSaturation_17U_16U_if_acc_1_nl[2:0];
  assign cvt_5_IntSaturation_17U_16U_if_acc_1_itm_2_1 = readslicef_3_1_2((cvt_5_IntSaturation_17U_16U_if_acc_1_nl));
  assign nl_cvt_6_IntSaturation_17U_16U_if_acc_2_nl = conv_s2u_2_3({(~ IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_mx0w0[14]))}) + 3'b1;
  assign cvt_6_IntSaturation_17U_16U_if_acc_2_nl = nl_cvt_6_IntSaturation_17U_16U_if_acc_2_nl[2:0];
  assign cvt_6_IntSaturation_17U_16U_if_acc_2_itm_2_1 = readslicef_3_1_2((cvt_6_IntSaturation_17U_16U_if_acc_2_nl));
  assign cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl = (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[62])
      & ((IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[0]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[1])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[2]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[3])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[4]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[5])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[6]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[7])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[8]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[9])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[10]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[11])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[12]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[13])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[14]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[15])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[16]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[17])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[18]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[19])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[20]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[21])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[22]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[23])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[24]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[25])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[26]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[27])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[28]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[29])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[30]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[31])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[32]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[33])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[34]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[35])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[36]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[37])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[38]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[39])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[40]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[41])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[42]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[43])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[44]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[45])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[46]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[47])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[48]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[49])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[50]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[51])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[52]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[53])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[54]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[55])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[56]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[57])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[58]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[59])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[60]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[61])
      | (~ (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[111])));
  assign nl_cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp = conv_s2s_49_50(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_6_sva[111:63])
      + conv_u2s_1_50(cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl);
  assign cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp = nl_cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49:0];
  assign cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp = (cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49])
      & (~((cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[48:16]==33'b111111111111111111111111111111111)));
  assign cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp = ~((cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49])
      | (~((cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[48:16]!=33'b000000000000000000000000000000000))));
  assign nl_cvt_7_IntSaturation_17U_16U_if_acc_2_nl = conv_s2u_2_3({(~ IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_mx0w0[14]))}) + 3'b1;
  assign cvt_7_IntSaturation_17U_16U_if_acc_2_nl = nl_cvt_7_IntSaturation_17U_16U_if_acc_2_nl[2:0];
  assign cvt_7_IntSaturation_17U_16U_if_acc_2_itm_2_1 = readslicef_3_1_2((cvt_7_IntSaturation_17U_16U_if_acc_2_nl));
  assign nl_cvt_8_IntSaturation_17U_16U_if_acc_3_nl = conv_s2u_2_3({(~ IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_mx0w0[14]))}) + 3'b1;
  assign cvt_8_IntSaturation_17U_16U_if_acc_3_nl = nl_cvt_8_IntSaturation_17U_16U_if_acc_3_nl[2:0];
  assign cvt_8_IntSaturation_17U_16U_if_acc_3_itm_2_1 = readslicef_3_1_2((cvt_8_IntSaturation_17U_16U_if_acc_3_nl));
  assign cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_and_6_nl = (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[62])
      & ((IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[0]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[1])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[2]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[3])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[4]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[5])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[6]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[7])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[8]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[9])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[10]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[11])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[12]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[13])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[14]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[15])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[16]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[17])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[18]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[19])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[20]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[21])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[22]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[23])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[24]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[25])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[26]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[27])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[28]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[29])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[30]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[31])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[32]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[33])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[34]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[35])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[36]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[37])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[38]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[39])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[40]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[41])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[42]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[43])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[44]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[45])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[46]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[47])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[48]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[49])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[50]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[51])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[52]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[53])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[54]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[55])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[56]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[57])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[58]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[59])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[60]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[61])
      | (~ (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[111])));
  assign nl_cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp = conv_s2s_49_50(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_8_sva[111:63])
      + conv_u2s_1_50(cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_and_6_nl);
  assign cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp = nl_cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[49:0];
  assign cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp = (cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[49])
      & (~((cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[48:16]==33'b111111111111111111111111111111111)));
  assign cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp = ~((cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[49])
      | (~((cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[48:16]!=33'b000000000000000000000000000000000))));
  assign cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl = (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[62])
      & ((IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[0]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[1])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[2]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[3])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[4]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[5])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[6]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[7])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[8]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[9])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[10]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[11])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[12]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[13])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[14]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[15])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[16]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[17])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[18]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[19])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[20]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[21])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[22]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[23])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[24]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[25])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[26]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[27])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[28]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[29])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[30]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[31])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[32]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[33])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[34]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[35])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[36]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[37])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[38]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[39])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[40]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[41])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[42]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[43])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[44]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[45])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[46]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[47])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[48]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[49])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[50]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[51])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[52]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[53])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[54]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[55])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[56]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[57])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[58]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[59])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[60]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[61])
      | (~ (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[111])));
  assign nl_cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp = conv_s2s_49_50(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_7_sva[111:63])
      + conv_u2s_1_50(cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl);
  assign cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp = nl_cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49:0];
  assign cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp = (cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49])
      & (~((cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[48:16]==33'b111111111111111111111111111111111)));
  assign cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp = ~((cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49])
      | (~((cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[48:16]!=33'b000000000000000000000000000000000))));
  assign cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_and_2_nl = (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[62])
      & ((IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[0]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[1])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[2]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[3])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[4]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[5])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[6]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[7])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[8]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[9])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[10]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[11])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[12]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[13])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[14]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[15])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[16]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[17])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[18]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[19])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[20]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[21])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[22]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[23])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[24]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[25])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[26]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[27])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[28]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[29])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[30]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[31])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[32]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[33])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[34]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[35])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[36]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[37])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[38]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[39])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[40]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[41])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[42]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[43])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[44]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[45])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[46]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[47])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[48]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[49])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[50]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[51])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[52]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[53])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[54]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[55])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[56]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[57])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[58]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[59])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[60]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[61])
      | (~ (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[111])));
  assign nl_cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp = conv_s2s_49_50(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_5_sva[111:63])
      + conv_u2s_1_50(cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_and_2_nl);
  assign cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp = nl_cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[49:0];
  assign cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp = (cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[49])
      & (~((cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[48:16]==33'b111111111111111111111111111111111)));
  assign cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp = ~((cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[49])
      | (~((cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[48:16]!=33'b000000000000000000000000000000000))));
  assign nl_cvt_9_IntSaturation_17U_16U_if_acc_1_nl = conv_s2u_2_3({(~ IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_mx0w0[14]))}) + 3'b1;
  assign cvt_9_IntSaturation_17U_16U_if_acc_1_nl = nl_cvt_9_IntSaturation_17U_16U_if_acc_1_nl[2:0];
  assign cvt_9_IntSaturation_17U_16U_if_acc_1_itm_2_1 = readslicef_3_1_2((cvt_9_IntSaturation_17U_16U_if_acc_1_nl));
  assign nl_cvt_10_IntSaturation_17U_16U_if_acc_2_nl = conv_s2u_2_3({(~ IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_mx0w0[14]))}) + 3'b1;
  assign cvt_10_IntSaturation_17U_16U_if_acc_2_nl = nl_cvt_10_IntSaturation_17U_16U_if_acc_2_nl[2:0];
  assign cvt_10_IntSaturation_17U_16U_if_acc_2_itm_2_1 = readslicef_3_1_2((cvt_10_IntSaturation_17U_16U_if_acc_2_nl));
  assign cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl = (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[62])
      & ((IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[0]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[1])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[2]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[3])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[4]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[5])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[6]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[7])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[8]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[9])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[10]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[11])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[12]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[13])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[14]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[15])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[16]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[17])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[18]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[19])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[20]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[21])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[22]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[23])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[24]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[25])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[26]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[27])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[28]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[29])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[30]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[31])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[32]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[33])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[34]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[35])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[36]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[37])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[38]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[39])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[40]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[41])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[42]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[43])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[44]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[45])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[46]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[47])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[48]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[49])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[50]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[51])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[52]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[53])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[54]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[55])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[56]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[57])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[58]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[59])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[60]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[61])
      | (~ (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[111])));
  assign nl_cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp = conv_s2s_49_50(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_10_sva[111:63])
      + conv_u2s_1_50(cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl);
  assign cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp = nl_cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49:0];
  assign cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp = (cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49])
      & (~((cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[48:16]==33'b111111111111111111111111111111111)));
  assign cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp = ~((cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49])
      | (~((cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[48:16]!=33'b000000000000000000000000000000000))));
  assign nl_cvt_11_IntSaturation_17U_16U_if_acc_2_nl = conv_s2u_2_3({(~ IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_mx0w0[14]))}) + 3'b1;
  assign cvt_11_IntSaturation_17U_16U_if_acc_2_nl = nl_cvt_11_IntSaturation_17U_16U_if_acc_2_nl[2:0];
  assign cvt_11_IntSaturation_17U_16U_if_acc_2_itm_2_1 = readslicef_3_1_2((cvt_11_IntSaturation_17U_16U_if_acc_2_nl));
  assign nl_cvt_12_IntSaturation_17U_16U_if_acc_3_nl = conv_s2u_2_3({(~ IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_mx0w0[14]))}) + 3'b1;
  assign cvt_12_IntSaturation_17U_16U_if_acc_3_nl = nl_cvt_12_IntSaturation_17U_16U_if_acc_3_nl[2:0];
  assign cvt_12_IntSaturation_17U_16U_if_acc_3_itm_2_1 = readslicef_3_1_2((cvt_12_IntSaturation_17U_16U_if_acc_3_nl));
  assign cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_and_6_nl = (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[62])
      & ((IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[0]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[1])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[2]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[3])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[4]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[5])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[6]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[7])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[8]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[9])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[10]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[11])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[12]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[13])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[14]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[15])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[16]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[17])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[18]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[19])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[20]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[21])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[22]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[23])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[24]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[25])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[26]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[27])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[28]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[29])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[30]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[31])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[32]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[33])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[34]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[35])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[36]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[37])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[38]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[39])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[40]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[41])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[42]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[43])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[44]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[45])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[46]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[47])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[48]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[49])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[50]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[51])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[52]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[53])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[54]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[55])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[56]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[57])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[58]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[59])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[60]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[61])
      | (~ (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[111])));
  assign nl_cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp = conv_s2s_49_50(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_12_sva[111:63])
      + conv_u2s_1_50(cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_and_6_nl);
  assign cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp = nl_cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[49:0];
  assign cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp = (cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[49])
      & (~((cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[48:16]==33'b111111111111111111111111111111111)));
  assign cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp = ~((cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[49])
      | (~((cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[48:16]!=33'b000000000000000000000000000000000))));
  assign cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl = (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[62])
      & ((IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[0]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[1])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[2]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[3])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[4]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[5])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[6]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[7])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[8]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[9])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[10]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[11])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[12]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[13])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[14]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[15])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[16]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[17])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[18]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[19])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[20]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[21])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[22]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[23])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[24]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[25])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[26]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[27])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[28]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[29])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[30]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[31])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[32]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[33])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[34]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[35])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[36]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[37])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[38]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[39])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[40]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[41])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[42]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[43])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[44]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[45])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[46]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[47])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[48]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[49])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[50]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[51])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[52]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[53])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[54]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[55])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[56]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[57])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[58]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[59])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[60]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[61])
      | (~ (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[111])));
  assign nl_cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp = conv_s2s_49_50(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_11_sva[111:63])
      + conv_u2s_1_50(cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl);
  assign cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp = nl_cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49:0];
  assign cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp = (cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49])
      & (~((cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[48:16]==33'b111111111111111111111111111111111)));
  assign cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp = ~((cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49])
      | (~((cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[48:16]!=33'b000000000000000000000000000000000))));
  assign nl_cvt_13_IntSaturation_17U_16U_if_acc_2_nl = conv_s2u_2_3({(~ IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_mx0w0[14]))}) + 3'b1;
  assign cvt_13_IntSaturation_17U_16U_if_acc_2_nl = nl_cvt_13_IntSaturation_17U_16U_if_acc_2_nl[2:0];
  assign cvt_13_IntSaturation_17U_16U_if_acc_2_itm_2_1 = readslicef_3_1_2((cvt_13_IntSaturation_17U_16U_if_acc_2_nl));
  assign nl_cvt_14_IntSaturation_17U_16U_if_acc_3_nl = conv_s2u_2_3({(~ IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_mx0w0[14]))}) + 3'b1;
  assign cvt_14_IntSaturation_17U_16U_if_acc_3_nl = nl_cvt_14_IntSaturation_17U_16U_if_acc_3_nl[2:0];
  assign cvt_14_IntSaturation_17U_16U_if_acc_3_itm_2_1 = readslicef_3_1_2((cvt_14_IntSaturation_17U_16U_if_acc_3_nl));
  assign cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_and_6_nl = (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[62])
      & ((IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[0]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[1])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[2]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[3])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[4]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[5])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[6]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[7])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[8]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[9])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[10]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[11])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[12]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[13])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[14]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[15])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[16]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[17])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[18]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[19])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[20]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[21])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[22]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[23])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[24]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[25])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[26]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[27])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[28]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[29])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[30]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[31])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[32]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[33])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[34]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[35])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[36]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[37])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[38]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[39])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[40]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[41])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[42]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[43])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[44]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[45])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[46]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[47])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[48]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[49])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[50]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[51])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[52]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[53])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[54]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[55])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[56]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[57])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[58]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[59])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[60]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[61])
      | (~ (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[111])));
  assign nl_cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp = conv_s2s_49_50(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_14_sva[111:63])
      + conv_u2s_1_50(cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_and_6_nl);
  assign cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp = nl_cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[49:0];
  assign cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp = (cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[49])
      & (~((cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[48:16]==33'b111111111111111111111111111111111)));
  assign cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp = ~((cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[49])
      | (~((cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[48:16]!=33'b000000000000000000000000000000000))));
  assign nl_cvt_15_IntSaturation_17U_16U_if_acc_3_nl = conv_s2u_2_3({(~ IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_mx0w0[14]))}) + 3'b1;
  assign cvt_15_IntSaturation_17U_16U_if_acc_3_nl = nl_cvt_15_IntSaturation_17U_16U_if_acc_3_nl[2:0];
  assign cvt_15_IntSaturation_17U_16U_if_acc_3_itm_2_1 = readslicef_3_1_2((cvt_15_IntSaturation_17U_16U_if_acc_3_nl));
  assign nl_cvt_16_IntSaturation_17U_16U_if_acc_4_nl = conv_s2u_2_3({(~ IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_sva_mx0w0[14]))}) + 3'b1;
  assign cvt_16_IntSaturation_17U_16U_if_acc_4_nl = nl_cvt_16_IntSaturation_17U_16U_if_acc_4_nl[2:0];
  assign cvt_16_IntSaturation_17U_16U_if_acc_4_itm_2_1 = readslicef_3_1_2((cvt_16_IntSaturation_17U_16U_if_acc_4_nl));
  assign cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_and_8_nl = (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[62])
      & ((IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[0]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[1])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[2]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[3])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[4]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[5])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[6]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[7])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[8]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[9])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[10]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[11])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[12]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[13])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[14]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[15])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[16]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[17])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[18]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[19])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[20]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[21])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[22]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[23])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[24]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[25])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[26]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[27])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[28]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[29])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[30]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[31])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[32]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[33])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[34]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[35])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[36]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[37])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[38]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[39])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[40]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[41])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[42]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[43])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[44]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[45])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[46]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[47])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[48]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[49])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[50]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[51])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[52]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[53])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[54]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[55])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[56]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[57])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[58]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[59])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[60]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[61])
      | (~ (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[111])));
  assign nl_cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_acc_4_tmp = conv_s2s_49_50(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_sva[111:63])
      + conv_u2s_1_50(cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_and_8_nl);
  assign cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_acc_4_tmp = nl_cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_acc_4_tmp[49:0];
  assign cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_and_9_tmp = (cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_acc_4_tmp[49])
      & (~((cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_acc_4_tmp[48:16]==33'b111111111111111111111111111111111)));
  assign cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_nor_20_tmp = ~((cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_acc_4_tmp[49])
      | (~((cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_acc_4_tmp[48:16]!=33'b000000000000000000000000000000000))));
  assign cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_and_6_nl = (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[62])
      & ((IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[0]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[1])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[2]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[3])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[4]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[5])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[6]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[7])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[8]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[9])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[10]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[11])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[12]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[13])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[14]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[15])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[16]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[17])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[18]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[19])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[20]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[21])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[22]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[23])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[24]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[25])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[26]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[27])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[28]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[29])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[30]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[31])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[32]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[33])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[34]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[35])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[36]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[37])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[38]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[39])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[40]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[41])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[42]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[43])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[44]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[45])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[46]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[47])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[48]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[49])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[50]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[51])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[52]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[53])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[54]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[55])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[56]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[57])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[58]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[59])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[60]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[61])
      | (~ (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[111])));
  assign nl_cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp = conv_s2s_49_50(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_15_sva[111:63])
      + conv_u2s_1_50(cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_and_6_nl);
  assign cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp = nl_cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[49:0];
  assign cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp = (cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[49])
      & (~((cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[48:16]==33'b111111111111111111111111111111111)));
  assign cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp = ~((cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[49])
      | (~((cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[48:16]!=33'b000000000000000000000000000000000))));
  assign cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl = (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[62])
      & ((IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[0]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[1])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[2]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[3])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[4]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[5])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[6]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[7])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[8]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[9])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[10]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[11])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[12]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[13])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[14]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[15])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[16]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[17])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[18]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[19])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[20]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[21])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[22]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[23])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[24]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[25])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[26]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[27])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[28]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[29])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[30]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[31])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[32]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[33])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[34]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[35])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[36]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[37])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[38]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[39])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[40]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[41])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[42]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[43])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[44]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[45])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[46]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[47])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[48]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[49])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[50]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[51])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[52]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[53])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[54]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[55])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[56]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[57])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[58]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[59])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[60]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[61])
      | (~ (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[111])));
  assign nl_cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp = conv_s2s_49_50(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_13_sva[111:63])
      + conv_u2s_1_50(cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_and_4_nl);
  assign cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp = nl_cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49:0];
  assign cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp = (cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49])
      & (~((cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[48:16]==33'b111111111111111111111111111111111)));
  assign cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp = ~((cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[49])
      | (~((cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[48:16]!=33'b000000000000000000000000000000000))));
  assign cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_and_2_nl = (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[62])
      & ((IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[0]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[1])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[2]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[3])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[4]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[5])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[6]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[7])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[8]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[9])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[10]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[11])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[12]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[13])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[14]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[15])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[16]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[17])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[18]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[19])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[20]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[21])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[22]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[23])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[24]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[25])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[26]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[27])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[28]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[29])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[30]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[31])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[32]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[33])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[34]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[35])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[36]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[37])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[38]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[39])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[40]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[41])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[42]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[43])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[44]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[45])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[46]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[47])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[48]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[49])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[50]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[51])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[52]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[53])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[54]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[55])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[56]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[57])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[58]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[59])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[60]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[61])
      | (~ (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[111])));
  assign nl_cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp = conv_s2s_49_50(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_9_sva[111:63])
      + conv_u2s_1_50(cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_and_2_nl);
  assign cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp = nl_cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[49:0];
  assign cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp = (cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[49])
      & (~((cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[48:16]==33'b111111111111111111111111111111111)));
  assign cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp = ~((cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[49])
      | (~((cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[48:16]!=33'b000000000000000000000000000000000))));
  assign cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_and_nl = (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[62])
      & ((IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[0]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[1])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[2]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[3])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[4]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[5])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[6]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[7])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[8]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[9])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[10]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[11])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[12]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[13])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[14]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[15])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[16]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[17])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[18]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[19])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[20]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[21])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[22]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[23])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[24]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[25])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[26]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[27])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[28]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[29])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[30]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[31])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[32]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[33])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[34]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[35])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[36]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[37])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[38]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[39])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[40]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[41])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[42]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[43])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[44]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[45])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[46]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[47])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[48]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[49])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[50]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[51])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[52]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[53])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[54]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[55])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[56]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[57])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[58]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[59])
      | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[60]) | (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[61])
      | (~ (IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[111])));
  assign nl_cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_acc_tmp = conv_s2s_49_50(IntShiftRight_49U_6U_17U_obits_fixed_asn_rndi_1_sva[111:63])
      + conv_u2s_1_50(cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_and_nl);
  assign cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_acc_tmp = nl_cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_acc_tmp[49:0];
  assign cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_and_1_tmp = (cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_acc_tmp[49])
      & (~((cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_acc_tmp[48:16]==33'b111111111111111111111111111111111)));
  assign cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_nor_tmp = ~((cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_acc_tmp[49])
      | (~((cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_acc_tmp[48:16]!=33'b000000000000000000000000000000000))));
  assign cvt_1_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_nl = (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[30])
      & ((IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[0]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[1])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[2]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[3])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[4]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[5])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[6]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[7])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[8]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[9])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[10]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[11])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[12]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[13])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[14]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[15])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[16]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[17])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[18]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[19])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[20]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[21])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[22]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[23])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[24]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[25])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[26]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[27])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[28]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[29])
      | (~ (IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[74])));
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_1_sva = conv_s2s_44_45(IntSignedShiftRight_12U_6U_26U_mbits_fixed_1_sva[74:31])
      + conv_u2s_1_45(cvt_1_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_nl);
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_1_sva = nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_1_sva[44:0];
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_1_sva = (IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_1_sva[44])
      & (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_1_sva[43:25]==19'b1111111111111111111)));
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_1_sva = ~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_1_sva[44])
      | (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_1_sva[43:25]!=19'b0000000000000000000))));
  assign cvt_1_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_2_nl = ~(MUX_v_24_2_2((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_1_sva[24:1]),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_1_sva));
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_1_sva = ~(MUX_v_24_2_2((cvt_1_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_2_nl),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_1_sva));
  assign cvt_2_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_2_nl = (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[30])
      & ((IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[0]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[1])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[2]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[3])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[4]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[5])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[6]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[7])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[8]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[9])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[10]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[11])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[12]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[13])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[14]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[15])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[16]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[17])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[18]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[19])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[20]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[21])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[22]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[23])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[24]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[25])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[26]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[27])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[28]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[29])
      | (~ (IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[74])));
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_2_sva = conv_s2s_44_45(IntSignedShiftRight_12U_6U_26U_mbits_fixed_2_sva[74:31])
      + conv_u2s_1_45(cvt_2_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_2_nl);
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_2_sva = nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_2_sva[44:0];
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_2_sva = (IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_2_sva[44])
      & (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_2_sva[43:25]==19'b1111111111111111111)));
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_2_sva = ~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_2_sva[44])
      | (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_2_sva[43:25]!=19'b0000000000000000000))));
  assign cvt_2_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_7_nl = ~(MUX_v_24_2_2((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_2_sva[24:1]),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_2_sva));
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_2_sva = ~(MUX_v_24_2_2((cvt_2_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_7_nl),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_2_sva));
  assign cvt_3_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_2_nl = (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[30])
      & ((IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[0]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[1])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[2]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[3])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[4]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[5])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[6]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[7])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[8]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[9])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[10]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[11])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[12]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[13])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[14]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[15])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[16]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[17])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[18]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[19])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[20]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[21])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[22]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[23])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[24]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[25])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[26]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[27])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[28]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[29])
      | (~ (IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[74])));
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_3_sva = conv_s2s_44_45(IntSignedShiftRight_12U_6U_26U_mbits_fixed_3_sva[74:31])
      + conv_u2s_1_45(cvt_3_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_2_nl);
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_3_sva = nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_3_sva[44:0];
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_3_sva = (IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_3_sva[44])
      & (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_3_sva[43:25]==19'b1111111111111111111)));
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_3_sva = ~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_3_sva[44])
      | (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_3_sva[43:25]!=19'b0000000000000000000))));
  assign cvt_3_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_7_nl = ~(MUX_v_24_2_2((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_3_sva[24:1]),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_3_sva));
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_3_sva = ~(MUX_v_24_2_2((cvt_3_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_7_nl),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_3_sva));
  assign cvt_4_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl = (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[30])
      & ((IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[0]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[1])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[2]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[3])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[4]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[5])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[6]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[7])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[8]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[9])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[10]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[11])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[12]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[13])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[14]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[15])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[16]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[17])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[18]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[19])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[20]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[21])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[22]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[23])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[24]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[25])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[26]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[27])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[28]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[29])
      | (~ (IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[74])));
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_4_sva = conv_s2s_44_45(IntSignedShiftRight_12U_6U_26U_mbits_fixed_4_sva[74:31])
      + conv_u2s_1_45(cvt_4_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl);
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_4_sva = nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_4_sva[44:0];
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_4_sva = (IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_4_sva[44])
      & (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_4_sva[43:25]==19'b1111111111111111111)));
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_4_sva = ~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_4_sva[44])
      | (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_4_sva[43:25]!=19'b0000000000000000000))));
  assign cvt_4_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl = ~(MUX_v_24_2_2((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_4_sva[24:1]),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_4_sva));
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_4_sva = ~(MUX_v_24_2_2((cvt_4_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_4_sva));
  assign cvt_5_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_2_nl = (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[30])
      & ((IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[0]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[1])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[2]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[3])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[4]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[5])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[6]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[7])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[8]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[9])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[10]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[11])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[12]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[13])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[14]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[15])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[16]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[17])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[18]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[19])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[20]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[21])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[22]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[23])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[24]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[25])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[26]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[27])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[28]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[29])
      | (~ (IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[74])));
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_5_sva = conv_s2s_44_45(IntSignedShiftRight_12U_6U_26U_mbits_fixed_5_sva[74:31])
      + conv_u2s_1_45(cvt_5_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_2_nl);
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_5_sva = nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_5_sva[44:0];
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_5_sva = (IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_5_sva[44])
      & (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_5_sva[43:25]==19'b1111111111111111111)));
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_5_sva = ~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_5_sva[44])
      | (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_5_sva[43:25]!=19'b0000000000000000000))));
  assign cvt_5_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_7_nl = ~(MUX_v_24_2_2((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_5_sva[24:1]),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_5_sva));
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_5_sva = ~(MUX_v_24_2_2((cvt_5_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_7_nl),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_5_sva));
  assign cvt_6_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl = (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[30])
      & ((IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[0]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[1])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[2]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[3])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[4]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[5])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[6]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[7])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[8]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[9])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[10]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[11])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[12]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[13])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[14]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[15])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[16]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[17])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[18]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[19])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[20]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[21])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[22]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[23])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[24]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[25])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[26]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[27])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[28]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[29])
      | (~ (IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[74])));
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_6_sva = conv_s2s_44_45(IntSignedShiftRight_12U_6U_26U_mbits_fixed_6_sva[74:31])
      + conv_u2s_1_45(cvt_6_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl);
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_6_sva = nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_6_sva[44:0];
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_6_sva = (IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_6_sva[44])
      & (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_6_sva[43:25]==19'b1111111111111111111)));
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_6_sva = ~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_6_sva[44])
      | (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_6_sva[43:25]!=19'b0000000000000000000))));
  assign cvt_6_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl = ~(MUX_v_24_2_2((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_6_sva[24:1]),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_6_sva));
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_6_sva = ~(MUX_v_24_2_2((cvt_6_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_6_sva));
  assign cvt_7_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl = (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[30])
      & ((IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[0]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[1])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[2]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[3])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[4]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[5])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[6]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[7])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[8]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[9])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[10]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[11])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[12]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[13])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[14]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[15])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[16]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[17])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[18]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[19])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[20]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[21])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[22]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[23])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[24]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[25])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[26]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[27])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[28]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[29])
      | (~ (IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[74])));
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_7_sva = conv_s2s_44_45(IntSignedShiftRight_12U_6U_26U_mbits_fixed_7_sva[74:31])
      + conv_u2s_1_45(cvt_7_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl);
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_7_sva = nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_7_sva[44:0];
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_7_sva = (IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_7_sva[44])
      & (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_7_sva[43:25]==19'b1111111111111111111)));
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_7_sva = ~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_7_sva[44])
      | (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_7_sva[43:25]!=19'b0000000000000000000))));
  assign cvt_7_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl = ~(MUX_v_24_2_2((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_7_sva[24:1]),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_7_sva));
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_7_sva = ~(MUX_v_24_2_2((cvt_7_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_7_sva));
  assign cvt_8_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_6_nl = (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[30])
      & ((IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[0]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[1])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[2]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[3])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[4]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[5])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[6]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[7])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[8]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[9])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[10]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[11])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[12]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[13])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[14]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[15])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[16]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[17])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[18]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[19])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[20]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[21])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[22]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[23])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[24]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[25])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[26]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[27])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[28]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[29])
      | (~ (IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[74])));
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_8_sva = conv_s2s_44_45(IntSignedShiftRight_12U_6U_26U_mbits_fixed_8_sva[74:31])
      + conv_u2s_1_45(cvt_8_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_6_nl);
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_8_sva = nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_8_sva[44:0];
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_8_sva = (IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_8_sva[44])
      & (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_8_sva[43:25]==19'b1111111111111111111)));
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_8_sva = ~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_8_sva[44])
      | (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_8_sva[43:25]!=19'b0000000000000000000))));
  assign cvt_8_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_17_nl = ~(MUX_v_24_2_2((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_8_sva[24:1]),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_8_sva));
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_8_sva = ~(MUX_v_24_2_2((cvt_8_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_17_nl),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_8_sva));
  assign cvt_9_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_2_nl = (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[30])
      & ((IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[0]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[1])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[2]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[3])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[4]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[5])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[6]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[7])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[8]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[9])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[10]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[11])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[12]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[13])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[14]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[15])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[16]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[17])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[18]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[19])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[20]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[21])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[22]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[23])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[24]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[25])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[26]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[27])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[28]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[29])
      | (~ (IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[74])));
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_9_sva = conv_s2s_44_45(IntSignedShiftRight_12U_6U_26U_mbits_fixed_9_sva[74:31])
      + conv_u2s_1_45(cvt_9_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_2_nl);
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_9_sva = nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_9_sva[44:0];
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_9_sva = (IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_9_sva[44])
      & (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_9_sva[43:25]==19'b1111111111111111111)));
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_9_sva = ~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_9_sva[44])
      | (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_9_sva[43:25]!=19'b0000000000000000000))));
  assign cvt_9_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_7_nl = ~(MUX_v_24_2_2((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_9_sva[24:1]),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_9_sva));
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_9_sva = ~(MUX_v_24_2_2((cvt_9_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_7_nl),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_9_sva));
  assign cvt_10_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl = (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[30])
      & ((IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[0]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[1])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[2]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[3])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[4]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[5])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[6]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[7])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[8]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[9])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[10]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[11])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[12]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[13])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[14]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[15])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[16]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[17])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[18]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[19])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[20]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[21])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[22]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[23])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[24]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[25])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[26]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[27])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[28]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[29])
      | (~ (IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[74])));
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_10_sva = conv_s2s_44_45(IntSignedShiftRight_12U_6U_26U_mbits_fixed_10_sva[74:31])
      + conv_u2s_1_45(cvt_10_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl);
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_10_sva = nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_10_sva[44:0];
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_10_sva = (IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_10_sva[44])
      & (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_10_sva[43:25]==19'b1111111111111111111)));
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_10_sva = ~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_10_sva[44])
      | (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_10_sva[43:25]!=19'b0000000000000000000))));
  assign cvt_10_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl = ~(MUX_v_24_2_2((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_10_sva[24:1]),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_10_sva));
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_10_sva = ~(MUX_v_24_2_2((cvt_10_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_10_sva));
  assign cvt_11_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl = (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[30])
      & ((IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[0]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[1])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[2]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[3])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[4]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[5])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[6]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[7])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[8]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[9])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[10]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[11])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[12]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[13])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[14]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[15])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[16]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[17])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[18]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[19])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[20]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[21])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[22]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[23])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[24]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[25])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[26]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[27])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[28]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[29])
      | (~ (IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[74])));
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_11_sva = conv_s2s_44_45(IntSignedShiftRight_12U_6U_26U_mbits_fixed_11_sva[74:31])
      + conv_u2s_1_45(cvt_11_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl);
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_11_sva = nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_11_sva[44:0];
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_11_sva = (IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_11_sva[44])
      & (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_11_sva[43:25]==19'b1111111111111111111)));
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_11_sva = ~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_11_sva[44])
      | (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_11_sva[43:25]!=19'b0000000000000000000))));
  assign cvt_11_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl = ~(MUX_v_24_2_2((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_11_sva[24:1]),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_11_sva));
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_11_sva = ~(MUX_v_24_2_2((cvt_11_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_11_sva));
  assign cvt_12_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_6_nl = (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[30])
      & ((IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[0]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[1])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[2]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[3])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[4]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[5])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[6]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[7])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[8]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[9])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[10]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[11])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[12]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[13])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[14]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[15])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[16]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[17])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[18]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[19])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[20]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[21])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[22]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[23])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[24]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[25])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[26]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[27])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[28]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[29])
      | (~ (IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[74])));
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_12_sva = conv_s2s_44_45(IntSignedShiftRight_12U_6U_26U_mbits_fixed_12_sva[74:31])
      + conv_u2s_1_45(cvt_12_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_6_nl);
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_12_sva = nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_12_sva[44:0];
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_12_sva = (IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_12_sva[44])
      & (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_12_sva[43:25]==19'b1111111111111111111)));
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_12_sva = ~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_12_sva[44])
      | (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_12_sva[43:25]!=19'b0000000000000000000))));
  assign cvt_12_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_17_nl = ~(MUX_v_24_2_2((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_12_sva[24:1]),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_12_sva));
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_12_sva = ~(MUX_v_24_2_2((cvt_12_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_17_nl),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_12_sva));
  assign cvt_13_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl = (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[30])
      & ((IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[0]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[1])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[2]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[3])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[4]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[5])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[6]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[7])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[8]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[9])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[10]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[11])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[12]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[13])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[14]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[15])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[16]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[17])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[18]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[19])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[20]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[21])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[22]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[23])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[24]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[25])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[26]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[27])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[28]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[29])
      | (~ (IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[74])));
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_13_sva = conv_s2s_44_45(IntSignedShiftRight_12U_6U_26U_mbits_fixed_13_sva[74:31])
      + conv_u2s_1_45(cvt_13_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_4_nl);
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_13_sva = nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_13_sva[44:0];
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_13_sva = (IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_13_sva[44])
      & (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_13_sva[43:25]==19'b1111111111111111111)));
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_13_sva = ~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_13_sva[44])
      | (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_13_sva[43:25]!=19'b0000000000000000000))));
  assign cvt_13_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl = ~(MUX_v_24_2_2((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_13_sva[24:1]),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_13_sva));
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_13_sva = ~(MUX_v_24_2_2((cvt_13_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_12_nl),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_13_sva));
  assign cvt_14_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_6_nl = (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[30])
      & ((IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[0]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[1])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[2]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[3])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[4]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[5])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[6]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[7])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[8]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[9])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[10]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[11])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[12]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[13])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[14]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[15])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[16]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[17])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[18]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[19])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[20]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[21])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[22]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[23])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[24]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[25])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[26]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[27])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[28]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[29])
      | (~ (IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[74])));
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_14_sva = conv_s2s_44_45(IntSignedShiftRight_12U_6U_26U_mbits_fixed_14_sva[74:31])
      + conv_u2s_1_45(cvt_14_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_6_nl);
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_14_sva = nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_14_sva[44:0];
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_14_sva = (IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_14_sva[44])
      & (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_14_sva[43:25]==19'b1111111111111111111)));
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_14_sva = ~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_14_sva[44])
      | (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_14_sva[43:25]!=19'b0000000000000000000))));
  assign cvt_14_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_17_nl = ~(MUX_v_24_2_2((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_14_sva[24:1]),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_14_sva));
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_14_sva = ~(MUX_v_24_2_2((cvt_14_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_17_nl),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_14_sva));
  assign cvt_15_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_6_nl = (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[30])
      & ((IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[0]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[1])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[2]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[3])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[4]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[5])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[6]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[7])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[8]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[9])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[10]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[11])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[12]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[13])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[14]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[15])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[16]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[17])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[18]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[19])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[20]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[21])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[22]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[23])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[24]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[25])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[26]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[27])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[28]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[29])
      | (~ (IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[74])));
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_15_sva = conv_s2s_44_45(IntSignedShiftRight_12U_6U_26U_mbits_fixed_15_sva[74:31])
      + conv_u2s_1_45(cvt_15_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_6_nl);
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_15_sva = nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_15_sva[44:0];
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_15_sva = (IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_15_sva[44])
      & (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_15_sva[43:25]==19'b1111111111111111111)));
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_15_sva = ~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_15_sva[44])
      | (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_15_sva[43:25]!=19'b0000000000000000000))));
  assign cvt_15_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_17_nl = ~(MUX_v_24_2_2((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_15_sva[24:1]),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_15_sva));
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_15_sva = ~(MUX_v_24_2_2((cvt_15_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_17_nl),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_15_sva));
  assign cvt_16_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_8_nl = (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[30])
      & ((IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[0]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[1])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[2]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[3])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[4]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[5])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[6]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[7])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[8]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[9])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[10]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[11])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[12]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[13])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[14]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[15])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[16]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[17])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[18]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[19])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[20]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[21])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[22]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[23])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[24]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[25])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[26]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[27])
      | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[28]) | (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[29])
      | (~ (IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[74])));
  assign nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_sva = conv_s2s_44_45(IntSignedShiftRight_12U_6U_26U_mbits_fixed_sva[74:31])
      + conv_u2s_1_45(cvt_16_IntSignedShiftRight_12U_6U_26U_obits_fixed_and_8_nl);
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_sva = nl_IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_sva[44:0];
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_sva = (IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_sva[44])
      & (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_sva[43:25]==19'b1111111111111111111)));
  assign IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_sva = ~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_sva[44])
      | (~((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_sva[43:25]!=19'b0000000000000000000))));
  assign cvt_16_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_22_nl = ~(MUX_v_24_2_2((IntSignedShiftRight_12U_6U_26U_obits_fixed_acc_sat_sva[24:1]),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_ovfl_sva));
  assign FpFloatToInt_16U_5U_10U_internal_int_24_1_sva = ~(MUX_v_24_2_2((cvt_16_IntSignedShiftRight_12U_6U_26U_obits_fixed_nor_22_nl),
      24'b111111111111111111111111, IntSignedShiftRight_12U_6U_26U_obits_fixed_and_unfl_sva));
  assign nl_cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_1_nl = ({1'b1 , (~
      (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_16[4:1]))})
      + 5'b1;
  assign cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_1_nl = nl_cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_1_nl[4:0];
  assign cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_1_itm_4 = readslicef_5_1_4((cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_1_nl));
  assign FpMantRNE_17U_11U_else_carry_1_sva = (FpIntToFloat_17U_5U_10U_else_int_mant_1_sva[5])
      & ((FpIntToFloat_17U_5U_10U_else_int_mant_1_sva[0]) | (FpIntToFloat_17U_5U_10U_else_int_mant_1_sva[1])
      | (FpIntToFloat_17U_5U_10U_else_int_mant_1_sva[2]) | (FpIntToFloat_17U_5U_10U_else_int_mant_1_sva[3])
      | (FpIntToFloat_17U_5U_10U_else_int_mant_1_sva[4]) | (FpIntToFloat_17U_5U_10U_else_int_mant_1_sva[6]));
  assign nl_cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl = ({1'b1 , (~
      (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_17[4:1]))})
      + 5'b1;
  assign cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl = nl_cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl[4:0];
  assign cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4 = readslicef_5_1_4((cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl));
  assign FpMantRNE_17U_11U_else_carry_2_sva = (FpIntToFloat_17U_5U_10U_else_int_mant_2_sva[5])
      & ((FpIntToFloat_17U_5U_10U_else_int_mant_2_sva[0]) | (FpIntToFloat_17U_5U_10U_else_int_mant_2_sva[1])
      | (FpIntToFloat_17U_5U_10U_else_int_mant_2_sva[2]) | (FpIntToFloat_17U_5U_10U_else_int_mant_2_sva[3])
      | (FpIntToFloat_17U_5U_10U_else_int_mant_2_sva[4]) | (FpIntToFloat_17U_5U_10U_else_int_mant_2_sva[6]));
  assign nl_cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl = ({1'b1 , (~
      (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_18[4:1]))})
      + 5'b1;
  assign cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl = nl_cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl[4:0];
  assign cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4 = readslicef_5_1_4((cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl));
  assign FpMantRNE_17U_11U_else_carry_3_sva = (cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[5])
      & ((cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[0]) | (cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[1])
      | (cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[2]) | (cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[3])
      | (cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[4]) | (cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[6]));
  assign nl_cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl = ({1'b1 , (~
      (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_19[4:1]))})
      + 5'b1;
  assign cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl = nl_cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4:0];
  assign cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4 = readslicef_5_1_4((cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl));
  assign FpMantRNE_17U_11U_else_carry_4_sva = (cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[5])
      & ((cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[0]) | (cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[1])
      | (cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[2]) | (cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[3])
      | (cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[4]) | (cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[6]));
  assign nl_cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl = ({1'b1 , (~
      (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_20[4:1]))})
      + 5'b1;
  assign cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl = nl_cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl[4:0];
  assign cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4 = readslicef_5_1_4((cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl));
  assign FpMantRNE_17U_11U_else_carry_5_sva = (cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[5])
      & ((cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[0]) | (cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[1])
      | (cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[2]) | (cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[3])
      | (cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[4]) | (cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[6]));
  assign nl_cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl = ({1'b1 , (~
      (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_21[4:1]))})
      + 5'b1;
  assign cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl = nl_cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4:0];
  assign cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4 = readslicef_5_1_4((cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl));
  assign FpMantRNE_17U_11U_else_carry_6_sva = (cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[5])
      & ((cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[0]) | (cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[1])
      | (cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[2]) | (cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[3])
      | (cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[4]) | (cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[6]));
  assign nl_cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl = ({1'b1 , (~
      (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_22[4:1]))})
      + 5'b1;
  assign cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl = nl_cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4:0];
  assign cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4 = readslicef_5_1_4((cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl));
  assign FpMantRNE_17U_11U_else_carry_7_sva = (cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[5])
      & ((cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[0]) | (cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[1])
      | (cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[2]) | (cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[3])
      | (cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[4]) | (cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[6]));
  assign nl_cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl = ({1'b1 , (~
      (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_23[4:1]))})
      + 5'b1;
  assign cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl = nl_cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl[4:0];
  assign cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4 = readslicef_5_1_4((cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl));
  assign FpMantRNE_17U_11U_else_carry_8_sva = (cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[5])
      & ((cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[0]) | (cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[1])
      | (cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[2]) | (cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[3])
      | (cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[4]) | (cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[6]));
  assign nl_cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl = ({1'b1 , (~
      (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_24[4:1]))})
      + 5'b1;
  assign cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl = nl_cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl[4:0];
  assign cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4 = readslicef_5_1_4((cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_nl));
  assign FpMantRNE_17U_11U_else_carry_9_sva = (FpIntToFloat_17U_5U_10U_else_int_mant_9_sva[5])
      & ((FpIntToFloat_17U_5U_10U_else_int_mant_9_sva[0]) | (FpIntToFloat_17U_5U_10U_else_int_mant_9_sva[1])
      | (FpIntToFloat_17U_5U_10U_else_int_mant_9_sva[2]) | (FpIntToFloat_17U_5U_10U_else_int_mant_9_sva[3])
      | (FpIntToFloat_17U_5U_10U_else_int_mant_9_sva[4]) | (FpIntToFloat_17U_5U_10U_else_int_mant_9_sva[6]));
  assign nl_cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl = ({1'b1 ,
      (~ (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_25[4:1]))})
      + 5'b1;
  assign cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl = nl_cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4:0];
  assign cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4 = readslicef_5_1_4((cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl));
  assign FpMantRNE_17U_11U_else_carry_10_sva = (cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[5])
      & ((cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[0]) | (cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[1])
      | (cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[2]) | (cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[3])
      | (cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[4]) | (cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[6]));
  assign nl_cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl = ({1'b1 ,
      (~ (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_26[4:1]))})
      + 5'b1;
  assign cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl = nl_cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4:0];
  assign cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4 = readslicef_5_1_4((cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl));
  assign FpMantRNE_17U_11U_else_carry_11_sva = (cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[5])
      & ((cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[0]) | (cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[1])
      | (cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[2]) | (cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[3])
      | (cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[4]) | (cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[6]));
  assign nl_cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl = ({1'b1 ,
      (~ (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_27[4:1]))})
      + 5'b1;
  assign cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl = nl_cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl[4:0];
  assign cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4 = readslicef_5_1_4((cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl));
  assign FpMantRNE_17U_11U_else_carry_12_sva = (cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[5])
      & ((cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[0]) | (cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[1])
      | (cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[2]) | (cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[3])
      | (cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[4]) | (cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[6]));
  assign nl_cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl = ({1'b1 ,
      (~ (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_28[4:1]))})
      + 5'b1;
  assign cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl = nl_cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl[4:0];
  assign cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4 = readslicef_5_1_4((cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_nl));
  assign FpMantRNE_17U_11U_else_carry_13_sva = (cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[5])
      & ((cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[0]) | (cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[1])
      | (cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[2]) | (cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[3])
      | (cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[4]) | (cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[6]));
  assign nl_cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl = ({1'b1 ,
      (~ (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_29[4:1]))})
      + 5'b1;
  assign cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl = nl_cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl[4:0];
  assign cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4 = readslicef_5_1_4((cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl));
  assign FpMantRNE_17U_11U_else_carry_14_sva = (cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[5])
      & ((cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[0]) | (cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[1])
      | (cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[2]) | (cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[3])
      | (cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[4]) | (cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[6]));
  assign nl_cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl = ({1'b1 ,
      (~ (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_30[4:1]))})
      + 5'b1;
  assign cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl = nl_cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl[4:0];
  assign cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4 = readslicef_5_1_4((cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_nl));
  assign FpMantRNE_17U_11U_else_carry_15_sva = (cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[5])
      & ((cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[0]) | (cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[1])
      | (cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[2]) | (cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[3])
      | (cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[4]) | (cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[6]));
  assign nl_cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_8_nl = ({1'b1 ,
      (~ (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_31[4:1]))})
      + 5'b1;
  assign cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_8_nl = nl_cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_8_nl[4:0];
  assign cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_8_tmp_4 = readslicef_5_1_4((cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_8_nl));
  assign FpMantRNE_17U_11U_else_carry_sva = (cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_tmp[5])
      & ((cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_tmp[0]) | (cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_tmp[1])
      | (cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_tmp[2]) | (cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_tmp[3])
      | (cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_tmp[4]) | (cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_tmp[6]));
  assign cvt_if_unequal_tmp = ~((cfg_out_precision_1_sva_6==2'b01));
  assign FpIntToFloat_17U_5U_10U_o_mant_1_lpi_1_dfm_1 = MUX_v_10_2_2(reg_chn_idata_data_sva_3_15_0_2_reg,
      10'b1111111111, FpIntToFloat_17U_5U_10U_is_inf_1_lpi_1_dfm_6);
  assign nl_cvt_1_IntSaturation_17U_8U_else_if_acc_nl = conv_s2u_10_11({IntShiftRightSat_49U_6U_17U_o_16_1_sva_4
      , reg_chn_idata_data_sva_3_15_0_1_reg , (reg_chn_idata_data_sva_3_15_0_2_reg[9:6])})
      + 11'b1;
  assign cvt_1_IntSaturation_17U_8U_else_if_acc_nl = nl_cvt_1_IntSaturation_17U_8U_else_if_acc_nl[10:0];
  assign cvt_1_IntSaturation_17U_8U_else_if_acc_itm_10 = readslicef_11_1_10((cvt_1_IntSaturation_17U_8U_else_if_acc_nl));
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_nl = ~(cvt_1_IntSaturation_17U_8U_else_if_acc_itm_10
      | FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_2);
  assign IntSaturation_17U_8U_and_1_nl = cvt_1_IntSaturation_17U_8U_else_if_acc_itm_10
      & (~ FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_2);
  assign IntSaturation_17U_8U_o_7_1_1_lpi_1_dfm_1 = MUX1HOT_v_7_3_2((reg_chn_idata_data_sva_3_15_0_2_reg[6:0]),
      7'b1000000, 7'b111111, {(IntSaturation_17U_8U_IntSaturation_17U_8U_nor_nl)
      , (IntSaturation_17U_8U_and_1_nl) , FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_2});
  assign FpIntToFloat_17U_5U_10U_o_mant_2_lpi_1_dfm_1 = MUX_v_10_2_2(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_1_reg,
      10'b1111111111, FpIntToFloat_17U_5U_10U_is_inf_2_lpi_1_dfm_6);
  assign nl_cvt_2_IntSaturation_17U_8U_else_if_acc_1_nl = conv_s2u_10_11({IntShiftRightSat_49U_6U_17U_o_16_2_sva_3
      , reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_reg , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_1_reg[9:6])})
      + 11'b1;
  assign cvt_2_IntSaturation_17U_8U_else_if_acc_1_nl = nl_cvt_2_IntSaturation_17U_8U_else_if_acc_1_nl[10:0];
  assign cvt_2_IntSaturation_17U_8U_else_if_acc_1_itm_10 = readslicef_11_1_10((cvt_2_IntSaturation_17U_8U_else_if_acc_1_nl));
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_1_nl = ~(cvt_2_IntSaturation_17U_8U_else_if_acc_1_itm_10
      | FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_2);
  assign IntSaturation_17U_8U_and_3_nl = cvt_2_IntSaturation_17U_8U_else_if_acc_1_itm_10
      & (~ FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_2);
  assign IntSaturation_17U_8U_o_7_1_2_lpi_1_dfm_1 = MUX1HOT_v_7_3_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_1_reg[6:0]),
      7'b1000000, 7'b111111, {(IntSaturation_17U_8U_IntSaturation_17U_8U_nor_1_nl)
      , (IntSaturation_17U_8U_and_3_nl) , FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_2});
  assign and_2136_cse = (cfg_out_precision_1_sva_6==2'b11);
  assign cvt_else_nor_dfs = ~(cvt_else_equal_tmp | cvt_else_equal_tmp_1 | and_2136_cse);
  assign cvt_else_equal_tmp_1 = ~((cfg_out_precision_1_sva_6!=2'b00));
  assign cvt_else_equal_tmp = (cfg_out_precision_1_sva_6==2'b01);
  assign FpIntToFloat_17U_5U_10U_o_mant_3_lpi_1_dfm_1 = MUX_v_10_2_2(FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_7_itm_1,
      10'b1111111111, FpIntToFloat_17U_5U_10U_is_inf_3_lpi_1_dfm_7);
  assign nl_cvt_3_IntSaturation_17U_8U_else_if_acc_1_nl = conv_s2u_10_11({IntShiftRightSat_49U_6U_17U_o_16_3_sva_4
      , reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_reg , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_1_reg[9:6])})
      + 11'b1;
  assign cvt_3_IntSaturation_17U_8U_else_if_acc_1_nl = nl_cvt_3_IntSaturation_17U_8U_else_if_acc_1_nl[10:0];
  assign cvt_3_IntSaturation_17U_8U_else_if_acc_1_itm_10 = readslicef_11_1_10((cvt_3_IntSaturation_17U_8U_else_if_acc_1_nl));
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_2_nl = ~(cvt_3_IntSaturation_17U_8U_else_if_acc_1_itm_10
      | FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_2);
  assign IntSaturation_17U_8U_and_5_nl = cvt_3_IntSaturation_17U_8U_else_if_acc_1_itm_10
      & (~ FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_2);
  assign IntSaturation_17U_8U_o_7_1_3_lpi_1_dfm_1 = MUX1HOT_v_7_3_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_1_reg[6:0]),
      7'b1000000, 7'b111111, {(IntSaturation_17U_8U_IntSaturation_17U_8U_nor_2_nl)
      , (IntSaturation_17U_8U_and_5_nl) , FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_2});
  assign FpIntToFloat_17U_5U_10U_o_mant_4_lpi_1_dfm_1 = MUX_v_10_2_2(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_1_reg,
      10'b1111111111, FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_7);
  assign nl_cvt_4_IntSaturation_17U_8U_else_if_acc_2_nl = conv_s2u_10_11({IntShiftRightSat_49U_6U_17U_o_16_4_sva_3
      , (FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5[14:6])}) + 11'b1;
  assign cvt_4_IntSaturation_17U_8U_else_if_acc_2_nl = nl_cvt_4_IntSaturation_17U_8U_else_if_acc_2_nl[10:0];
  assign cvt_4_IntSaturation_17U_8U_else_if_acc_2_itm_10 = readslicef_11_1_10((cvt_4_IntSaturation_17U_8U_else_if_acc_2_nl));
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_3_nl = ~(cvt_4_IntSaturation_17U_8U_else_if_acc_2_itm_10
      | FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_2);
  assign IntSaturation_17U_8U_and_7_nl = cvt_4_IntSaturation_17U_8U_else_if_acc_2_itm_10
      & (~ FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_2);
  assign IntSaturation_17U_8U_o_7_1_4_lpi_1_dfm_1 = MUX1HOT_v_7_3_2((FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5[6:0]),
      7'b1000000, 7'b111111, {(IntSaturation_17U_8U_IntSaturation_17U_8U_nor_3_nl)
      , (IntSaturation_17U_8U_and_7_nl) , FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_2});
  assign FpIntToFloat_17U_5U_10U_o_mant_5_lpi_1_dfm_1 = MUX_v_10_2_2(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_1_reg,
      10'b1111111111, FpIntToFloat_17U_5U_10U_is_inf_5_lpi_1_dfm_7);
  assign nl_cvt_5_IntSaturation_17U_8U_else_if_acc_1_nl = conv_s2u_10_11({IntShiftRightSat_49U_6U_17U_o_16_5_sva_4
      , reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_reg , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_1_reg[9:6])})
      + 11'b1;
  assign cvt_5_IntSaturation_17U_8U_else_if_acc_1_nl = nl_cvt_5_IntSaturation_17U_8U_else_if_acc_1_nl[10:0];
  assign cvt_5_IntSaturation_17U_8U_else_if_acc_1_itm_10 = readslicef_11_1_10((cvt_5_IntSaturation_17U_8U_else_if_acc_1_nl));
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_4_nl = ~(cvt_5_IntSaturation_17U_8U_else_if_acc_1_itm_10
      | FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_2);
  assign IntSaturation_17U_8U_and_9_nl = cvt_5_IntSaturation_17U_8U_else_if_acc_1_itm_10
      & (~ FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_2);
  assign IntSaturation_17U_8U_o_7_1_5_lpi_1_dfm_1 = MUX1HOT_v_7_3_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_1_reg[6:0]),
      7'b1000000, 7'b111111, {(IntSaturation_17U_8U_IntSaturation_17U_8U_nor_4_nl)
      , (IntSaturation_17U_8U_and_9_nl) , FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_2});
  assign FpIntToFloat_17U_5U_10U_o_mant_6_lpi_1_dfm_1 = MUX_v_10_2_2(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_1_reg,
      10'b1111111111, FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_7);
  assign nl_cvt_6_IntSaturation_17U_8U_else_if_acc_2_nl = conv_s2u_10_11({IntShiftRightSat_49U_6U_17U_o_16_6_sva_3
      , reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_reg , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_1_reg[9:6])})
      + 11'b1;
  assign cvt_6_IntSaturation_17U_8U_else_if_acc_2_nl = nl_cvt_6_IntSaturation_17U_8U_else_if_acc_2_nl[10:0];
  assign cvt_6_IntSaturation_17U_8U_else_if_acc_2_itm_10 = readslicef_11_1_10((cvt_6_IntSaturation_17U_8U_else_if_acc_2_nl));
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_5_nl = ~(cvt_6_IntSaturation_17U_8U_else_if_acc_2_itm_10
      | FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_2);
  assign IntSaturation_17U_8U_and_11_nl = cvt_6_IntSaturation_17U_8U_else_if_acc_2_itm_10
      & (~ FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_2);
  assign IntSaturation_17U_8U_o_7_1_6_lpi_1_dfm_1 = MUX1HOT_v_7_3_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_1_reg[6:0]),
      7'b1000000, 7'b111111, {(IntSaturation_17U_8U_IntSaturation_17U_8U_nor_5_nl)
      , (IntSaturation_17U_8U_and_11_nl) , FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_2});
  assign FpIntToFloat_17U_5U_10U_o_mant_7_lpi_1_dfm_1 = MUX_v_10_2_2(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_1_reg,
      10'b1111111111, FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_7);
  assign nl_cvt_7_IntSaturation_17U_8U_else_if_acc_2_nl = conv_s2u_10_11({IntShiftRightSat_49U_6U_17U_o_16_7_sva_3
      , reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_reg , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_1_reg[9:6])})
      + 11'b1;
  assign cvt_7_IntSaturation_17U_8U_else_if_acc_2_nl = nl_cvt_7_IntSaturation_17U_8U_else_if_acc_2_nl[10:0];
  assign cvt_7_IntSaturation_17U_8U_else_if_acc_2_itm_10 = readslicef_11_1_10((cvt_7_IntSaturation_17U_8U_else_if_acc_2_nl));
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_6_nl = ~(cvt_7_IntSaturation_17U_8U_else_if_acc_2_itm_10
      | FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_2);
  assign IntSaturation_17U_8U_and_13_nl = cvt_7_IntSaturation_17U_8U_else_if_acc_2_itm_10
      & (~ FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_2);
  assign IntSaturation_17U_8U_o_7_1_7_lpi_1_dfm_1 = MUX1HOT_v_7_3_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_1_reg[6:0]),
      7'b1000000, 7'b111111, {(IntSaturation_17U_8U_IntSaturation_17U_8U_nor_6_nl)
      , (IntSaturation_17U_8U_and_13_nl) , FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_2});
  assign FpIntToFloat_17U_5U_10U_o_mant_8_lpi_1_dfm_1 = MUX_v_10_2_2(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_1_reg,
      10'b1111111111, FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_8);
  assign nl_cvt_8_IntSaturation_17U_8U_else_if_acc_3_nl = conv_s2u_10_11({IntShiftRightSat_49U_6U_17U_o_16_8_sva_3
      , reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_reg , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_1_reg[9:6])})
      + 11'b1;
  assign cvt_8_IntSaturation_17U_8U_else_if_acc_3_nl = nl_cvt_8_IntSaturation_17U_8U_else_if_acc_3_nl[10:0];
  assign cvt_8_IntSaturation_17U_8U_else_if_acc_3_itm_10 = readslicef_11_1_10((cvt_8_IntSaturation_17U_8U_else_if_acc_3_nl));
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_7_nl = ~(cvt_8_IntSaturation_17U_8U_else_if_acc_3_itm_10
      | FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_2);
  assign IntSaturation_17U_8U_and_15_nl = cvt_8_IntSaturation_17U_8U_else_if_acc_3_itm_10
      & (~ FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_2);
  assign IntSaturation_17U_8U_o_7_1_8_lpi_1_dfm_1 = MUX1HOT_v_7_3_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_1_reg[6:0]),
      7'b1000000, 7'b111111, {(IntSaturation_17U_8U_IntSaturation_17U_8U_nor_7_nl)
      , (IntSaturation_17U_8U_and_15_nl) , FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_2});
  assign FpIntToFloat_17U_5U_10U_o_mant_9_lpi_1_dfm_1 = MUX_v_10_2_2(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_1_reg,
      10'b1111111111, FpIntToFloat_17U_5U_10U_is_inf_9_lpi_1_dfm_7);
  assign nl_cvt_9_IntSaturation_17U_8U_else_if_acc_1_nl = conv_s2u_10_11({IntShiftRightSat_49U_6U_17U_o_16_9_sva_4
      , reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_reg , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_1_reg[9:6])})
      + 11'b1;
  assign cvt_9_IntSaturation_17U_8U_else_if_acc_1_nl = nl_cvt_9_IntSaturation_17U_8U_else_if_acc_1_nl[10:0];
  assign cvt_9_IntSaturation_17U_8U_else_if_acc_1_itm_10 = readslicef_11_1_10((cvt_9_IntSaturation_17U_8U_else_if_acc_1_nl));
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_8_nl = ~(cvt_9_IntSaturation_17U_8U_else_if_acc_1_itm_10
      | FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_2);
  assign IntSaturation_17U_8U_and_17_nl = cvt_9_IntSaturation_17U_8U_else_if_acc_1_itm_10
      & (~ FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_2);
  assign IntSaturation_17U_8U_o_7_1_9_lpi_1_dfm_1 = MUX1HOT_v_7_3_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_1_reg[6:0]),
      7'b1000000, 7'b111111, {(IntSaturation_17U_8U_IntSaturation_17U_8U_nor_8_nl)
      , (IntSaturation_17U_8U_and_17_nl) , FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_2});
  assign FpIntToFloat_17U_5U_10U_o_mant_10_lpi_1_dfm_1 = MUX_v_10_2_2(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_1_reg,
      10'b1111111111, FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_7);
  assign nl_cvt_10_IntSaturation_17U_8U_else_if_acc_2_nl = conv_s2u_10_11({IntShiftRightSat_49U_6U_17U_o_16_10_sva_3
      , reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_reg , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_1_reg[9:6])})
      + 11'b1;
  assign cvt_10_IntSaturation_17U_8U_else_if_acc_2_nl = nl_cvt_10_IntSaturation_17U_8U_else_if_acc_2_nl[10:0];
  assign cvt_10_IntSaturation_17U_8U_else_if_acc_2_itm_10 = readslicef_11_1_10((cvt_10_IntSaturation_17U_8U_else_if_acc_2_nl));
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_9_nl = ~(cvt_10_IntSaturation_17U_8U_else_if_acc_2_itm_10
      | FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_2);
  assign IntSaturation_17U_8U_and_19_nl = cvt_10_IntSaturation_17U_8U_else_if_acc_2_itm_10
      & (~ FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_2);
  assign IntSaturation_17U_8U_o_7_1_10_lpi_1_dfm_1 = MUX1HOT_v_7_3_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_1_reg[6:0]),
      7'b1000000, 7'b111111, {(IntSaturation_17U_8U_IntSaturation_17U_8U_nor_9_nl)
      , (IntSaturation_17U_8U_and_19_nl) , FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_2});
  assign FpIntToFloat_17U_5U_10U_o_mant_11_lpi_1_dfm_1 = MUX_v_10_2_2(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_1_reg,
      10'b1111111111, FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_7);
  assign nl_cvt_11_IntSaturation_17U_8U_else_if_acc_2_nl = conv_s2u_10_11({IntShiftRightSat_49U_6U_17U_o_16_11_sva_3
      , reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_reg , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_1_reg[9:6])})
      + 11'b1;
  assign cvt_11_IntSaturation_17U_8U_else_if_acc_2_nl = nl_cvt_11_IntSaturation_17U_8U_else_if_acc_2_nl[10:0];
  assign cvt_11_IntSaturation_17U_8U_else_if_acc_2_itm_10 = readslicef_11_1_10((cvt_11_IntSaturation_17U_8U_else_if_acc_2_nl));
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_10_nl = ~(cvt_11_IntSaturation_17U_8U_else_if_acc_2_itm_10
      | FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_2);
  assign IntSaturation_17U_8U_and_21_nl = cvt_11_IntSaturation_17U_8U_else_if_acc_2_itm_10
      & (~ FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_2);
  assign IntSaturation_17U_8U_o_7_1_11_lpi_1_dfm_1 = MUX1HOT_v_7_3_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_1_reg[6:0]),
      7'b1000000, 7'b111111, {(IntSaturation_17U_8U_IntSaturation_17U_8U_nor_10_nl)
      , (IntSaturation_17U_8U_and_21_nl) , FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_2});
  assign FpIntToFloat_17U_5U_10U_o_mant_12_lpi_1_dfm_1 = MUX_v_10_2_2(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_1_reg,
      10'b1111111111, FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_8);
  assign nl_cvt_12_IntSaturation_17U_8U_else_if_acc_3_nl = conv_s2u_10_11({IntShiftRightSat_49U_6U_17U_o_16_12_sva_3
      , reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_reg , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_1_reg[9:6])})
      + 11'b1;
  assign cvt_12_IntSaturation_17U_8U_else_if_acc_3_nl = nl_cvt_12_IntSaturation_17U_8U_else_if_acc_3_nl[10:0];
  assign cvt_12_IntSaturation_17U_8U_else_if_acc_3_itm_10 = readslicef_11_1_10((cvt_12_IntSaturation_17U_8U_else_if_acc_3_nl));
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_11_nl = ~(cvt_12_IntSaturation_17U_8U_else_if_acc_3_itm_10
      | FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_2);
  assign IntSaturation_17U_8U_and_23_nl = cvt_12_IntSaturation_17U_8U_else_if_acc_3_itm_10
      & (~ FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_2);
  assign IntSaturation_17U_8U_o_7_1_12_lpi_1_dfm_1 = MUX1HOT_v_7_3_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_1_reg[6:0]),
      7'b1000000, 7'b111111, {(IntSaturation_17U_8U_IntSaturation_17U_8U_nor_11_nl)
      , (IntSaturation_17U_8U_and_23_nl) , FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_2});
  assign FpIntToFloat_17U_5U_10U_o_mant_13_lpi_1_dfm_1 = MUX_v_10_2_2(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_1_reg,
      10'b1111111111, FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_7);
  assign nl_cvt_13_IntSaturation_17U_8U_else_if_acc_2_nl = conv_s2u_10_11({IntShiftRightSat_49U_6U_17U_o_16_13_sva_3
      , reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_reg , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_1_reg[9:6])})
      + 11'b1;
  assign cvt_13_IntSaturation_17U_8U_else_if_acc_2_nl = nl_cvt_13_IntSaturation_17U_8U_else_if_acc_2_nl[10:0];
  assign cvt_13_IntSaturation_17U_8U_else_if_acc_2_itm_10 = readslicef_11_1_10((cvt_13_IntSaturation_17U_8U_else_if_acc_2_nl));
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_12_nl = ~(cvt_13_IntSaturation_17U_8U_else_if_acc_2_itm_10
      | FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_2);
  assign IntSaturation_17U_8U_and_25_nl = cvt_13_IntSaturation_17U_8U_else_if_acc_2_itm_10
      & (~ FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_2);
  assign IntSaturation_17U_8U_o_7_1_13_lpi_1_dfm_1 = MUX1HOT_v_7_3_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_1_reg[6:0]),
      7'b1000000, 7'b111111, {(IntSaturation_17U_8U_IntSaturation_17U_8U_nor_12_nl)
      , (IntSaturation_17U_8U_and_25_nl) , FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_2});
  assign FpIntToFloat_17U_5U_10U_o_mant_14_lpi_1_dfm_1 = MUX_v_10_2_2(reg_IntShiftRightSat_49U_6U_17U_o_15_1_14_3_reg,
      10'b1111111111, FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_8);
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_13_nl = ~(cvt_14_IntSaturation_17U_8U_else_if_acc_3_itm_10
      | cvt_14_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_3_svs_1);
  assign IntSaturation_17U_8U_and_27_nl = cvt_14_IntSaturation_17U_8U_else_if_acc_3_itm_10
      & (~ cvt_14_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_3_svs_1);
  assign IntSaturation_17U_8U_o_7_1_14_lpi_1_dfm_1 = MUX1HOT_v_7_3_2((reg_IntShiftRightSat_49U_6U_17U_o_15_1_14_3_reg[6:0]),
      7'b1000000, 7'b111111, {(IntSaturation_17U_8U_IntSaturation_17U_8U_nor_13_nl)
      , (IntSaturation_17U_8U_and_27_nl) , cvt_14_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_3_svs_1});
  assign FpIntToFloat_17U_5U_10U_o_mant_15_lpi_1_dfm_1 = MUX_v_10_2_2(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_1_reg,
      10'b1111111111, FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_8);
  assign nl_cvt_15_IntSaturation_17U_8U_else_if_acc_3_nl = conv_s2u_10_11({IntShiftRightSat_49U_6U_17U_o_16_15_sva_3
      , reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_reg , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_1_reg[9:6])})
      + 11'b1;
  assign cvt_15_IntSaturation_17U_8U_else_if_acc_3_nl = nl_cvt_15_IntSaturation_17U_8U_else_if_acc_3_nl[10:0];
  assign cvt_15_IntSaturation_17U_8U_else_if_acc_3_itm_10 = readslicef_11_1_10((cvt_15_IntSaturation_17U_8U_else_if_acc_3_nl));
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_14_nl = ~(cvt_15_IntSaturation_17U_8U_else_if_acc_3_itm_10
      | FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_2);
  assign IntSaturation_17U_8U_and_29_nl = cvt_15_IntSaturation_17U_8U_else_if_acc_3_itm_10
      & (~ FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_2);
  assign IntSaturation_17U_8U_o_7_1_15_lpi_1_dfm_1 = MUX1HOT_v_7_3_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_1_reg[6:0]),
      7'b1000000, 7'b111111, {(IntSaturation_17U_8U_IntSaturation_17U_8U_nor_14_nl)
      , (IntSaturation_17U_8U_and_29_nl) , FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_2});
  assign FpIntToFloat_17U_5U_10U_o_mant_lpi_1_dfm_1 = MUX_v_10_2_2(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_1_reg,
      10'b1111111111, FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_9);
  assign nl_cvt_16_IntSaturation_17U_8U_else_if_acc_4_nl = conv_s2u_10_11({IntShiftRightSat_49U_6U_17U_o_16_sva_3
      , reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_reg , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_1_reg[9:6])})
      + 11'b1;
  assign cvt_16_IntSaturation_17U_8U_else_if_acc_4_nl = nl_cvt_16_IntSaturation_17U_8U_else_if_acc_4_nl[10:0];
  assign cvt_16_IntSaturation_17U_8U_else_if_acc_4_itm_10 = readslicef_11_1_10((cvt_16_IntSaturation_17U_8U_else_if_acc_4_nl));
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_nor_15_nl = ~(cvt_16_IntSaturation_17U_8U_else_if_acc_4_itm_10
      | FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_2);
  assign IntSaturation_17U_8U_and_31_nl = cvt_16_IntSaturation_17U_8U_else_if_acc_4_itm_10
      & (~ FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_2);
  assign IntSaturation_17U_8U_o_7_1_lpi_1_dfm_1 = MUX1HOT_v_7_3_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_1_reg[6:0]),
      7'b1000000, 7'b111111, {(IntSaturation_17U_8U_IntSaturation_17U_8U_nor_15_nl)
      , (IntSaturation_17U_8U_and_31_nl) , FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_2});
  assign nl_cvt_14_IntSaturation_17U_8U_else_if_acc_3_nl = conv_s2u_10_11({IntShiftRightSat_49U_6U_17U_o_16_14_sva_3
      , reg_IntShiftRightSat_49U_6U_17U_o_15_1_14_1_reg , (reg_IntShiftRightSat_49U_6U_17U_o_15_1_14_3_reg[9:6])})
      + 11'b1;
  assign cvt_14_IntSaturation_17U_8U_else_if_acc_3_nl = nl_cvt_14_IntSaturation_17U_8U_else_if_acc_3_nl[10:0];
  assign cvt_14_IntSaturation_17U_8U_else_if_acc_3_itm_10 = readslicef_11_1_10((cvt_14_IntSaturation_17U_8U_else_if_acc_3_nl));
  assign cvt_and_147_m1c = (~ cfg_mode_eql_1_sva_6) & cvt_unequal_tmp_21;
  assign main_stage_en_1 = chn_in_rsci_bawt & or_5189_cse;
  assign FpFloatToInt_16U_5U_10U_if_qr_1_lpi_1_dfm_mx0 = MUX_v_16_2_2(16'b111111111111111,
      16'b1000000000000000, chn_idata_data_sva_2_47_31_1[0]);
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_1_sva = ({(~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_1_sva[14:0]))
      , (~ FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_mx0w0)}) + 16'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_1_sva = nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_1_sva[15:0];
  assign FpFloatToInt_16U_5U_10U_if_qr_2_lpi_1_dfm_mx0 = MUX_v_16_2_2(16'b111111111111111,
      16'b1000000000000000, chn_idata_data_sva_2_79_63_1[0]);
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_2_sva = ({(~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_2_sva[14:0]))
      , (~ FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_mx0w0)}) + 16'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_2_sva = nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_2_sva[15:0];
  assign FpFloatToInt_16U_5U_10U_if_qr_3_lpi_1_dfm_mx0 = MUX_v_16_2_2(16'b111111111111111,
      16'b1000000000000000, chn_idata_data_sva_2_111_95_1[0]);
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_3_sva = ({(~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_3_sva[14:0]))
      , (~ FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_mx0w0)}) + 16'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_3_sva = nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_3_sva[15:0];
  assign FpFloatToInt_16U_5U_10U_if_qr_4_lpi_1_dfm_mx0 = MUX_v_16_2_2(16'b111111111111111,
      16'b1000000000000000, chn_idata_data_sva_2_143_127_1[0]);
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_4_sva = ({(~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_4_sva[14:0]))
      , (~ FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_mx0w0)}) + 16'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_4_sva = nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_4_sva[15:0];
  assign FpFloatToInt_16U_5U_10U_if_qr_5_lpi_1_dfm_mx0 = MUX_v_16_2_2(16'b111111111111111,
      16'b1000000000000000, chn_idata_data_sva_2_175_159_1[0]);
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_5_sva = ({(~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_5_sva[14:0]))
      , (~ FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_mx0w0)}) + 16'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_5_sva = nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_5_sva[15:0];
  assign FpFloatToInt_16U_5U_10U_if_qr_6_lpi_1_dfm_mx0 = MUX_v_16_2_2(16'b111111111111111,
      16'b1000000000000000, chn_idata_data_sva_2_207_191_1[0]);
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_6_sva = ({(~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_6_sva[14:0]))
      , (~ FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_mx0w0)}) + 16'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_6_sva = nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_6_sva[15:0];
  assign FpFloatToInt_16U_5U_10U_if_qr_7_lpi_1_dfm_mx0 = MUX_v_16_2_2(16'b111111111111111,
      16'b1000000000000000, chn_idata_data_sva_2_239_223_1[0]);
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_7_sva = ({(~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_7_sva[14:0]))
      , (~ FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_mx0w0)}) + 16'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_7_sva = nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_7_sva[15:0];
  assign FpFloatToInt_16U_5U_10U_if_qr_8_lpi_1_dfm_mx0 = MUX_v_16_2_2(16'b111111111111111,
      16'b1000000000000000, chn_idata_data_sva_2_271_255_1[0]);
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_8_sva = ({(~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_8_sva[14:0]))
      , (~ FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_mx0w0)}) + 16'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_8_sva = nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_8_sva[15:0];
  assign FpFloatToInt_16U_5U_10U_if_qr_9_lpi_1_dfm_mx0 = MUX_v_16_2_2(16'b111111111111111,
      16'b1000000000000000, chn_idata_data_sva_2_303_287_1[0]);
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_9_sva = ({(~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_9_sva[14:0]))
      , (~ FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_mx0w0)}) + 16'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_9_sva = nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_9_sva[15:0];
  assign FpFloatToInt_16U_5U_10U_if_qr_10_lpi_1_dfm_mx0 = MUX_v_16_2_2(16'b111111111111111,
      16'b1000000000000000, chn_idata_data_sva_2_335_319_1[0]);
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_10_sva = ({(~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_10_sva[14:0]))
      , (~ FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_mx0w0)}) + 16'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_10_sva = nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_10_sva[15:0];
  assign FpFloatToInt_16U_5U_10U_if_qr_11_lpi_1_dfm_mx0 = MUX_v_16_2_2(16'b111111111111111,
      16'b1000000000000000, chn_idata_data_sva_2_367_351_1[0]);
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_11_sva = ({(~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_11_sva[14:0]))
      , (~ FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_mx0w0)}) + 16'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_11_sva = nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_11_sva[15:0];
  assign FpFloatToInt_16U_5U_10U_if_qr_12_lpi_1_dfm_mx0 = MUX_v_16_2_2(16'b111111111111111,
      16'b1000000000000000, chn_idata_data_sva_2_399_383_1[0]);
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_12_sva = ({(~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_12_sva[14:0]))
      , (~ FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_mx0w0)}) + 16'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_12_sva = nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_12_sva[15:0];
  assign FpFloatToInt_16U_5U_10U_if_qr_13_lpi_1_dfm_mx0 = MUX_v_16_2_2(16'b111111111111111,
      16'b1000000000000000, chn_idata_data_sva_2_431_415_1[0]);
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_13_sva = ({(~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_13_sva[14:0]))
      , (~ FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_mx0w0)}) + 16'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_13_sva = nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_13_sva[15:0];
  assign FpFloatToInt_16U_5U_10U_if_qr_14_lpi_1_dfm_mx0 = MUX_v_16_2_2(16'b111111111111111,
      16'b1000000000000000, chn_idata_data_sva_2_463_447_1[0]);
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_14_sva = ({(~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_14_sva[14:0]))
      , (~ FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_mx0w0)}) + 16'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_14_sva = nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_14_sva[15:0];
  assign FpFloatToInt_16U_5U_10U_if_qr_15_lpi_1_dfm_mx0 = MUX_v_16_2_2(16'b111111111111111,
      16'b1000000000000000, chn_idata_data_sva_2_495_479_1[0]);
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_15_sva = ({(~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_15_sva[14:0]))
      , (~ FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_mx0w0)}) + 16'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_15_sva = nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_15_sva[15:0];
  assign FpFloatToInt_16U_5U_10U_if_qr_lpi_1_dfm_mx0 = MUX_v_16_2_2(16'b111111111111111,
      16'b1000000000000000, chn_idata_data_sva_2_511_1);
  assign nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_sva = ({(~ (FpFloatToInt_16U_5U_10U_internal_int_24_1_sva[14:0]))
      , (~ FpFloatToInt_16U_5U_10U_internal_int_0_sva_mx0w0)}) + 16'b1;
  assign FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_sva = nl_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_sva[15:0];
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_lpi_1_dfm_5_mx0 = MUX_v_10_2_2(FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_15_mx0w1,
      (chn_idata_data_sva_1_507_479_1[10:1]), IsNaN_8U_23U_land_lpi_1_dfm_3);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_15_lpi_1_dfm_5_mx0 = MUX_v_10_2_2(FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_14_mx0w1,
      (chn_idata_data_sva_1_475_447_1[10:1]), IsNaN_8U_23U_land_15_lpi_1_dfm_3);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_14_lpi_1_dfm_5_mx0 = MUX_v_10_2_2(FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_13_mx0w1,
      (chn_idata_data_sva_1_443_415_1[10:1]), IsNaN_8U_23U_land_14_lpi_1_dfm_3);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_13_lpi_1_dfm_5_mx0 = MUX_v_10_2_2(FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_12_mx0w1,
      (chn_idata_data_sva_1_411_383_1[10:1]), IsNaN_8U_23U_land_13_lpi_1_dfm_3);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_12_lpi_1_dfm_5_mx0 = MUX_v_10_2_2(FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_11_mx0w1,
      (chn_idata_data_sva_1_379_351_1[10:1]), IsNaN_8U_23U_land_12_lpi_1_dfm_3);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_11_lpi_1_dfm_5_mx0 = MUX_v_10_2_2(FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_10_mx0w1,
      (chn_idata_data_sva_1_347_319_1[10:1]), IsNaN_8U_23U_land_11_lpi_1_dfm_3);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_10_lpi_1_dfm_5_mx0 = MUX_v_10_2_2(FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_9_mx0w1,
      (chn_idata_data_sva_1_315_287_1[10:1]), IsNaN_8U_23U_land_10_lpi_1_dfm_3);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_9_lpi_1_dfm_5_mx0 = MUX_v_10_2_2(FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_8_mx0w1,
      (chn_idata_data_sva_1_283_255_1[10:1]), IsNaN_8U_23U_land_9_lpi_1_dfm_3);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_8_lpi_1_dfm_5_mx0 = MUX_v_10_2_2(FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_7_mx0w1,
      (chn_idata_data_sva_1_251_223_1[10:1]), IsNaN_8U_23U_land_8_lpi_1_dfm_3);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_7_lpi_1_dfm_5_mx0 = MUX_v_10_2_2(FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_6_mx0w1,
      (chn_idata_data_sva_1_219_191_1[10:1]), IsNaN_8U_23U_land_7_lpi_1_dfm_3);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_6_lpi_1_dfm_5_mx0 = MUX_v_10_2_2(FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_5_mx0w1,
      (chn_idata_data_sva_1_187_159_1[10:1]), IsNaN_8U_23U_land_6_lpi_1_dfm_3);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_5_lpi_1_dfm_5_mx0 = MUX_v_10_2_2((chn_idata_data_sva_1_155_127_1[10:1]),
      FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_4_mx0w1,
      or_tmp_2469);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_4_lpi_1_dfm_5_mx0 = MUX_v_10_2_2(FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_3_mx0w1,
      (chn_idata_data_sva_1_123_95_1[10:1]), IsNaN_8U_23U_land_4_lpi_1_dfm_3);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_3_lpi_1_dfm_5_mx0 = MUX_v_10_2_2(FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_2_mx0w1,
      (chn_idata_data_sva_1_91_63_1[10:1]), IsNaN_8U_23U_land_3_lpi_1_dfm_3);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_2_lpi_1_dfm_5_mx0 = MUX_v_10_2_2(FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_1_mx0w1,
      (chn_idata_data_sva_1_59_31_1[10:1]), IsNaN_8U_23U_land_2_lpi_1_dfm_3);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_1_lpi_1_dfm_5_mx0 = MUX_v_10_2_2(FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_mx0w1,
      (chn_idata_data_sva_1_27_0_1[9:0]), IsNaN_8U_23U_land_1_lpi_1_dfm_3);
  assign cvt_1_FpMantDecShiftRight_23U_8U_10U_carry_and_nl = ((FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_1_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_guard_mask_1_sva[23])) & ((FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_1_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_1_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_mask_1_sva[23]));
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_1_sva = (cvt_1_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_itm[23:13])
      + conv_u2u_1_11(cvt_1_FpMantDecShiftRight_23U_8U_10U_carry_and_nl);
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_1_sva = nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_1_sva[10:0];
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_1_sva = (chn_idata_data_sva_1_27_0_1[22:0])
      & (FpMantDecShiftRight_23U_8U_10U_guard_mask_1_sva[22:0]);
  assign nl_cvt_1_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl = (FpMantDecShiftRight_23U_8U_10U_guard_mask_1_sva[22:0])
      + 23'b11111111111111111111111;
  assign cvt_1_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl = nl_cvt_1_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_1_sva = (chn_idata_data_sva_1_27_0_1[22:0])
      & (cvt_1_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_nl);
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_1_sva = (chn_idata_data_sva_1_27_0_1[22:0])
      & (FpMantDecShiftRight_23U_8U_10U_least_mask_1_sva[22:0]);
  assign cvt_2_FpMantDecShiftRight_23U_8U_10U_carry_and_1_nl = ((FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_2_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_guard_mask_2_sva[23])) & ((FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_2_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_2_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_mask_2_sva[23]));
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_2_sva = (cvt_2_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_itm[23:13])
      + conv_u2u_1_11(cvt_2_FpMantDecShiftRight_23U_8U_10U_carry_and_1_nl);
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_2_sva = nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_2_sva[10:0];
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_2_sva = (chn_idata_data_sva_1_59_31_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_guard_mask_2_sva[22:0]);
  assign nl_cvt_2_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl = (FpMantDecShiftRight_23U_8U_10U_guard_mask_2_sva[22:0])
      + 23'b11111111111111111111111;
  assign cvt_2_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl = nl_cvt_2_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_2_sva = (chn_idata_data_sva_1_59_31_1[23:1])
      & (cvt_2_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl);
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_2_sva = (chn_idata_data_sva_1_59_31_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_least_mask_2_sva[22:0]);
  assign cvt_3_FpMantDecShiftRight_23U_8U_10U_carry_and_1_nl = ((FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_3_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_guard_mask_3_sva[23])) & ((FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_3_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_3_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_mask_3_sva[23]));
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_3_sva = (cvt_3_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_itm[23:13])
      + conv_u2u_1_11(cvt_3_FpMantDecShiftRight_23U_8U_10U_carry_and_1_nl);
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_3_sva = nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_3_sva[10:0];
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_3_sva = (chn_idata_data_sva_1_91_63_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_guard_mask_3_sva[22:0]);
  assign nl_cvt_3_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl = (FpMantDecShiftRight_23U_8U_10U_guard_mask_3_sva[22:0])
      + 23'b11111111111111111111111;
  assign cvt_3_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl = nl_cvt_3_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_3_sva = (chn_idata_data_sva_1_91_63_1[23:1])
      & (cvt_3_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl);
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_3_sva = (chn_idata_data_sva_1_91_63_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_least_mask_3_sva[22:0]);
  assign cvt_4_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl = ((FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_4_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_guard_mask_4_sva[23])) & ((FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_4_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_4_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_mask_4_sva[23]));
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_4_sva = (cvt_4_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm[23:13])
      + conv_u2u_1_11(cvt_4_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl);
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_4_sva = nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_4_sva[10:0];
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_4_sva = (chn_idata_data_sva_1_123_95_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_guard_mask_4_sva[22:0]);
  assign nl_cvt_4_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl = (FpMantDecShiftRight_23U_8U_10U_guard_mask_4_sva[22:0])
      + 23'b11111111111111111111111;
  assign cvt_4_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl = nl_cvt_4_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_4_sva = (chn_idata_data_sva_1_123_95_1[23:1])
      & (cvt_4_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl);
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_4_sva = (chn_idata_data_sva_1_123_95_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_least_mask_4_sva[22:0]);
  assign cvt_5_FpMantDecShiftRight_23U_8U_10U_carry_and_1_nl = ((FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_5_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_guard_mask_5_sva[23])) & ((FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_5_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_5_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_mask_5_sva[23]));
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_5_sva = (cvt_5_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_itm[23:13])
      + conv_u2u_1_11(cvt_5_FpMantDecShiftRight_23U_8U_10U_carry_and_1_nl);
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_5_sva = nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_5_sva[10:0];
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_5_sva = (chn_idata_data_sva_1_155_127_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_guard_mask_5_sva[22:0]);
  assign nl_cvt_5_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl = (FpMantDecShiftRight_23U_8U_10U_guard_mask_5_sva[22:0])
      + 23'b11111111111111111111111;
  assign cvt_5_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl = nl_cvt_5_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_5_sva = (chn_idata_data_sva_1_155_127_1[23:1])
      & (cvt_5_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl);
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_5_sva = (chn_idata_data_sva_1_155_127_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_least_mask_5_sva[22:0]);
  assign cvt_6_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl = ((FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_6_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_guard_mask_6_sva[23])) & ((FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_6_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_6_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_mask_6_sva[23]));
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_6_sva = (cvt_6_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm[23:13])
      + conv_u2u_1_11(cvt_6_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl);
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_6_sva = nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_6_sva[10:0];
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_6_sva = (chn_idata_data_sva_1_187_159_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_guard_mask_6_sva[22:0]);
  assign nl_cvt_6_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl = (FpMantDecShiftRight_23U_8U_10U_guard_mask_6_sva[22:0])
      + 23'b11111111111111111111111;
  assign cvt_6_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl = nl_cvt_6_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_6_sva = (chn_idata_data_sva_1_187_159_1[23:1])
      & (cvt_6_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl);
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_6_sva = (chn_idata_data_sva_1_187_159_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_least_mask_6_sva[22:0]);
  assign cvt_7_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl = ((FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_7_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_guard_mask_7_sva[23])) & ((FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_7_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_7_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_mask_7_sva[23]));
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_7_sva = (cvt_7_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm[23:13])
      + conv_u2u_1_11(cvt_7_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl);
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_7_sva = nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_7_sva[10:0];
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_7_sva = (chn_idata_data_sva_1_219_191_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_guard_mask_7_sva[22:0]);
  assign nl_cvt_7_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl = (FpMantDecShiftRight_23U_8U_10U_guard_mask_7_sva[22:0])
      + 23'b11111111111111111111111;
  assign cvt_7_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl = nl_cvt_7_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_7_sva = (chn_idata_data_sva_1_219_191_1[23:1])
      & (cvt_7_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl);
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_7_sva = (chn_idata_data_sva_1_219_191_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_least_mask_7_sva[22:0]);
  assign cvt_8_FpMantDecShiftRight_23U_8U_10U_carry_and_3_nl = ((FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_8_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_guard_mask_8_sva[23])) & ((FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_8_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_8_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_mask_8_sva[23]));
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_8_sva = (cvt_8_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_itm[23:13])
      + conv_u2u_1_11(cvt_8_FpMantDecShiftRight_23U_8U_10U_carry_and_3_nl);
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_8_sva = nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_8_sva[10:0];
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_8_sva = (chn_idata_data_sva_1_251_223_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_guard_mask_8_sva[22:0]);
  assign nl_cvt_8_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl = (FpMantDecShiftRight_23U_8U_10U_guard_mask_8_sva[22:0])
      + 23'b11111111111111111111111;
  assign cvt_8_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl = nl_cvt_8_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_8_sva = (chn_idata_data_sva_1_251_223_1[23:1])
      & (cvt_8_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl);
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_8_sva = (chn_idata_data_sva_1_251_223_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_least_mask_8_sva[22:0]);
  assign cvt_9_FpMantDecShiftRight_23U_8U_10U_carry_and_1_nl = ((FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_9_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_guard_mask_9_sva[23])) & ((FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_9_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_9_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_mask_9_sva[23]));
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_9_sva = (cvt_9_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_1_itm[23:13])
      + conv_u2u_1_11(cvt_9_FpMantDecShiftRight_23U_8U_10U_carry_and_1_nl);
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_9_sva = nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_9_sva[10:0];
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_9_sva = (chn_idata_data_sva_1_283_255_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_guard_mask_9_sva[22:0]);
  assign nl_cvt_9_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl = (FpMantDecShiftRight_23U_8U_10U_guard_mask_9_sva[22:0])
      + 23'b11111111111111111111111;
  assign cvt_9_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl = nl_cvt_9_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_9_sva = (chn_idata_data_sva_1_283_255_1[23:1])
      & (cvt_9_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_1_nl);
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_9_sva = (chn_idata_data_sva_1_283_255_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_least_mask_9_sva[22:0]);
  assign cvt_10_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl = ((FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_10_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_guard_mask_10_sva[23])) & ((FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_10_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_10_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_mask_10_sva[23]));
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_10_sva = (cvt_10_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm[23:13])
      + conv_u2u_1_11(cvt_10_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl);
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_10_sva = nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_10_sva[10:0];
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_10_sva = (chn_idata_data_sva_1_315_287_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_guard_mask_10_sva[22:0]);
  assign nl_cvt_10_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl = (FpMantDecShiftRight_23U_8U_10U_guard_mask_10_sva[22:0])
      + 23'b11111111111111111111111;
  assign cvt_10_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl = nl_cvt_10_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_10_sva = (chn_idata_data_sva_1_315_287_1[23:1])
      & (cvt_10_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl);
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_10_sva = (chn_idata_data_sva_1_315_287_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_least_mask_10_sva[22:0]);
  assign cvt_11_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl = ((FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_11_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_guard_mask_11_sva[23])) & ((FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_11_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_11_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_mask_11_sva[23]));
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_11_sva = (cvt_11_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm[23:13])
      + conv_u2u_1_11(cvt_11_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl);
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_11_sva = nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_11_sva[10:0];
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_11_sva = (chn_idata_data_sva_1_347_319_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_guard_mask_11_sva[22:0]);
  assign nl_cvt_11_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl = (FpMantDecShiftRight_23U_8U_10U_guard_mask_11_sva[22:0])
      + 23'b11111111111111111111111;
  assign cvt_11_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl = nl_cvt_11_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_11_sva = (chn_idata_data_sva_1_347_319_1[23:1])
      & (cvt_11_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl);
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_11_sva = (chn_idata_data_sva_1_347_319_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_least_mask_11_sva[22:0]);
  assign cvt_12_FpMantDecShiftRight_23U_8U_10U_carry_and_3_nl = ((FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_12_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_guard_mask_12_sva[23])) & ((FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_12_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_12_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_mask_12_sva[23]));
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_12_sva = (cvt_12_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_itm[23:13])
      + conv_u2u_1_11(cvt_12_FpMantDecShiftRight_23U_8U_10U_carry_and_3_nl);
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_12_sva = nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_12_sva[10:0];
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_12_sva = (chn_idata_data_sva_1_379_351_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_guard_mask_12_sva[22:0]);
  assign nl_cvt_12_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl = (FpMantDecShiftRight_23U_8U_10U_guard_mask_12_sva[22:0])
      + 23'b11111111111111111111111;
  assign cvt_12_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl = nl_cvt_12_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_12_sva = (chn_idata_data_sva_1_379_351_1[23:1])
      & (cvt_12_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl);
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_12_sva = (chn_idata_data_sva_1_379_351_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_least_mask_12_sva[22:0]);
  assign cvt_13_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl = ((FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_13_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_guard_mask_13_sva[23])) & ((FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_13_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_13_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_mask_13_sva[23]));
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_13_sva = (cvt_13_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_2_itm[23:13])
      + conv_u2u_1_11(cvt_13_FpMantDecShiftRight_23U_8U_10U_carry_and_2_nl);
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_13_sva = nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_13_sva[10:0];
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_13_sva = (chn_idata_data_sva_1_411_383_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_guard_mask_13_sva[22:0]);
  assign nl_cvt_13_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl = (FpMantDecShiftRight_23U_8U_10U_guard_mask_13_sva[22:0])
      + 23'b11111111111111111111111;
  assign cvt_13_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl = nl_cvt_13_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_13_sva = (chn_idata_data_sva_1_411_383_1[23:1])
      & (cvt_13_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_2_nl);
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_13_sva = (chn_idata_data_sva_1_411_383_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_least_mask_13_sva[22:0]);
  assign cvt_14_FpMantDecShiftRight_23U_8U_10U_carry_and_3_nl = ((FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_14_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_guard_mask_14_sva[23])) & ((FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_14_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_14_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_mask_14_sva[23]));
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_14_sva = (cvt_14_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_itm[23:13])
      + conv_u2u_1_11(cvt_14_FpMantDecShiftRight_23U_8U_10U_carry_and_3_nl);
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_14_sva = nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_14_sva[10:0];
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_14_sva = (chn_idata_data_sva_1_443_415_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_guard_mask_14_sva[22:0]);
  assign nl_cvt_14_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl = (FpMantDecShiftRight_23U_8U_10U_guard_mask_14_sva[22:0])
      + 23'b11111111111111111111111;
  assign cvt_14_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl = nl_cvt_14_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_14_sva = (chn_idata_data_sva_1_443_415_1[23:1])
      & (cvt_14_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl);
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_14_sva = (chn_idata_data_sva_1_443_415_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_least_mask_14_sva[22:0]);
  assign cvt_15_FpMantDecShiftRight_23U_8U_10U_carry_and_3_nl = ((FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_15_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_guard_mask_15_sva[23])) & ((FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_15_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_15_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_mask_15_sva[23]));
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_15_sva = (cvt_15_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_3_itm[23:13])
      + conv_u2u_1_11(cvt_15_FpMantDecShiftRight_23U_8U_10U_carry_and_3_nl);
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_15_sva = nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_15_sva[10:0];
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_15_sva = (chn_idata_data_sva_1_475_447_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_guard_mask_15_sva[22:0]);
  assign nl_cvt_15_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl = (FpMantDecShiftRight_23U_8U_10U_guard_mask_15_sva[22:0])
      + 23'b11111111111111111111111;
  assign cvt_15_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl = nl_cvt_15_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_15_sva = (chn_idata_data_sva_1_475_447_1[23:1])
      & (cvt_15_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_3_nl);
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_15_sva = (chn_idata_data_sva_1_475_447_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_least_mask_15_sva[22:0]);
  assign cvt_16_FpMantDecShiftRight_23U_8U_10U_carry_and_4_nl = ((FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_guard_mask_sva[23])) & ((FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_sva!=23'b00000000000000000000000)
      | (FpMantDecShiftRight_23U_8U_10U_least_mask_sva[23]));
  assign nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva = (cvt_16_FpMantDecShiftRight_23U_8U_10U_i_mant_s_rshift_4_itm[23:13])
      + conv_u2u_1_11(cvt_16_FpMantDecShiftRight_23U_8U_10U_carry_and_4_nl);
  assign FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva = nl_FpMantDecShiftRight_23U_8U_10U_o_mant_sum_sva[10:0];
  assign FpMantDecShiftRight_23U_8U_10U_guard_bits_22_0_sva = (chn_idata_data_sva_1_507_479_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_guard_mask_sva[22:0]);
  assign nl_cvt_16_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_4_nl = (FpMantDecShiftRight_23U_8U_10U_guard_mask_sva[22:0])
      + 23'b11111111111111111111111;
  assign cvt_16_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_4_nl = nl_cvt_16_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_4_nl[22:0];
  assign FpMantDecShiftRight_23U_8U_10U_stick_bits_22_0_sva = (chn_idata_data_sva_1_507_479_1[23:1])
      & (cvt_16_FpMantDecShiftRight_23U_8U_10U_stick_mask_acc_4_nl);
  assign FpMantDecShiftRight_23U_8U_10U_least_bits_22_0_sva = (chn_idata_data_sva_1_507_479_1[23:1])
      & (FpMantDecShiftRight_23U_8U_10U_least_mask_sva[22:0]);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_2
      & cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_4_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_15_ssc
      = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_15_tmp | nand_133_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_31_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_15_tmp
      & (~ nand_133_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_15_tmp = cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_2
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_15_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_2
      & cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_14_ssc
      = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_14_tmp | nand_135_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_29_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_14_tmp
      & (~ nand_135_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_14_tmp = cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_14_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_2
      & cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_13_ssc
      = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_13_tmp | nand_137_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_27_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_13_tmp
      & (~ nand_137_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_13_tmp = cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_13_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_2
      & cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_12_ssc
      = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_12_tmp | nand_139_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_25_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_12_tmp
      & (~ nand_139_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_12_tmp = cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_12_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_2
      & cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_11_ssc
      = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_11_tmp | nand_141_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_23_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_11_tmp
      & (~ nand_141_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_11_tmp = cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_11_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_2
      & cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_10_ssc
      = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_10_tmp | nand_143_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_21_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_10_tmp
      & (~ nand_143_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_10_tmp = cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_10_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_2
      & cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_9_ssc
      = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_9_tmp | nand_145_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_19_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_9_tmp
      & (~ nand_145_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_9_tmp = cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_9_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_2
      & cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_8_ssc
      = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_8_tmp | nand_147_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_17_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_8_tmp
      & (~ nand_147_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_8_tmp = cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_8_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_2
      & cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_7_ssc
      = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_7_tmp | nand_149_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_15_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_7_tmp
      & (~ nand_149_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_7_tmp = cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_7_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_2
      & cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_6_ssc
      = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_6_tmp | nand_151_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_13_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_6_tmp
      & (~ nand_151_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_6_tmp = cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_6_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_2
      & cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_5_ssc
      = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_5_tmp | nand_153_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_11_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_5_tmp
      & (~ nand_153_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_5_tmp = cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_5_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_2
      & cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_4_ssc
      = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_4_tmp | nand_156_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_9_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_4_tmp
      & (~ nand_156_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_4_tmp = cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_4_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_2
      & cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_3_ssc
      = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_3_tmp | nand_158_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_7_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_3_tmp
      & (~ nand_158_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_3_tmp = cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_3_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_2
      & cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_2_ssc
      = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_2_tmp | nand_160_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_5_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_2_tmp
      & (~ nand_160_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_2_tmp = cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_2_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_2
      & cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_1_ssc
      = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_1_tmp | nand_162_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_3_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_1_tmp
      & (~ nand_162_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_1_tmp = cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_2);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_is_zero_1_lpi_1_dfm = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_2
      & cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_2;
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_FpWidthDec_8U_23U_5U_10U_1U_1U_nor_ssc =
      ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_tmp | nand_164_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_and_1_m1c = FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_tmp
      & (~ nand_164_cse);
  assign FpWidthDec_8U_23U_5U_10U_1U_1U_else_and_tmp = cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_2
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_2);
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_1_sva = conv_u2u_16_17({(~
      IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_mx0w0) , (~ IntShiftRightSat_49U_6U_17U_o_0_1_sva_mx0w0)})
      + 17'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_1_sva = nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_1_sva[16:0];
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_2_sva = conv_u2u_16_17({(~
      IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_mx0w0) , (~ IntShiftRightSat_49U_6U_17U_o_0_2_sva_mx0w0)})
      + 17'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_2_sva = nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_2_sva[16:0];
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_3_sva = conv_u2u_16_17({(~
      IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_mx0w0) , (~ IntShiftRightSat_49U_6U_17U_o_0_3_sva_mx0w0)})
      + 17'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_3_sva = nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_3_sva[16:0];
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_4_sva = conv_u2u_16_17({(~
      IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_mx0w0) , (~ IntShiftRightSat_49U_6U_17U_o_0_4_sva_mx0w0)})
      + 17'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_4_sva = nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_4_sva[16:0];
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_5_sva = conv_u2u_16_17({(~
      IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_mx0w0) , (~ IntShiftRightSat_49U_6U_17U_o_0_5_sva_mx0w0)})
      + 17'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_5_sva = nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_5_sva[16:0];
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_6_sva = conv_u2u_16_17({(~
      IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_mx0w0) , (~ IntShiftRightSat_49U_6U_17U_o_0_6_sva_mx0w0)})
      + 17'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_6_sva = nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_6_sva[16:0];
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_7_sva = conv_u2u_16_17({(~
      IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_mx0w0) , (~ IntShiftRightSat_49U_6U_17U_o_0_7_sva_mx0w0)})
      + 17'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_7_sva = nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_7_sva[16:0];
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_8_sva = conv_u2u_16_17({(~
      IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_mx0w0) , (~ IntShiftRightSat_49U_6U_17U_o_0_8_sva_mx0w0)})
      + 17'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_8_sva = nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_8_sva[16:0];
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_9_sva = conv_u2u_16_17({(~
      IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_mx0w0) , (~ IntShiftRightSat_49U_6U_17U_o_0_9_sva_mx0w0)})
      + 17'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_9_sva = nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_9_sva[16:0];
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_10_sva = conv_u2u_16_17({(~
      IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_mx0w0) , (~ IntShiftRightSat_49U_6U_17U_o_0_10_sva_mx0w0)})
      + 17'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_10_sva = nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_10_sva[16:0];
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_11_sva = conv_u2u_16_17({(~
      IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_mx0w0) , (~ IntShiftRightSat_49U_6U_17U_o_0_11_sva_mx0w0)})
      + 17'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_11_sva = nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_11_sva[16:0];
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_12_sva = conv_u2u_16_17({(~
      IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_mx0w0) , (~ IntShiftRightSat_49U_6U_17U_o_0_12_sva_mx0w0)})
      + 17'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_12_sva = nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_12_sva[16:0];
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_13_sva = conv_u2u_16_17({(~
      IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_mx0w0) , (~ IntShiftRightSat_49U_6U_17U_o_0_13_sva_mx0w0)})
      + 17'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_13_sva = nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_13_sva[16:0];
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_14_sva = conv_u2u_16_17({(~
      IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_mx0w0) , (~ IntShiftRightSat_49U_6U_17U_o_0_14_sva_mx0w0)})
      + 17'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_14_sva = nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_14_sva[16:0];
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_15_sva = conv_u2u_16_17({(~
      IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_mx0w0) , (~ IntShiftRightSat_49U_6U_17U_o_0_15_sva_mx0w0)})
      + 17'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_15_sva = nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_15_sva[16:0];
  assign nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_sva = conv_u2u_16_17({(~
      IntShiftRightSat_49U_6U_17U_o_15_1_sva_mx0w0) , (~ IntShiftRightSat_49U_6U_17U_o_0_sva_mx0w0)})
      + 17'b1;
  assign FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_sva = nl_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_sva[16:0];
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_m1c = ~(cvt_1_FpFloatToInt_16U_5U_10U_if_acc_itm_11_1
      | IsNaN_5U_10U_land_1_lpi_1_dfm_mx0w0);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_1_m1c = ~(cvt_2_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1
      | IsNaN_5U_10U_land_2_lpi_1_dfm_mx0w0);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_2_m1c = ~(cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1
      | IsNaN_5U_10U_land_3_lpi_1_dfm_4);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_3_m1c = ~(cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1
      | IsNaN_5U_10U_land_4_lpi_1_dfm_4);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_4_m1c = ~(cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1
      | IsNaN_5U_10U_land_5_lpi_1_dfm_4);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_5_m1c = ~(cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1
      | IsNaN_5U_10U_land_6_lpi_1_dfm_4);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_6_m1c = ~(cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1
      | IsNaN_5U_10U_land_7_lpi_1_dfm_5);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_7_m1c = ~(cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1
      | IsNaN_5U_10U_land_8_lpi_1_dfm_4);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_8_m1c = ~(cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1
      | IsNaN_5U_10U_land_9_lpi_1_dfm_4);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_9_m1c = ~(cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1
      | IsNaN_5U_10U_land_10_lpi_1_dfm_4);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_10_m1c = ~(cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1
      | IsNaN_5U_10U_land_11_lpi_1_dfm_4);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_11_m1c = ~(cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1
      | IsNaN_5U_10U_land_12_lpi_1_dfm_4);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_12_m1c = ~(cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1
      | IsNaN_5U_10U_land_13_lpi_1_dfm_4);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_13_m1c = ~(cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1
      | IsNaN_5U_10U_land_14_lpi_1_dfm_5);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_14_m1c = ~(cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1
      | IsNaN_5U_10U_land_15_lpi_1_dfm_mx0w0);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_15_m1c = ~(cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_itm_11_1
      | IsNaN_5U_10U_land_lpi_1_dfm_4);
  assign nl_cvt_1_IntSaturation_17U_16U_else_if_acc_nl = conv_s2u_2_3({IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0
      , (IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_mx0w0[14])}) + 3'b1;
  assign cvt_1_IntSaturation_17U_16U_else_if_acc_nl = nl_cvt_1_IntSaturation_17U_16U_else_if_acc_nl[2:0];
  assign cvt_1_IntSaturation_17U_16U_else_if_acc_itm_2_1 = readslicef_3_1_2((cvt_1_IntSaturation_17U_16U_else_if_acc_nl));
  assign nl_cvt_2_IntSaturation_17U_16U_else_if_acc_1_nl = conv_s2u_2_3({IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0
      , (IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_mx0w0[14])}) + 3'b1;
  assign cvt_2_IntSaturation_17U_16U_else_if_acc_1_nl = nl_cvt_2_IntSaturation_17U_16U_else_if_acc_1_nl[2:0];
  assign cvt_2_IntSaturation_17U_16U_else_if_acc_1_itm_2_1 = readslicef_3_1_2((cvt_2_IntSaturation_17U_16U_else_if_acc_1_nl));
  assign nl_cvt_3_IntSaturation_17U_16U_else_if_acc_1_nl = conv_s2u_2_3({IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0
      , (IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_mx0w0[14])}) + 3'b1;
  assign cvt_3_IntSaturation_17U_16U_else_if_acc_1_nl = nl_cvt_3_IntSaturation_17U_16U_else_if_acc_1_nl[2:0];
  assign cvt_3_IntSaturation_17U_16U_else_if_acc_1_itm_2_1 = readslicef_3_1_2((cvt_3_IntSaturation_17U_16U_else_if_acc_1_nl));
  assign nl_cvt_4_IntSaturation_17U_16U_else_if_acc_2_nl = conv_s2u_2_3({IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0
      , (IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_mx0w0[14])}) + 3'b1;
  assign cvt_4_IntSaturation_17U_16U_else_if_acc_2_nl = nl_cvt_4_IntSaturation_17U_16U_else_if_acc_2_nl[2:0];
  assign cvt_4_IntSaturation_17U_16U_else_if_acc_2_itm_2_1 = readslicef_3_1_2((cvt_4_IntSaturation_17U_16U_else_if_acc_2_nl));
  assign nl_cvt_5_IntSaturation_17U_16U_else_if_acc_1_nl = conv_s2u_2_3({IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0
      , (IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_mx0w0[14])}) + 3'b1;
  assign cvt_5_IntSaturation_17U_16U_else_if_acc_1_nl = nl_cvt_5_IntSaturation_17U_16U_else_if_acc_1_nl[2:0];
  assign cvt_5_IntSaturation_17U_16U_else_if_acc_1_itm_2_1 = readslicef_3_1_2((cvt_5_IntSaturation_17U_16U_else_if_acc_1_nl));
  assign nl_cvt_6_IntSaturation_17U_16U_else_if_acc_2_nl = conv_s2u_2_3({IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0
      , (IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_mx0w0[14])}) + 3'b1;
  assign cvt_6_IntSaturation_17U_16U_else_if_acc_2_nl = nl_cvt_6_IntSaturation_17U_16U_else_if_acc_2_nl[2:0];
  assign cvt_6_IntSaturation_17U_16U_else_if_acc_2_itm_2_1 = readslicef_3_1_2((cvt_6_IntSaturation_17U_16U_else_if_acc_2_nl));
  assign nl_cvt_7_IntSaturation_17U_16U_else_if_acc_2_nl = conv_s2u_2_3({IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0
      , (IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_mx0w0[14])}) + 3'b1;
  assign cvt_7_IntSaturation_17U_16U_else_if_acc_2_nl = nl_cvt_7_IntSaturation_17U_16U_else_if_acc_2_nl[2:0];
  assign cvt_7_IntSaturation_17U_16U_else_if_acc_2_itm_2_1 = readslicef_3_1_2((cvt_7_IntSaturation_17U_16U_else_if_acc_2_nl));
  assign nl_cvt_8_IntSaturation_17U_16U_else_if_acc_3_nl = conv_s2u_2_3({IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0
      , (IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_mx0w0[14])}) + 3'b1;
  assign cvt_8_IntSaturation_17U_16U_else_if_acc_3_nl = nl_cvt_8_IntSaturation_17U_16U_else_if_acc_3_nl[2:0];
  assign cvt_8_IntSaturation_17U_16U_else_if_acc_3_itm_2_1 = readslicef_3_1_2((cvt_8_IntSaturation_17U_16U_else_if_acc_3_nl));
  assign nl_cvt_9_IntSaturation_17U_16U_else_if_acc_1_nl = conv_s2u_2_3({IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0
      , (IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_mx0w0[14])}) + 3'b1;
  assign cvt_9_IntSaturation_17U_16U_else_if_acc_1_nl = nl_cvt_9_IntSaturation_17U_16U_else_if_acc_1_nl[2:0];
  assign cvt_9_IntSaturation_17U_16U_else_if_acc_1_itm_2_1 = readslicef_3_1_2((cvt_9_IntSaturation_17U_16U_else_if_acc_1_nl));
  assign nl_cvt_10_IntSaturation_17U_16U_else_if_acc_2_nl = conv_s2u_2_3({IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0
      , (IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_mx0w0[14])}) + 3'b1;
  assign cvt_10_IntSaturation_17U_16U_else_if_acc_2_nl = nl_cvt_10_IntSaturation_17U_16U_else_if_acc_2_nl[2:0];
  assign cvt_10_IntSaturation_17U_16U_else_if_acc_2_itm_2_1 = readslicef_3_1_2((cvt_10_IntSaturation_17U_16U_else_if_acc_2_nl));
  assign nl_cvt_11_IntSaturation_17U_16U_else_if_acc_2_nl = conv_s2u_2_3({IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0
      , (IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_mx0w0[14])}) + 3'b1;
  assign cvt_11_IntSaturation_17U_16U_else_if_acc_2_nl = nl_cvt_11_IntSaturation_17U_16U_else_if_acc_2_nl[2:0];
  assign cvt_11_IntSaturation_17U_16U_else_if_acc_2_itm_2_1 = readslicef_3_1_2((cvt_11_IntSaturation_17U_16U_else_if_acc_2_nl));
  assign nl_cvt_12_IntSaturation_17U_16U_else_if_acc_3_nl = conv_s2u_2_3({IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0
      , (IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_mx0w0[14])}) + 3'b1;
  assign cvt_12_IntSaturation_17U_16U_else_if_acc_3_nl = nl_cvt_12_IntSaturation_17U_16U_else_if_acc_3_nl[2:0];
  assign cvt_12_IntSaturation_17U_16U_else_if_acc_3_itm_2_1 = readslicef_3_1_2((cvt_12_IntSaturation_17U_16U_else_if_acc_3_nl));
  assign nl_cvt_13_IntSaturation_17U_16U_else_if_acc_2_nl = conv_s2u_2_3({IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0
      , (IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_mx0w0[14])}) + 3'b1;
  assign cvt_13_IntSaturation_17U_16U_else_if_acc_2_nl = nl_cvt_13_IntSaturation_17U_16U_else_if_acc_2_nl[2:0];
  assign cvt_13_IntSaturation_17U_16U_else_if_acc_2_itm_2_1 = readslicef_3_1_2((cvt_13_IntSaturation_17U_16U_else_if_acc_2_nl));
  assign nl_cvt_15_IntSaturation_17U_16U_else_if_acc_3_nl = conv_s2u_2_3({IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0
      , (IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_mx0w0[14])}) + 3'b1;
  assign cvt_15_IntSaturation_17U_16U_else_if_acc_3_nl = nl_cvt_15_IntSaturation_17U_16U_else_if_acc_3_nl[2:0];
  assign cvt_15_IntSaturation_17U_16U_else_if_acc_3_itm_2_1 = readslicef_3_1_2((cvt_15_IntSaturation_17U_16U_else_if_acc_3_nl));
  assign nl_cvt_16_IntSaturation_17U_16U_else_if_acc_4_nl = conv_s2u_2_3({IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0
      , (IntShiftRightSat_49U_6U_17U_o_15_1_sva_mx0w0[14])}) + 3'b1;
  assign cvt_16_IntSaturation_17U_16U_else_if_acc_4_nl = nl_cvt_16_IntSaturation_17U_16U_else_if_acc_4_nl[2:0];
  assign cvt_16_IntSaturation_17U_16U_else_if_acc_4_itm_2_1 = readslicef_3_1_2((cvt_16_IntSaturation_17U_16U_else_if_acc_4_nl));
  assign nl_cvt_14_IntSaturation_17U_16U_else_if_acc_3_nl = conv_s2u_2_3({IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0
      , (IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_mx0w0[14])}) + 3'b1;
  assign cvt_14_IntSaturation_17U_16U_else_if_acc_3_nl = nl_cvt_14_IntSaturation_17U_16U_else_if_acc_3_nl[2:0];
  assign cvt_14_IntSaturation_17U_16U_else_if_acc_3_itm_2_1 = readslicef_3_1_2((cvt_14_IntSaturation_17U_16U_else_if_acc_3_nl));
  assign cvt_asn_319 = ~(cvt_if_unequal_tmp | cfg_mode_eql_1_sva_6 | cvt_unequal_tmp_21);
  assign cvt_asn_321 = cvt_if_unequal_tmp & (~ cfg_mode_eql_1_sva_6) & (~ cvt_unequal_tmp_21);
  assign cvt_asn_323 = cvt_else_nor_dfs & (~ cfg_mode_eql_1_sva_6) & cvt_unequal_tmp_21;
  assign cvt_asn_327 = cvt_else_equal_tmp_1 & (~ cfg_mode_eql_1_sva_6) & cvt_unequal_tmp_21;
  assign cvt_asn_329 = cvt_else_nor_dfs_1_mx1 & (~ cfg_mode_eql_1_sva_6) & cvt_unequal_tmp_21;
  assign cvt_asn_333 = cvt_else_equal_tmp_4_mx1 & (~ cfg_mode_eql_1_sva_6) & cvt_unequal_tmp_21;
  assign cvt_asn_335 = cvt_else_nor_dfs_3_mx1 & (~ cfg_mode_eql_1_sva_6) & cvt_unequal_tmp_21;
  assign cvt_asn_339 = cvt_else_equal_tmp_10_mx0 & (~ cfg_mode_eql_1_sva_6) & cvt_unequal_tmp_21;
  assign cvt_asn_341 = cvt_else_nor_dfs_15_mx1 & cvt_unequal_tmp_21 & (~ cfg_mode_eql_1_sva_6);
  assign cvt_asn_345 = cvt_else_equal_tmp_46_mx1 & cvt_unequal_tmp_21 & (~ cfg_mode_eql_1_sva_6);
  assign cvt_asn_347 = cvt_else_nor_dfs_14_mx1 & (~ cfg_mode_eql_1_sva_6) & cvt_unequal_tmp_21;
  assign cvt_asn_351 = cvt_else_equal_tmp_43_mx0 & (~ cfg_mode_eql_1_sva_6) & cvt_unequal_tmp_21;
  assign cvt_asn_353 = cvt_else_nor_dfs_5_mx1 & (~ cfg_mode_eql_1_sva_6) & cvt_unequal_tmp_21;
  assign cvt_asn_357 = cvt_else_equal_tmp_16_mx1 & (~ cfg_mode_eql_1_sva_6) & cvt_unequal_tmp_21;
  assign cvt_asn_359 = cvt_else_nor_dfs_13_mx1 & (~ cfg_mode_eql_1_sva_6) & cvt_unequal_tmp_21;
  assign cvt_asn_363 = cvt_else_equal_tmp_40_mx1 & (~ cfg_mode_eql_1_sva_6) & cvt_unequal_tmp_21;
  assign cvt_asn_365 = cvt_else_nor_dfs_6_mx1 & (~ cfg_mode_eql_1_sva_6) & cvt_unequal_tmp_21;
  assign cvt_asn_369 = cvt_else_equal_tmp_19_mx0 & (~ cfg_mode_eql_1_sva_6) & cvt_unequal_tmp_21;
  assign cvt_asn_371 = cvt_else_nor_dfs_9_mx1 & (~ cfg_mode_eql_1_sva_6) & cvt_unequal_tmp_21;
  assign cvt_asn_375 = cvt_else_equal_tmp_37_mx0 & (~ cfg_mode_eql_1_sva_6) & cvt_unequal_tmp_21;
  assign cvt_asn_377 = cvt_else_nor_dfs_7_mx1 & cvt_and_147_m1c;
  assign cvt_asn_381 = cvt_else_equal_tmp_22_mx1 & cvt_and_147_m1c;
  assign cvt_asn_383 = cvt_else_nor_dfs_11_mx1 & (~ cfg_mode_eql_1_sva_6) & cvt_unequal_tmp_21;
  assign cvt_asn_387 = cvt_else_equal_tmp_34_mx1 & (~ cfg_mode_eql_1_sva_6) & cvt_unequal_tmp_21;
  assign cvt_asn_389 = cvt_else_nor_dfs_10_mx1 & (~ cfg_mode_eql_1_sva_6) & cvt_unequal_tmp_21;
  assign cvt_asn_393 = cvt_else_equal_tmp_31_mx0 & (~ cfg_mode_eql_1_sva_6) & cvt_unequal_tmp_21;
  assign cvt_asn_399 = cvt_else_equal_tmp_28_mx1 & (~ cfg_mode_eql_1_sva_6) & cvt_unequal_tmp_21;
  assign and_dcpl_3 = (cfg_proc_precision_1_sva_st_64==2'b10);
  assign and_dcpl_4 = and_dcpl_3 & or_5189_cse;
  assign and_dcpl_70 = chn_in_rsci_bawt & (cfg_proc_precision_rsci_d[1]);
  assign and_dcpl_71 = and_dcpl_70 & (~ (cfg_proc_precision_rsci_d[0]));
  assign and_dcpl_73 = chn_out_rsci_bawt & reg_chn_out_rsci_ld_core_psct_cse;
  assign and_dcpl_75 = or_5189_cse & (~ (cfg_out_precision_rsci_d[1]));
  assign and_dcpl_77 = or_4524_cse & chn_in_rsci_bawt & (cfg_out_precision_rsci_d[0]);
  assign and_dcpl_80 = (~ (cfg_out_precision_rsci_d[1])) & chn_out_rsci_bawt & reg_chn_out_rsci_ld_core_psct_cse;
  assign and_dcpl_83 = or_4524_cse & chn_in_rsci_bawt & (~ (cfg_out_precision_rsci_d[0]));
  assign or_tmp_19 = (cfg_proc_precision_rsci_d[0]) | (~ and_dcpl_70);
  assign or_23_nl = (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_tmp_6 = MUX_s_1_2_2((or_23_nl), or_tmp_19, or_5189_cse);
  assign or_tmp_24 = nor_2040_cse | (cfg_proc_precision_rsci_d[0]) | (~ and_dcpl_70);
  assign or_86_nl = (~ cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_st_2
      | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_tmp_39 = MUX_s_1_2_2((or_86_nl), or_tmp_19, or_5189_cse);
  assign mux_109_nl = MUX_s_1_2_2(or_186_cse, (~ or_4550_cse), reg_cfg_proc_precision_1_sva_st_40_cse[1]);
  assign mux_110_cse = MUX_s_1_2_2((mux_109_nl), or_186_cse, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign and_tmp_8 = main_stage_v_1 & mux_110_cse;
  assign and_tmp_11 = main_stage_v_1 & or_4550_cse;
  assign mux_tmp_114 = MUX_s_1_2_2(and_tmp_11, and_2186_cse, or_5189_cse);
  assign and_tmp_12 = or_183_cse_1 & or_4550_cse;
  assign nor_2056_nl = ~((reg_cfg_proc_precision_1_sva_st_40_cse[1]) | (~ and_tmp_12));
  assign mux_tmp_117 = MUX_s_1_2_2((nor_2056_nl), and_tmp_12, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign and_tmp_16 = main_stage_v_1 & mux_tmp_117;
  assign or_tmp_213 = (cfg_out_precision_rsci_d!=2'b10) | (~ and_2186_cse);
  assign nor_2055_nl = ~((reg_cfg_proc_precision_1_sva_st_40_cse[1]) | and_dcpl_3);
  assign mux_tmp_120 = MUX_s_1_2_2((nor_2055_nl), or_4550_cse, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign not_tmp_119 = ~((cfg_out_precision_1_sva_st_154[1]) & main_stage_v_1 & mux_tmp_120);
  assign or_tmp_218 = (cfg_out_precision_1_sva_st_154[0]) | not_tmp_119;
  assign and_tmp_18 = main_stage_v_1 & mux_tmp_120;
  assign mux_tmp_122 = MUX_s_1_2_2(and_tmp_18, and_2186_cse, or_5189_cse);
  assign nor_2054_nl = ~((reg_cfg_proc_precision_1_sva_st_40_cse[1]) | (~ mux_tmp_120));
  assign mux_tmp_123 = MUX_s_1_2_2((nor_2054_nl), mux_tmp_120, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign and_tmp_19 = main_stage_v_1 & mux_tmp_123;
  assign nor_2052_nl = ~((reg_cfg_proc_precision_1_sva_st_40_cse[1]) | (~ and_tmp_19));
  assign mux_tmp_129 = MUX_s_1_2_2((nor_2052_nl), and_tmp_19, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign nor_2050_nl = ~((reg_cfg_proc_precision_1_sva_st_40_cse[1]) | (~ mux_tmp_117));
  assign mux_148_nl = MUX_s_1_2_2((nor_2050_nl), mux_tmp_117, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign and_tmp_33 = main_stage_v_1 & (mux_148_nl);
  assign nor_2049_nl = ~((reg_cfg_proc_precision_1_sva_st_40_cse[1]) | (~ and_tmp_33));
  assign mux_tmp_151 = MUX_s_1_2_2((nor_2049_nl), and_tmp_33, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign mux_tmp_161 = MUX_s_1_2_2(main_stage_v_2, main_stage_v_1, or_5189_cse);
  assign or_tmp_306 = (~ main_stage_v_2) | (cfg_proc_precision_1_sva_st_65!=2'b10);
  assign nor_2029_nl = ~((cfg_proc_precision_1_sva_st_64[1]) | (~ cfg_mode_eql_1_sva_4));
  assign mux_188_nl = MUX_s_1_2_2((nor_2029_nl), cfg_mode_eql_1_sva_4, cfg_proc_precision_1_sva_st_64[0]);
  assign nand_nl = ~(main_stage_v_1 & (~ (mux_188_nl)));
  assign or_378_nl = (~ main_stage_v_1) | cfg_mode_eql_1_sva_4;
  assign nor_48_nl = ~((cfg_out_precision_1_sva_st_154!=2'b01));
  assign mux_tmp_189 = MUX_s_1_2_2((or_378_nl), (nand_nl), nor_48_nl);
  assign or_tmp_378 = (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b01)
      | (cfg_proc_precision_1_sva_st_65!=2'b10);
  assign nor_2027_nl = ~((cfg_proc_precision_1_sva_st_89[1]) | (~ main_stage_v_2));
  assign mux_tmp_199 = MUX_s_1_2_2((nor_2027_nl), main_stage_v_2, cfg_proc_precision_1_sva_st_89[0]);
  assign nor_2028_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ mux_tmp_199));
  assign mux_tmp_200 = MUX_s_1_2_2((nor_2028_nl), mux_tmp_199, cfg_proc_precision_1_sva_st_101[0]);
  assign or_tmp_389 = (cfg_proc_precision_1_sva_st_89[0]) | (~((cfg_proc_precision_1_sva_st_89[1])
      & or_4862_cse));
  assign nor_2022_nl = ~((cfg_proc_precision_1_sva_st_64[1]) | (~ main_stage_v_1));
  assign mux_tmp_236 = MUX_s_1_2_2((nor_2022_nl), main_stage_v_1, cfg_proc_precision_1_sva_st_64[0]);
  assign nor_2021_nl = ~((cfg_proc_precision_1_sva_st_65[1]) | (~ main_stage_v_2));
  assign mux_tmp_239 = MUX_s_1_2_2((nor_2021_nl), main_stage_v_2, cfg_proc_precision_1_sva_st_65[0]);
  assign or_429_nl = cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_tmp
      | (cfg_out_precision_1_sva_st_154!=2'b10) | (~ and_tmp_11);
  assign or_431_nl = (~ main_stage_v_2) | cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_svs_st_2
      | (~ or_4862_cse);
  assign mux_244_nl = MUX_s_1_2_2((or_431_nl), (or_429_nl), or_5189_cse);
  assign or_434_nl = nor_2040_cse | cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_tmp
      | (cfg_out_precision_1_sva_st_154!=2'b10) | (~ and_tmp_11);
  assign mux_tmp_245 = MUX_s_1_2_2((or_434_nl), (mux_244_nl), nor_57_cse);
  assign and_tmp_50 = or_4714_cse & or_4862_cse;
  assign and_tmp_52 = main_stage_v_2 & (IntShiftRightSat_49U_6U_17U_lor_3_lpi_1_dfm
      | cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2)
      & and_tmp_50;
  assign or_448_nl = (cfg_proc_precision_1_sva_st_64[0]) | (~((cfg_proc_precision_1_sva_st_64[1])
      & or_513_cse));
  assign mux_tmp_249 = MUX_s_1_2_2((~ or_513_cse), (or_448_nl), or_183_cse_1);
  assign mux_250_nl = MUX_s_1_2_2((~ or_513_cse), mux_tmp_249, cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp);
  assign and_152_nl = main_stage_v_1 & (mux_250_nl);
  assign and_153_nl = main_stage_v_1 & mux_tmp_249;
  assign or_445_nl = (cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp
      & (cfg_out_precision_1_sva_st_154[1])) | (cfg_out_precision_1_sva_st_154[0]);
  assign mux_tmp_251 = MUX_s_1_2_2((and_153_nl), (and_152_nl), or_445_nl);
  assign mux_252_nl = MUX_s_1_2_2(main_stage_v_2, and_tmp_52, or_451_cse);
  assign mux_tmp_253 = MUX_s_1_2_2((mux_252_nl), mux_tmp_251, or_5189_cse);
  assign nor_2015_nl = ~((reg_cfg_proc_precision_1_sva_st_40_cse[1]) | (~ mux_tmp_236));
  assign mux_tmp_259 = MUX_s_1_2_2((nor_2015_nl), mux_tmp_236, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign nor_2013_nl = ~((cfg_proc_precision_1_sva_st_89[1]) | (~ mux_tmp_239));
  assign mux_tmp_263 = MUX_s_1_2_2((nor_2013_nl), mux_tmp_239, cfg_proc_precision_1_sva_st_89[0]);
  assign nor_2007_nl = ~((~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp | (~ mux_344_cse));
  assign nor_2009_nl = ~(nor_2219_cse | (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 |
      nor_50_cse);
  assign not_tmp_249 = MUX_s_1_2_2((nor_2009_nl), (nor_2007_nl), or_5189_cse);
  assign nor_1995_nl = ~((~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp | (~ mux_344_cse));
  assign nor_1997_nl = ~(nor_2219_cse | (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 |
      nor_50_cse);
  assign not_tmp_269 = MUX_s_1_2_2((nor_1997_nl), (nor_1995_nl), or_5189_cse);
  assign not_tmp_270 = ~((cfg_out_precision_1_sva_st_154[1]) & main_stage_v_1 & and_tmp_12);
  assign or_510_cse = IntShiftRightSat_49U_6U_17U_lor_5_lpi_1_dfm | cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2;
  assign and_tmp_67 = or_510_cse & and_tmp_50;
  assign nor_1988_nl = ~(((cfg_out_precision_1_sva_st_154[1]) & cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp)
      | (cfg_out_precision_1_sva_st_154[0]) | (~ mux_tmp_259));
  assign mux_tmp_294 = MUX_s_1_2_2((nor_1988_nl), mux_tmp_259, cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp);
  assign nor_1987_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ mux_tmp_239));
  assign mux_tmp_298 = MUX_s_1_2_2((nor_1987_nl), mux_tmp_239, cfg_proc_precision_1_sva_st_101[0]);
  assign and_167_nl = or_510_cse & mux_tmp_298;
  assign or_520_nl = ((cfg_out_precision_1_sva_st_149[1]) & FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_3)
      | (cfg_out_precision_1_sva_st_149[0]);
  assign mux_tmp_299 = MUX_s_1_2_2(mux_tmp_298, (and_167_nl), or_520_nl);
  assign nor_1983_nl = ~((reg_cfg_proc_precision_1_sva_st_40_cse[1]) | (~ mux_tmp_259));
  assign mux_tmp_305 = MUX_s_1_2_2((nor_1983_nl), mux_tmp_259, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign or_tmp_533 = (~ cvt_unequal_tmp_20) | cfg_mode_eql_1_sva_5 | (cfg_out_precision_1_sva_st_113!=2'b00)
      | (~ main_stage_v_2);
  assign mux_308_nl = MUX_s_1_2_2(main_stage_v_2, (~ or_tmp_533), cfg_proc_precision_1_sva_st_65[1]);
  assign mux_tmp_309 = MUX_s_1_2_2((mux_308_nl), main_stage_v_2, cfg_proc_precision_1_sva_st_65[0]);
  assign mux_310_nl = MUX_s_1_2_2(mux_tmp_309, (~ or_tmp_533), cfg_proc_precision_1_sva_st_101[1]);
  assign mux_tmp_311 = MUX_s_1_2_2((mux_310_nl), mux_tmp_309, cfg_proc_precision_1_sva_st_101[0]);
  assign mux_312_nl = MUX_s_1_2_2((~ or_tmp_533), mux_tmp_311, or_510_cse);
  assign mux_tmp_313 = MUX_s_1_2_2(mux_tmp_311, (mux_312_nl), or_461_cse);
  assign mux_tmp_317 = MUX_s_1_2_2((~ (reg_cfg_proc_precision_1_sva_st_40_cse[1])),
      or_183_cse_1, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign nor_1975_nl = ~((~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp | (~ mux_474_cse));
  assign nor_1977_nl = ~(nor_151_cse | nor_2219_cse | (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_3 | nor_50_cse);
  assign not_tmp_312 = MUX_s_1_2_2((nor_1977_nl), (nor_1975_nl), or_5189_cse);
  assign nor_1974_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ and_tmp_50));
  assign mux_tmp_321 = MUX_s_1_2_2((nor_1974_nl), and_tmp_50, cfg_proc_precision_1_sva_st_101[0]);
  assign and_tmp_71 = main_stage_v_1 & cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp
      & mux_tmp_120;
  assign nor_1964_nl = ~((~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp | (~ mux_344_cse));
  assign nor_1966_nl = ~(nor_2219_cse | (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 |
      nor_50_cse);
  assign not_tmp_336 = MUX_s_1_2_2((nor_1966_nl), (nor_1964_nl), or_5189_cse);
  assign nor_1959_nl = ~((cfg_proc_precision_1_sva_st_89[1]) | (~ or_400_cse_1));
  assign mux_tmp_345 = MUX_s_1_2_2((nor_1959_nl), or_400_cse_1, cfg_proc_precision_1_sva_st_89[0]);
  assign nor_1955_nl = ~(((cfg_out_precision_1_sva_st_154[1]) & cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp)
      | (cfg_out_precision_1_sva_st_154[0]) | (~ mux_tmp_259));
  assign mux_tmp_351 = MUX_s_1_2_2((nor_1955_nl), mux_tmp_259, cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp);
  assign or_600_cse = IntShiftRightSat_49U_6U_17U_lor_7_lpi_1_dfm | cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2;
  assign and_176_nl = or_600_cse & mux_tmp_298;
  assign or_599_nl = ((cfg_out_precision_1_sva_st_149[1]) & FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_3)
      | (cfg_out_precision_1_sva_st_149[0]);
  assign mux_tmp_356 = MUX_s_1_2_2(mux_tmp_298, (and_176_nl), or_599_nl);
  assign mux_369_nl = MUX_s_1_2_2((~ or_tmp_533), mux_tmp_311, or_600_cse);
  assign mux_tmp_370 = MUX_s_1_2_2(mux_tmp_311, (mux_369_nl), or_461_cse);
  assign nor_1942_nl = ~((~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp | (~ mux_344_cse));
  assign nor_1944_nl = ~(nor_151_cse | nor_2219_cse | (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_3 | nor_50_cse);
  assign not_tmp_388 = MUX_s_1_2_2((nor_1944_nl), (nor_1942_nl), or_5189_cse);
  assign and_tmp_79 = or_400_cse_1 & mux_1126_cse;
  assign nor_1935_nl = ~(((cfg_out_precision_1_sva_st_154[1]) & cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp)
      | (cfg_out_precision_1_sva_st_154[0]) | (~ mux_tmp_259));
  assign mux_tmp_386 = MUX_s_1_2_2((nor_1935_nl), mux_tmp_259, cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp);
  assign and_181_nl = or_4536_cse & mux_tmp_298;
  assign or_645_nl = ((cfg_out_precision_1_sva_st_149[1]) & FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_3)
      | (cfg_out_precision_1_sva_st_149[0]);
  assign mux_tmp_391 = MUX_s_1_2_2(mux_tmp_298, (and_181_nl), or_645_nl);
  assign mux_404_nl = MUX_s_1_2_2((~ or_tmp_533), mux_tmp_311, or_4536_cse);
  assign mux_tmp_405 = MUX_s_1_2_2(mux_tmp_311, (mux_404_nl), or_461_cse);
  assign nor_1922_nl = ~((~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp | (~ mux_344_cse));
  assign nor_1924_nl = ~(nor_151_cse | nor_2219_cse | (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_3 | nor_50_cse);
  assign not_tmp_436 = MUX_s_1_2_2((nor_1924_nl), (nor_1922_nl), or_5189_cse);
  assign mux_tmp_415 = MUX_s_1_2_2((~ (cfg_proc_precision_1_sva_st_101[1])), or_400_cse_1,
      cfg_proc_precision_1_sva_st_101[0]);
  assign nor_1919_nl = ~((cfg_proc_precision_1_sva_st_89[1]) | (~ mux_tmp_415));
  assign mux_tmp_416 = MUX_s_1_2_2((nor_1919_nl), mux_tmp_415, cfg_proc_precision_1_sva_st_89[0]);
  assign nor_1912_nl = ~(((cfg_out_precision_1_sva_st_154[1]) & cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp)
      | (cfg_out_precision_1_sva_st_154[0]) | (~ mux_tmp_259));
  assign mux_tmp_421 = MUX_s_1_2_2((nor_1912_nl), mux_tmp_259, cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp);
  assign nor_1915_nl = ~((reg_cfg_proc_precision_1_sva_st_40_cse[1]) | (~ mux_tmp_421));
  assign mux_tmp_422 = MUX_s_1_2_2((nor_1915_nl), mux_tmp_421, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign and_184_nl = or_4535_cse & mux_tmp_298;
  assign or_690_nl = ((cfg_out_precision_1_sva_st_149[1]) & FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_3)
      | (cfg_out_precision_1_sva_st_149[0]);
  assign mux_tmp_427 = MUX_s_1_2_2(mux_tmp_298, (and_184_nl), or_690_nl);
  assign nor_1911_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ mux_tmp_427));
  assign mux_tmp_428 = MUX_s_1_2_2((nor_1911_nl), mux_tmp_427, cfg_proc_precision_1_sva_st_101[0]);
  assign nor_1906_nl = ~((reg_cfg_proc_precision_1_sva_st_40_cse[1]) | (~ mux_tmp_305));
  assign mux_tmp_435 = MUX_s_1_2_2((nor_1906_nl), mux_tmp_305, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign nor_1901_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ mux_tmp_298));
  assign mux_tmp_440 = MUX_s_1_2_2((nor_1901_nl), mux_tmp_298, cfg_proc_precision_1_sva_st_101[0]);
  assign nor_1902_nl = ~((cfg_proc_precision_1_sva_st_89[1]) | (~ mux_tmp_440));
  assign mux_tmp_441 = MUX_s_1_2_2((nor_1902_nl), mux_tmp_440, cfg_proc_precision_1_sva_st_89[0]);
  assign nor_1892_nl = ~((~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp | (~ mux_344_cse));
  assign nor_1894_nl = ~(nor_151_cse | nor_2219_cse | (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_3 | nor_50_cse);
  assign not_tmp_497 = MUX_s_1_2_2((nor_1894_nl), (nor_1892_nl), or_5189_cse);
  assign and_tmp_93 = main_stage_v_1 & or_183_cse_1 & cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp
      & or_4550_cse;
  assign nor_1891_nl = ~((cfg_proc_precision_1_sva_st_89[1]) | (~ or_4862_cse));
  assign mux_tmp_455 = MUX_s_1_2_2((nor_1891_nl), or_4862_cse, cfg_proc_precision_1_sva_st_89[0]);
  assign and_tmp_94 = main_stage_v_2 & mux_tmp_455;
  assign nor_1882_nl = ~((~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp | (~ mux_344_cse));
  assign nor_1884_nl = ~((~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 |
      (~ mux_1126_cse));
  assign not_tmp_520 = MUX_s_1_2_2((nor_1884_nl), (nor_1882_nl), or_5189_cse);
  assign nor_1872_nl = ~(((cfg_out_precision_1_sva_st_154[1]) & cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp)
      | (cfg_out_precision_1_sva_st_154[0]) | (~ mux_tmp_259));
  assign mux_tmp_481 = MUX_s_1_2_2((nor_1872_nl), mux_tmp_259, cvt_10_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp);
  assign and_2218_nl = IntShiftRightSat_49U_6U_17U_lor_10_lpi_1_dfm & mux_tmp_298;
  assign or_784_nl = ((cfg_out_precision_1_sva_st_149[1]) & FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_3)
      | (cfg_out_precision_1_sva_st_149[0]);
  assign mux_486_nl = MUX_s_1_2_2(mux_tmp_298, (and_2218_nl), or_784_nl);
  assign mux_tmp_487 = MUX_s_1_2_2((mux_486_nl), mux_tmp_298, IntShiftRightSat_49U_6U_17U_lor_11_lpi_1_dfm);
  assign mux_500_nl = MUX_s_1_2_2((~ or_tmp_533), mux_tmp_311, IntShiftRightSat_49U_6U_17U_lor_10_lpi_1_dfm);
  assign or_795_nl = (~((cfg_out_precision_1_sva_st_149!=2'b00))) | IntShiftRightSat_49U_6U_17U_lor_11_lpi_1_dfm;
  assign mux_tmp_502 = MUX_s_1_2_2((mux_500_nl), mux_tmp_311, or_795_nl);
  assign nor_1858_nl = ~((~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp | (~
      mux_474_cse));
  assign nor_1860_nl = ~(nor_151_cse | (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_3 | (~ mux_1126_cse));
  assign not_tmp_580 = MUX_s_1_2_2((nor_1860_nl), (nor_1858_nl), or_5189_cse);
  assign nor_1851_nl = ~(((cfg_out_precision_1_sva_st_154[1]) & cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp)
      | (cfg_out_precision_1_sva_st_154[0]) | (~ mux_tmp_259));
  assign mux_tmp_519 = MUX_s_1_2_2((nor_1851_nl), mux_tmp_259, cvt_11_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp);
  assign and_2214_nl = IntShiftRightSat_49U_6U_17U_lor_12_lpi_1_dfm & mux_tmp_298;
  assign or_828_nl = ((cfg_out_precision_1_sva_st_149[1]) & FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_3)
      | (cfg_out_precision_1_sva_st_149[0]);
  assign mux_524_nl = MUX_s_1_2_2(mux_tmp_298, (and_2214_nl), or_828_nl);
  assign mux_tmp_525 = MUX_s_1_2_2((mux_524_nl), mux_tmp_298, IntShiftRightSat_49U_6U_17U_lor_2_lpi_1_dfm);
  assign mux_538_nl = MUX_s_1_2_2((~ or_tmp_533), mux_tmp_311, IntShiftRightSat_49U_6U_17U_lor_12_lpi_1_dfm);
  assign mux_540_nl = MUX_s_1_2_2(mux_tmp_311, (mux_538_nl), or_461_cse);
  assign mux_tmp_541 = MUX_s_1_2_2((mux_540_nl), mux_tmp_311, IntShiftRightSat_49U_6U_17U_lor_2_lpi_1_dfm);
  assign nor_1838_nl = ~((~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp | (~
      mux_474_cse));
  assign nor_1840_nl = ~(nor_151_cse | (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_3 | (~ mux_1126_cse));
  assign not_tmp_638 = MUX_s_1_2_2((nor_1840_nl), (nor_1838_nl), or_5189_cse);
  assign nor_1828_nl = ~(((cfg_out_precision_1_sva_st_154[1]) & cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp)
      | (cfg_out_precision_1_sva_st_154[0]) | (~ mux_tmp_305));
  assign mux_tmp_560 = MUX_s_1_2_2((nor_1828_nl), mux_tmp_305, cvt_12_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp);
  assign and_2210_nl = IntShiftRightSat_49U_6U_17U_lor_13_lpi_1_dfm & mux_tmp_298;
  assign or_871_nl = (~(((cfg_out_precision_1_sva_st_149[1]) & FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_3)
      | (cfg_out_precision_1_sva_st_149[0]))) | IsNaN_5U_10U_IsNaN_5U_10U_nand_14_itm_2;
  assign mux_tmp_565 = MUX_s_1_2_2((and_2210_nl), mux_tmp_298, or_871_nl);
  assign nor_1827_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ mux_tmp_565));
  assign mux_tmp_566 = MUX_s_1_2_2((nor_1827_nl), mux_tmp_565, cfg_proc_precision_1_sva_st_101[0]);
  assign and_2209_nl = IntShiftRightSat_49U_6U_17U_lor_13_lpi_1_dfm & main_stage_v_2;
  assign mux_576_nl = MUX_s_1_2_2(main_stage_v_2, (and_2209_nl), or_461_cse);
  assign mux_tmp_577 = MUX_s_1_2_2((mux_576_nl), main_stage_v_2, IsNaN_5U_10U_IsNaN_5U_10U_nand_14_itm_2);
  assign nor_1815_nl = ~((cfg_proc_precision_1_sva_st_65[1]) | (~ mux_tmp_577));
  assign mux_tmp_578 = MUX_s_1_2_2((nor_1815_nl), mux_tmp_577, cfg_proc_precision_1_sva_st_65[0]);
  assign nor_1816_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ mux_tmp_578));
  assign mux_tmp_579 = MUX_s_1_2_2((nor_1816_nl), mux_tmp_578, cfg_proc_precision_1_sva_st_101[0]);
  assign nor_1817_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ mux_tmp_579));
  assign mux_tmp_580 = MUX_s_1_2_2((nor_1817_nl), mux_tmp_579, cfg_proc_precision_1_sva_st_101[0]);
  assign or_894_nl = cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp
      | (cfg_out_precision_1_sva_st_154!=2'b10) | (~ and_1386_cse);
  assign or_898_nl = (~ main_stage_v_2) | FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_3
      | (cfg_out_precision_1_sva_st_149[0]) | (~((cfg_out_precision_1_sva_st_149[1])
      & mux_1142_cse));
  assign mux_tmp_585 = MUX_s_1_2_2((or_898_nl), (or_894_nl), or_5189_cse);
  assign and_2208_nl = IntShiftRightSat_49U_6U_17U_lor_14_lpi_1_dfm & or_400_cse_1;
  assign mux_tmp_591 = MUX_s_1_2_2((and_2208_nl), or_400_cse_1, IsNaN_5U_10U_IsNaN_5U_10U_nand_itm_2);
  assign nor_1810_nl = ~((cfg_proc_precision_1_sva_st_89[1]) | (~ mux_tmp_591));
  assign mux_tmp_592 = MUX_s_1_2_2((nor_1810_nl), mux_tmp_591, cfg_proc_precision_1_sva_st_89[0]);
  assign nor_1807_nl = ~((cfg_proc_precision_1_sva_st_64[1]) | (~ mux_1460_cse));
  assign mux_tmp_597 = MUX_s_1_2_2((nor_1807_nl), mux_1460_cse, cfg_proc_precision_1_sva_st_64[0]);
  assign and_2206_cse = IntShiftRightSat_49U_6U_17U_lor_14_lpi_1_dfm & main_stage_v_2;
  assign or_921_nl = (~(((cfg_out_precision_1_sva_st_149[1]) & FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_3)
      | (cfg_out_precision_1_sva_st_149[0]))) | IsNaN_5U_10U_IsNaN_5U_10U_nand_itm_2;
  assign mux_tmp_600 = MUX_s_1_2_2(and_2206_cse, main_stage_v_2, or_921_nl);
  assign nor_1803_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ mux_tmp_600));
  assign mux_tmp_601 = MUX_s_1_2_2((nor_1803_nl), mux_tmp_600, cfg_proc_precision_1_sva_st_101[0]);
  assign nor_1804_nl = ~((cfg_proc_precision_1_sva_st_89[1]) | (~ mux_tmp_601));
  assign mux_tmp_602 = MUX_s_1_2_2((nor_1804_nl), mux_tmp_601, cfg_proc_precision_1_sva_st_89[0]);
  assign mux_611_nl = MUX_s_1_2_2(main_stage_v_2, and_2206_cse, or_461_cse);
  assign mux_tmp_612 = MUX_s_1_2_2((mux_611_nl), main_stage_v_2, IsNaN_5U_10U_IsNaN_5U_10U_nand_itm_2);
  assign nor_1795_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ mux_tmp_612));
  assign mux_tmp_613 = MUX_s_1_2_2((nor_1795_nl), mux_tmp_612, cfg_proc_precision_1_sva_st_101[0]);
  assign nor_1796_nl = ~((cfg_proc_precision_1_sva_st_89[1]) | (~ mux_tmp_613));
  assign mux_tmp_614 = MUX_s_1_2_2((nor_1796_nl), mux_tmp_613, cfg_proc_precision_1_sva_st_89[0]);
  assign nor_1787_nl = ~((~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp | (~
      mux_474_cse));
  assign nor_1789_nl = ~((~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_3 | (~ mux_382_cse));
  assign not_tmp_757 = MUX_s_1_2_2((nor_1789_nl), (nor_1787_nl), or_5189_cse);
  assign nor_1780_nl = ~((cfg_proc_precision_1_sva_st_64[1]) | (~ mux_1489_cse));
  assign mux_tmp_634 = MUX_s_1_2_2((nor_1780_nl), mux_1489_cse, cfg_proc_precision_1_sva_st_64[0]);
  assign and_2202_nl = IntShiftRightSat_49U_6U_17U_lor_15_lpi_1_dfm & main_stage_v_2;
  assign mux_637_nl = MUX_s_1_2_2(main_stage_v_2, (and_2202_nl), or_461_cse);
  assign mux_tmp_638 = MUX_s_1_2_2((mux_637_nl), main_stage_v_2, IsNaN_5U_10U_nor_1_itm_2);
  assign nor_1774_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ mux_tmp_638));
  assign mux_tmp_639 = MUX_s_1_2_2((nor_1774_nl), mux_tmp_638, cfg_proc_precision_1_sva_st_101[0]);
  assign nor_1775_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ mux_tmp_639));
  assign mux_tmp_640 = MUX_s_1_2_2((nor_1775_nl), mux_tmp_639, cfg_proc_precision_1_sva_st_101[0]);
  assign nor_1776_nl = ~((cfg_proc_precision_1_sva_st_89[1]) | (~ mux_tmp_640));
  assign mux_tmp_641 = MUX_s_1_2_2((nor_1776_nl), mux_tmp_640, cfg_proc_precision_1_sva_st_89[0]);
  assign nor_1764_nl = ~((~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp | (~
      mux_474_cse));
  assign nor_1766_nl = ~((~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2 | (~ mux_417_cse));
  assign not_tmp_811 = MUX_s_1_2_2((nor_1766_nl), (nor_1764_nl), or_5189_cse);
  assign nor_1762_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ main_stage_v_2));
  assign mux_tmp_658 = MUX_s_1_2_2((nor_1762_nl), main_stage_v_2, cfg_proc_precision_1_sva_st_101[0]);
  assign and_2199_cse = IntShiftRightSat_49U_6U_17U_lor_16_lpi_1_dfm & main_stage_v_2;
  assign or_1015_nl = (~(((cfg_out_precision_1_sva_st_149[1]) & FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_3)
      | (cfg_out_precision_1_sva_st_149[0]))) | IsNaN_5U_10U_nor_14_itm_2;
  assign mux_tmp_678 = MUX_s_1_2_2(and_2199_cse, main_stage_v_2, or_1015_nl);
  assign nor_1748_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ mux_tmp_678));
  assign mux_tmp_679 = MUX_s_1_2_2((nor_1748_nl), mux_tmp_678, cfg_proc_precision_1_sva_st_101[0]);
  assign nor_1749_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ mux_tmp_679));
  assign mux_tmp_680 = MUX_s_1_2_2((nor_1749_nl), mux_tmp_679, cfg_proc_precision_1_sva_st_101[0]);
  assign nor_1750_nl = ~((cfg_proc_precision_1_sva_st_89[1]) | (~ mux_tmp_680));
  assign mux_tmp_681 = MUX_s_1_2_2((nor_1750_nl), mux_tmp_680, cfg_proc_precision_1_sva_st_89[0]);
  assign mux_691_nl = MUX_s_1_2_2(main_stage_v_2, and_2199_cse, or_461_cse);
  assign mux_tmp_692 = MUX_s_1_2_2((mux_691_nl), main_stage_v_2, IsNaN_5U_10U_nor_14_itm_2);
  assign nor_1738_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ mux_tmp_692));
  assign mux_tmp_693 = MUX_s_1_2_2((nor_1738_nl), mux_tmp_692, cfg_proc_precision_1_sva_st_101[0]);
  assign nor_1739_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ mux_tmp_693));
  assign mux_tmp_694 = MUX_s_1_2_2((nor_1739_nl), mux_tmp_693, cfg_proc_precision_1_sva_st_101[0]);
  assign nor_1740_nl = ~((cfg_proc_precision_1_sva_st_89[1]) | (~ mux_tmp_694));
  assign mux_tmp_695 = MUX_s_1_2_2((nor_1740_nl), mux_tmp_694, cfg_proc_precision_1_sva_st_89[0]);
  assign nor_1728_nl = ~((~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp | (~
      mux_474_cse));
  assign nor_1730_nl = ~((~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_3 | (~ mux_417_cse));
  assign not_tmp_899 = MUX_s_1_2_2((nor_1730_nl), (nor_1728_nl), or_5189_cse);
  assign nor_1718_nl = ~((reg_cfg_proc_precision_1_sva_st_40_cse[1]) | (~ mux_1489_cse));
  assign mux_tmp_719 = MUX_s_1_2_2((nor_1718_nl), mux_1489_cse, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign nor_1719_nl = ~((cfg_proc_precision_1_sva_st_64[1]) | (~ mux_tmp_719));
  assign mux_tmp_720 = MUX_s_1_2_2((nor_1719_nl), mux_tmp_719, cfg_proc_precision_1_sva_st_64[0]);
  assign and_2194_cse = IntShiftRightSat_49U_6U_17U_lor_lpi_1_dfm & main_stage_v_2;
  assign or_1072_nl = (~(((cfg_out_precision_1_sva_st_149[1]) & FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_3)
      | (cfg_out_precision_1_sva_st_149[0]))) | IsNaN_5U_10U_nor_itm_2;
  assign mux_tmp_723 = MUX_s_1_2_2(and_2194_cse, main_stage_v_2, or_1072_nl);
  assign nor_1711_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ mux_tmp_723));
  assign mux_tmp_724 = MUX_s_1_2_2((nor_1711_nl), mux_tmp_723, cfg_proc_precision_1_sva_st_101[0]);
  assign nor_1712_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ mux_tmp_724));
  assign mux_tmp_725 = MUX_s_1_2_2((nor_1712_nl), mux_tmp_724, cfg_proc_precision_1_sva_st_101[0]);
  assign nor_1713_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ mux_tmp_725));
  assign mux_tmp_726 = MUX_s_1_2_2((nor_1713_nl), mux_tmp_725, cfg_proc_precision_1_sva_st_101[0]);
  assign nor_1714_nl = ~((cfg_proc_precision_1_sva_st_89[1]) | (~ mux_tmp_726));
  assign mux_tmp_727 = MUX_s_1_2_2((nor_1714_nl), mux_tmp_726, cfg_proc_precision_1_sva_st_89[0]);
  assign mux_738_nl = MUX_s_1_2_2(main_stage_v_2, and_2194_cse, or_461_cse);
  assign mux_tmp_739 = MUX_s_1_2_2((mux_738_nl), main_stage_v_2, IsNaN_5U_10U_nor_itm_2);
  assign nor_1699_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ mux_tmp_739));
  assign mux_tmp_740 = MUX_s_1_2_2((nor_1699_nl), mux_tmp_739, cfg_proc_precision_1_sva_st_101[0]);
  assign nor_1700_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ mux_tmp_740));
  assign mux_tmp_741 = MUX_s_1_2_2((nor_1700_nl), mux_tmp_740, cfg_proc_precision_1_sva_st_101[0]);
  assign nor_1701_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ mux_tmp_741));
  assign mux_tmp_742 = MUX_s_1_2_2((nor_1701_nl), mux_tmp_741, cfg_proc_precision_1_sva_st_101[0]);
  assign nor_1702_nl = ~((cfg_proc_precision_1_sva_st_89[1]) | (~ mux_tmp_742));
  assign mux_tmp_743 = MUX_s_1_2_2((nor_1702_nl), mux_tmp_742, cfg_proc_precision_1_sva_st_89[0]);
  assign nor_1687_nl = ~((~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_tmp | (~
      mux_344_cse));
  assign nor_1689_nl = ~((~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_3 | (~ mux_417_cse));
  assign not_tmp_989 = MUX_s_1_2_2((nor_1689_nl), (nor_1687_nl), or_5189_cse);
  assign nor_1685_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ mux_tmp_658));
  assign mux_tmp_765 = MUX_s_1_2_2((nor_1685_nl), mux_tmp_658, cfg_proc_precision_1_sva_st_101[0]);
  assign nor_1686_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ mux_tmp_765));
  assign mux_tmp_766 = MUX_s_1_2_2((nor_1686_nl), mux_tmp_765, cfg_proc_precision_1_sva_st_101[0]);
  assign or_tmp_1375 = nor_1672_cse | (~ main_stage_v_3) | cfg_mode_eql_1_sva_6;
  assign or_tmp_1393 = ~(cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2
      & (cfg_out_precision_1_sva_st_113==2'b10) & mux_tmp_416);
  assign mux_tmp_944 = MUX_s_1_2_2(and_2186_cse, and_tmp_12, main_stage_v_1);
  assign mux_tmp_945 = MUX_s_1_2_2(mux_tmp_944, and_tmp_50, main_stage_v_2);
  assign and_tmp_165 = or_3538_cse & or_1159_cse;
  assign mux_tmp_946 = MUX_s_1_2_2(and_1386_cse, and_tmp_50, main_stage_v_2);
  assign mux_tmp_947 = MUX_s_1_2_2(mux_tmp_946, and_tmp_165, main_stage_v_3);
  assign and_tmp_166 = or_3542_cse & or_1159_cse;
  assign mux_tmp_960 = MUX_s_1_2_2(and_2186_cse, mux_tmp_123, main_stage_v_1);
  assign mux_tmp_961 = MUX_s_1_2_2(mux_tmp_960, and_tmp_79, main_stage_v_2);
  assign and_tmp_168 = or_3542_cse & and_tmp_165;
  assign mux_tmp_962 = MUX_s_1_2_2(and_tmp_19, and_tmp_79, main_stage_v_2);
  assign mux_tmp_963 = MUX_s_1_2_2(mux_tmp_962, and_tmp_168, main_stage_v_3);
  assign nor_1545_nl = ~((cfg_proc_precision_1_sva_st_102[1]) | (~ or_1159_cse));
  assign mux_969_nl = MUX_s_1_2_2((nor_1545_nl), or_1159_cse, cfg_proc_precision_1_sva_st_102[0]);
  assign and_tmp_169 = or_3538_cse & (mux_969_nl);
  assign nor_1534_nl = ~((cfg_proc_precision_1_sva_st_90[1]) | (~ or_1159_cse));
  assign mux_tmp_986 = MUX_s_1_2_2((nor_1534_nl), or_1159_cse, cfg_proc_precision_1_sva_st_90[0]);
  assign nor_1535_nl = ~((cfg_proc_precision_1_sva_st_102[1]) | (~ mux_tmp_986));
  assign mux_tmp_987 = MUX_s_1_2_2((nor_1535_nl), mux_tmp_986, cfg_proc_precision_1_sva_st_102[0]);
  assign mux_tmp_992 = MUX_s_1_2_2(mux_tmp_944, mux_1142_cse, main_stage_v_2);
  assign mux_tmp_994 = MUX_s_1_2_2(mux_989_cse, mux_tmp_987, main_stage_v_3);
  assign and_2247_nl = (~((cfg_out_precision_1_sva_6[1]) & (cfg_out_precision_1_sva_st_144[1])))
      & and_tmp_165;
  assign mux_1013_nl = MUX_s_1_2_2((and_2247_nl), and_tmp_165, or_1919_cse);
  assign mux_1014_nl = MUX_s_1_2_2(mux_tmp_946, (mux_1013_nl), main_stage_v_3);
  assign nor_208_nl = ~((cfg_out_precision_1_sva_st_144[0]) | (~ cvt_unequal_tmp_21));
  assign mux_tmp_1015 = MUX_s_1_2_2(mux_tmp_947, (mux_1014_nl), nor_208_nl);
  assign nor_1486_cse = ~((cfg_out_precision_1_sva_st_156[1]) | (~ mux_tmp_987));
  assign or_1644_nl = (~ cvt_unequal_tmp_21) | cfg_mode_eql_1_sva_6 | (cfg_out_precision_1_sva_6!=2'b10)
      | (cfg_out_precision_1_sva_st_156[0]);
  assign mux_tmp_1038 = MUX_s_1_2_2(nor_1486_cse, mux_tmp_987, or_1644_nl);
  assign nand_tmp_30 = (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt
      | (~ main_stage_v_3) | mux_tmp_1038;
  assign nor_1487_nl = ~((~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt
      | (main_stage_v_3 & (~ mux_tmp_1038)));
  assign or_1643_nl = (cfg_out_precision_1_sva_st_149!=2'b10) | (~ cvt_unequal_tmp_20)
      | cfg_mode_eql_1_sva_5 | (cfg_out_precision_1_sva_st_113!=2'b10);
  assign mux_tmp_1039 = MUX_s_1_2_2((nor_1487_nl), nand_tmp_30, or_1643_nl);
  assign and_tmp_171 = main_stage_v_3 & mux_tmp_1038;
  assign or_tmp_1650 = (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt
      | (~ and_tmp_171);
  assign mux_1040_nl = MUX_s_1_2_2(mux_tmp_1039, (~ or_tmp_1650), cfg_proc_precision_1_sva_st_65[1]);
  assign mux_tmp_1041 = MUX_s_1_2_2((mux_1040_nl), mux_tmp_1039, cfg_proc_precision_1_sva_st_65[0]);
  assign mux_1042_nl = MUX_s_1_2_2(mux_tmp_1041, (~ or_tmp_1650), cfg_proc_precision_1_sva_st_89[1]);
  assign mux_tmp_1043 = MUX_s_1_2_2((mux_1042_nl), mux_tmp_1041, cfg_proc_precision_1_sva_st_89[0]);
  assign mux_1046_nl = MUX_s_1_2_2(nand_tmp_30, (~ or_tmp_1650), reg_cfg_proc_precision_1_sva_st_40_cse[1]);
  assign mux_tmp_1047 = MUX_s_1_2_2((mux_1046_nl), nand_tmp_30, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign mux_1048_nl = MUX_s_1_2_2(mux_tmp_1047, (~ or_tmp_1650), reg_cfg_proc_precision_1_sva_st_40_cse[1]);
  assign mux_tmp_1049 = MUX_s_1_2_2((mux_1048_nl), mux_tmp_1047, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign nor_1464_nl = ~((cfg_out_precision_1_sva_6[1]) | (~ and_tmp_168));
  assign mux_1072_nl = MUX_s_1_2_2((nor_1464_nl), and_tmp_168, or_1919_cse);
  assign mux_1073_nl = MUX_s_1_2_2(mux_tmp_962, (mux_1072_nl), main_stage_v_3);
  assign nor_250_nl = ~((~ cvt_unequal_tmp_21) | (cfg_out_precision_1_sva_st_156!=2'b10));
  assign mux_tmp_1074 = MUX_s_1_2_2(mux_tmp_963, (mux_1073_nl), nor_250_nl);
  assign nor_1455_nl = ~((cfg_out_precision_1_sva_st_156[1]) | (~ and_tmp_169));
  assign or_1745_nl = cfg_mode_eql_1_sva_6 | (cfg_out_precision_1_sva_6!=2'b10) |
      (cfg_out_precision_1_sva_st_156[0]);
  assign mux_1086_nl = MUX_s_1_2_2((nor_1455_nl), and_tmp_169, or_1745_nl);
  assign mux_1087_nl = MUX_s_1_2_2(mux_tmp_962, (mux_1086_nl), main_stage_v_3);
  assign mux_976_nl = MUX_s_1_2_2(mux_tmp_962, and_tmp_169, main_stage_v_3);
  assign mux_tmp_1088 = MUX_s_1_2_2((mux_976_nl), (mux_1087_nl), cvt_unequal_tmp_21);
  assign or_1774_nl = nor_1589_cse | (~ cvt_unequal_tmp_21) | cfg_mode_eql_1_sva_6
      | (cfg_out_precision_1_sva_6!=2'b10) | (cfg_out_precision_1_sva_st_156[0]);
  assign mux_tmp_1100 = MUX_s_1_2_2(nor_1486_cse, mux_tmp_987, or_1774_nl);
  assign nand_tmp_36 = (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt
      | (~ main_stage_v_3) | mux_tmp_1100;
  assign nor_1446_nl = ~((~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt
      | (main_stage_v_3 & (~ mux_tmp_1100)));
  assign or_1773_nl = nor_151_cse | (cfg_out_precision_1_sva_st_149!=2'b10) | (~
      cvt_unequal_tmp_20) | cfg_mode_eql_1_sva_5 | (cfg_out_precision_1_sva_st_113!=2'b10);
  assign mux_tmp_1101 = MUX_s_1_2_2((nor_1446_nl), nand_tmp_36, or_1773_nl);
  assign and_tmp_175 = main_stage_v_3 & mux_tmp_1100;
  assign or_tmp_1780 = (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt
      | (~ and_tmp_175);
  assign mux_1102_nl = MUX_s_1_2_2(mux_tmp_1101, (~ or_tmp_1780), cfg_proc_precision_1_sva_st_65[1]);
  assign mux_tmp_1103 = MUX_s_1_2_2((mux_1102_nl), mux_tmp_1101, cfg_proc_precision_1_sva_st_65[0]);
  assign mux_1104_nl = MUX_s_1_2_2(mux_tmp_1103, (~ or_tmp_1780), cfg_proc_precision_1_sva_st_89[1]);
  assign mux_tmp_1105 = MUX_s_1_2_2((mux_1104_nl), mux_tmp_1103, cfg_proc_precision_1_sva_st_89[0]);
  assign mux_1108_nl = MUX_s_1_2_2(nand_tmp_36, (~ or_tmp_1780), reg_cfg_proc_precision_1_sva_st_40_cse[1]);
  assign mux_tmp_1109 = MUX_s_1_2_2((mux_1108_nl), nand_tmp_36, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign mux_1110_nl = MUX_s_1_2_2(mux_tmp_1109, (~ or_tmp_1780), reg_cfg_proc_precision_1_sva_st_40_cse[1]);
  assign mux_tmp_1111 = MUX_s_1_2_2((mux_1110_nl), mux_tmp_1109, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign mux_1151_nl = MUX_s_1_2_2(mux_tmp_1041, (~ or_tmp_1650), cfg_proc_precision_1_sva_st_101[1]);
  assign mux_tmp_1152 = MUX_s_1_2_2((mux_1151_nl), mux_tmp_1041, cfg_proc_precision_1_sva_st_101[0]);
  assign nor_1387_nl = ~((cfg_proc_precision_1_sva_st_102[1]) | (~ or_3538_cse));
  assign mux_tmp_1196 = MUX_s_1_2_2((nor_1387_nl), or_3538_cse, cfg_proc_precision_1_sva_st_102[0]);
  assign nor_1388_nl = ~((cfg_proc_precision_1_sva_st_66[1]) | (~ mux_tmp_1196));
  assign mux_tmp_1197 = MUX_s_1_2_2((nor_1388_nl), mux_tmp_1196, cfg_proc_precision_1_sva_st_66[0]);
  assign nand_202_cse = ~(main_stage_v_3 & mux_tmp_1197);
  assign or_tmp_1981 = (cfg_out_precision_1_sva_6!=2'b00) | nand_202_cse;
  assign or_tmp_1992 = (cfg_out_precision_1_sva_6!=2'b01) | nand_202_cse;
  assign nor_1371_nl = ~((cfg_proc_precision_1_sva_st_66[1]) | (~ main_stage_v_3));
  assign mux_tmp_1225 = MUX_s_1_2_2((nor_1371_nl), main_stage_v_3, cfg_proc_precision_1_sva_st_66[0]);
  assign nor_1372_nl = ~((cfg_proc_precision_1_sva_st_90[1]) | (~ mux_tmp_1225));
  assign mux_tmp_1226 = MUX_s_1_2_2((nor_1372_nl), mux_tmp_1225, cfg_proc_precision_1_sva_st_90[0]);
  assign nor_1373_nl = ~((cfg_proc_precision_1_sva_st_102[1]) | (~ mux_tmp_1226));
  assign mux_tmp_1227 = MUX_s_1_2_2((nor_1373_nl), mux_tmp_1226, cfg_proc_precision_1_sva_st_102[0]);
  assign mux_tmp_1264 = MUX_s_1_2_2(and_283_cse, and_tmp_94, or_5189_cse);
  assign or_tmp_2136 = (~ cvt_unequal_tmp_19) | cfg_mode_eql_1_sva_4 | (cfg_out_precision_1_sva_st_154!=2'b10)
      | (~ main_stage_v_1);
  assign or_tmp_2139 = main_stage_v_2 | (~ or_tmp_2136);
  assign mux_1269_nl = MUX_s_1_2_2(or_tmp_2139, (~ or_tmp_2136), cfg_proc_precision_1_sva_st_101[1]);
  assign mux_tmp_1270 = MUX_s_1_2_2((mux_1269_nl), or_tmp_2139, cfg_proc_precision_1_sva_st_101[0]);
  assign or_2140_cse = nor_50_cse | (cfg_out_precision_1_sva_st_149[0]);
  assign mux_1271_nl = MUX_s_1_2_2(mux_tmp_1270, (~ or_tmp_2136), cfg_proc_precision_1_sva_st_89[1]);
  assign mux_1272_nl = MUX_s_1_2_2((mux_1271_nl), mux_tmp_1270, cfg_proc_precision_1_sva_st_89[0]);
  assign mux_1273_nl = MUX_s_1_2_2(or_tmp_2136, (~ (mux_1272_nl)), cfg_out_precision_1_sva_st_149[1]);
  assign mux_1274_nl = MUX_s_1_2_2((mux_1273_nl), or_tmp_2136, or_2140_cse);
  assign mux_1275_nl = MUX_s_1_2_2((~ or_tmp_2139), (mux_1274_nl), or_1587_cse);
  assign mux_tmp_1276 = MUX_s_1_2_2((mux_1275_nl), or_tmp_2136, or_5189_cse);
  assign mux_tmp_1280 = MUX_s_1_2_2(mux_1464_cse, main_stage_v_1, or_5189_cse);
  assign mux_1281_nl = MUX_s_1_2_2(mux_tmp_1280, (~ mux_tmp_1276), reg_cfg_proc_precision_1_sva_st_40_cse[1]);
  assign mux_tmp_1282 = MUX_s_1_2_2((mux_1281_nl), mux_tmp_1280, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign mux_1325_nl = MUX_s_1_2_2(mux_tmp_1270, (~ or_tmp_2136), cfg_proc_precision_1_sva_st_101[1]);
  assign mux_tmp_1326 = MUX_s_1_2_2((mux_1325_nl), mux_tmp_1270, cfg_proc_precision_1_sva_st_101[0]);
  assign mux_1327_nl = MUX_s_1_2_2(mux_tmp_1326, (~ or_tmp_2136), cfg_proc_precision_1_sva_st_89[1]);
  assign mux_1328_nl = MUX_s_1_2_2((mux_1327_nl), mux_tmp_1326, cfg_proc_precision_1_sva_st_89[0]);
  assign mux_1329_nl = MUX_s_1_2_2(or_tmp_2136, (~ (mux_1328_nl)), cfg_out_precision_1_sva_st_149[1]);
  assign mux_1330_nl = MUX_s_1_2_2((mux_1329_nl), or_tmp_2136, or_2140_cse);
  assign mux_1331_nl = MUX_s_1_2_2((~ or_tmp_2139), (mux_1330_nl), or_1587_cse);
  assign mux_tmp_1332 = MUX_s_1_2_2((mux_1331_nl), or_tmp_2136, or_5189_cse);
  assign mux_tmp_1337 = MUX_s_1_2_2(mux_1494_cse, main_stage_v_1, or_5189_cse);
  assign mux_1338_nl = MUX_s_1_2_2(mux_tmp_1337, (~ mux_tmp_1332), reg_cfg_proc_precision_1_sva_st_40_cse[1]);
  assign mux_tmp_1339 = MUX_s_1_2_2((mux_1338_nl), mux_tmp_1337, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign mux_1340_nl = MUX_s_1_2_2(mux_tmp_1339, (~ mux_tmp_1332), reg_cfg_proc_precision_1_sva_st_40_cse[1]);
  assign mux_tmp_1341 = MUX_s_1_2_2((mux_1340_nl), mux_tmp_1339, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign nor_1320_cse = ~(main_stage_v_2 | (~ or_tmp_2136));
  assign and_2246_cse = nand_190_cse & or_tmp_2136;
  assign or_2232_nl = nor_151_cse | (cfg_out_precision_1_sva_st_149[0]);
  assign mux_1405_nl = MUX_s_1_2_2(and_2246_cse, or_tmp_2136, or_2232_nl);
  assign mux_1406_nl = MUX_s_1_2_2((mux_1405_nl), or_tmp_2136, nor_2219_cse);
  assign mux_1407_nl = MUX_s_1_2_2((mux_1406_nl), or_tmp_2136, nor_50_cse);
  assign mux_1408_nl = MUX_s_1_2_2(nor_1320_cse, (mux_1407_nl), or_1587_cse);
  assign mux_tmp_1409 = MUX_s_1_2_2((mux_1408_nl), or_tmp_2136, or_5189_cse);
  assign or_2245_nl = (~((cfg_out_precision_1_sva_st_149!=2'b10) | (~ main_stage_v_2)))
      | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt;
  assign mux_1416_nl = MUX_s_1_2_2((or_2245_nl), or_5189_cse, nor_151_cse);
  assign mux_1417_nl = MUX_s_1_2_2((mux_1416_nl), or_5189_cse, nor_2219_cse);
  assign mux_1418_nl = MUX_s_1_2_2((mux_1417_nl), or_5189_cse, nor_50_cse);
  assign or_2246_nl = main_stage_v_2 | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt;
  assign mux_tmp_1419 = MUX_s_1_2_2((or_2246_nl), (mux_1418_nl), or_1198_cse);
  assign not_tmp_1709 = ~(nor_8_cse | nor_2150_cse | (cfg_out_precision_1_sva_st_154!=2'b10)
      | mux_tmp_1419);
  assign nand_tmp_48 = ~(main_stage_v_1 & not_tmp_1709);
  assign mux_1430_nl = MUX_s_1_2_2(and_2246_cse, or_tmp_2136, cfg_out_precision_1_sva_st_149[0]);
  assign mux_1431_nl = MUX_s_1_2_2((mux_1430_nl), or_tmp_2136, nor_151_cse);
  assign mux_1432_nl = MUX_s_1_2_2((mux_1431_nl), or_tmp_2136, nor_2219_cse);
  assign mux_1433_nl = MUX_s_1_2_2((mux_1432_nl), or_tmp_2136, nor_50_cse);
  assign mux_1434_nl = MUX_s_1_2_2(nor_1320_cse, (mux_1433_nl), or_1587_cse);
  assign mux_tmp_1435 = MUX_s_1_2_2((mux_1434_nl), or_tmp_2136, or_5189_cse);
  assign and_306_nl = FpIntToFloat_17U_5U_10U_else_unequal_tmp_4 & (~(cvt_5_FpMantRNE_17U_11U_else_and_1_svs
      | (~ main_stage_v_2)));
  assign or_2306_nl = (~ cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2)
      | cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  assign mux_tmp_1469 = MUX_s_1_2_2((and_306_nl), main_stage_v_2, or_2306_nl);
  assign or_tmp_2432 = (~ chn_in_rsci_bawt) | cfg_mode_eql_rsci_d;
  assign or_tmp_2466 = IsNaN_8U_23U_IsNaN_8U_23U_nand_4_tmp | IsNaN_8U_23U_nor_4_tmp;
  assign or_tmp_2469 = IsNaN_8U_23U_nor_4_itm_2 | IsNaN_8U_23U_IsNaN_8U_23U_nand_4_itm_2;
  assign mux_tmp_1566 = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, cvt_16_FpMantRNE_24U_11U_else_and_4_svs_2);
  assign or_tmp_2569 = (~ cvt_16_FpMantRNE_24U_11U_else_and_4_svs_2) | (~ reg_chn_out_rsci_ld_core_psct_cse)
      | chn_out_rsci_bawt | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_tmp_1570 = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, cvt_15_FpMantRNE_24U_11U_else_and_3_svs_2);
  assign or_tmp_2571 = (~ cvt_15_FpMantRNE_24U_11U_else_and_3_svs_2) | (~ reg_chn_out_rsci_ld_core_psct_cse)
      | chn_out_rsci_bawt | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_tmp_1574 = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, cvt_14_FpMantRNE_24U_11U_else_and_3_svs_2);
  assign or_tmp_2573 = (~ cvt_14_FpMantRNE_24U_11U_else_and_3_svs_2) | (~ reg_chn_out_rsci_ld_core_psct_cse)
      | chn_out_rsci_bawt | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_tmp_1578 = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, cvt_13_FpMantRNE_24U_11U_else_and_2_svs_2);
  assign or_tmp_2575 = (~ cvt_13_FpMantRNE_24U_11U_else_and_2_svs_2) | (~ reg_chn_out_rsci_ld_core_psct_cse)
      | chn_out_rsci_bawt | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_tmp_1582 = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, cvt_12_FpMantRNE_24U_11U_else_and_3_svs_2);
  assign or_tmp_2577 = (~ cvt_12_FpMantRNE_24U_11U_else_and_3_svs_2) | (~ reg_chn_out_rsci_ld_core_psct_cse)
      | chn_out_rsci_bawt | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_tmp_1586 = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, cvt_11_FpMantRNE_24U_11U_else_and_2_svs_2);
  assign or_tmp_2579 = (~ cvt_11_FpMantRNE_24U_11U_else_and_2_svs_2) | (~ reg_chn_out_rsci_ld_core_psct_cse)
      | chn_out_rsci_bawt | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_tmp_1592 = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, cvt_9_FpMantRNE_24U_11U_else_and_1_svs_2);
  assign or_tmp_2588 = (~ cvt_9_FpMantRNE_24U_11U_else_and_1_svs_2) | (~ reg_chn_out_rsci_ld_core_psct_cse)
      | chn_out_rsci_bawt | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_tmp_1596 = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, cvt_8_FpMantRNE_24U_11U_else_and_3_svs_2);
  assign or_tmp_2590 = (~ cvt_8_FpMantRNE_24U_11U_else_and_3_svs_2) | (~ reg_chn_out_rsci_ld_core_psct_cse)
      | chn_out_rsci_bawt | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign nand_230_nl = ~(cvt_7_FpMantRNE_24U_11U_else_and_2_svs_2 & main_stage_v_1
      & (cfg_proc_precision_1_sva_st_64==2'b10));
  assign mux_tmp_1600 = MUX_s_1_2_2((nand_230_nl), or_tmp_19, or_5189_cse);
  assign or_tmp_2595 = (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt
      | (~ cvt_7_FpMantRNE_24U_11U_else_and_2_svs_2) | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_tmp_1606 = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, cvt_5_FpMantRNE_24U_11U_else_and_1_svs_2);
  assign or_tmp_2604 = (~ cvt_5_FpMantRNE_24U_11U_else_and_1_svs_2) | (~ reg_chn_out_rsci_ld_core_psct_cse)
      | chn_out_rsci_bawt | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_tmp_1610 = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, cvt_4_FpMantRNE_24U_11U_else_and_2_svs_2);
  assign or_tmp_2606 = (~ cvt_4_FpMantRNE_24U_11U_else_and_2_svs_2) | (~ reg_chn_out_rsci_ld_core_psct_cse)
      | chn_out_rsci_bawt | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_tmp_1614 = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, cvt_3_FpMantRNE_24U_11U_else_and_1_svs_2);
  assign or_tmp_2608 = (~ cvt_3_FpMantRNE_24U_11U_else_and_1_svs_2) | (~ reg_chn_out_rsci_ld_core_psct_cse)
      | chn_out_rsci_bawt | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_tmp_1618 = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, cvt_2_FpMantRNE_24U_11U_else_and_1_svs_2);
  assign or_tmp_2610 = (~ cvt_2_FpMantRNE_24U_11U_else_and_1_svs_2) | (~ reg_chn_out_rsci_ld_core_psct_cse)
      | chn_out_rsci_bawt | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_tmp_1622 = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, cvt_1_FpMantRNE_24U_11U_else_and_svs_2);
  assign or_tmp_2612 = (~ cvt_1_FpMantRNE_24U_11U_else_and_svs_2) | (~ reg_chn_out_rsci_ld_core_psct_cse)
      | chn_out_rsci_bawt | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign and_dcpl_93 = (~ chn_out_rsci_bawt) & reg_chn_out_rsci_ld_core_psct_cse;
  assign or_dcpl_4 = and_dcpl_93 | (~ main_stage_v_3);
  assign and_dcpl_98 = main_stage_v_3 & (~ cvt_unequal_tmp_21) & or_5189_cse;
  assign and_dcpl_102 = (~ cfg_mode_eql_1_sva_6) & main_stage_v_3 & or_5189_cse;
  assign and_dcpl_103 = or_5189_cse & main_stage_v_3;
  assign and_dcpl_105 = (~ main_stage_v_3) & chn_out_rsci_bawt & reg_chn_out_rsci_ld_core_psct_cse;
  assign and_dcpl_114 = or_5189_cse & main_stage_v_1;
  assign or_dcpl_15 = and_dcpl_3 | ((reg_cfg_proc_precision_1_sva_st_40_cse==2'b10));
  assign or_dcpl_16 = or_dcpl_15 | (~ main_stage_v_1);
  assign or_dcpl_30 = ~((~((reg_cfg_proc_precision_1_sva_st_40_cse==2'b10))) & main_stage_v_1);
  assign or_dcpl_32 = or_dcpl_15 | or_dcpl_30;
  assign and_dcpl_204 = or_4550_cse & or_5189_cse;
  assign and_dcpl_209 = (cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_nor_4_cse | cvt_1_IntShiftRight_49U_6U_17U_obits_fixed_nor_tmp)
      & or_5189_cse;
  assign and_dcpl_217 = (cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse | cvt_2_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp)
      & or_5189_cse;
  assign and_dcpl_224 = (cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse | cvt_3_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp)
      & or_5189_cse;
  assign or_dcpl_108 = (cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[16])
      | cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  assign and_dcpl_228 = (cfg_out_precision_1_sva_st_154==2'b10);
  assign or_dcpl_109 = cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse | cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  assign nor_tmp_636 = ~((~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt
      | (~ main_stage_v_2));
  assign or_dcpl_110 = (cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_acc_1_tmp[16])
      | cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_and_3_tmp;
  assign or_dcpl_111 = cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse | cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp;
  assign not_tmp_2254 = ~((cfg_out_precision_1_sva_st_154[1]) & and_tmp_12);
  assign or_tmp_2960 = (cfg_out_precision_1_sva_st_154[0]) | not_tmp_2254;
  assign or_dcpl_113 = cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp | (cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[16]);
  assign or_dcpl_114 = cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse | cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  assign and_tmp_225 = or_400_cse_1 & mux_tmp_455;
  assign or_dcpl_115 = (cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[16])
      | cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  assign or_dcpl_116 = cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse | cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  assign or_dcpl_119 = cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp | (cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[16]);
  assign or_dcpl_120 = cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse | cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp;
  assign and_dcpl_301 = (cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_nor_9_cse | cvt_9_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp)
      & or_5189_cse;
  assign or_dcpl_124 = cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp | (cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[16]);
  assign or_dcpl_125 = cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse | cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  assign or_dcpl_126 = (cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[16])
      | cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  assign or_dcpl_127 = cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse | cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  assign or_dcpl_130 = cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp | (cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[16]);
  assign or_dcpl_131 = cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse | cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp;
  assign or_dcpl_132 = (cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_acc_2_tmp[16])
      | cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_and_5_tmp;
  assign or_dcpl_133 = cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_nor_14_cse | cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp;
  assign or_tmp_3025 = nor_2219_cse | nor_50_cse | (cfg_out_precision_1_sva_st_149[0]);
  assign or_tmp_3032 = (cfg_out_precision_1_sva_st_154[0]) | not_tmp_270;
  assign or_dcpl_136 = cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp | (cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[16]);
  assign and_dcpl_363 = main_stage_v_1 & (cfg_out_precision_1_sva_st_154==2'b10);
  assign or_dcpl_137 = cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse | cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp;
  assign or_dcpl_139 = cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_and_7_tmp | (cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_acc_3_tmp[16]);
  assign or_dcpl_140 = cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_nor_19_cse | cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp;
  assign or_dcpl_143 = cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_and_9_tmp | (cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_acc_4_tmp[16]);
  assign or_dcpl_144 = cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_nor_24_cse | cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_nor_20_tmp;
  assign nor_1063_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ and_tmp_225));
  assign mux_tmp_1813 = MUX_s_1_2_2((nor_1063_nl), and_tmp_225, cfg_proc_precision_1_sva_st_101[0]);
  assign and_dcpl_401 = or_5189_cse & main_stage_v_2;
  assign and_dcpl_407 = (~ or_4862_cse) & (cfg_out_precision_1_sva_st_113[0]) & or_5189_cse
      & (~ (cfg_out_precision_1_sva_st_113[1]));
  assign and_dcpl_408 = or_5189_cse & (~ cvt_unequal_tmp_20);
  assign or_dcpl_147 = or_4862_cse | (cfg_out_precision_1_sva_st_113!=2'b01);
  assign and_dcpl_409 = or_dcpl_147 & and_dcpl_408;
  assign and_dcpl_411 = or_4862_cse & cvt_unequal_tmp_20 & or_5189_cse;
  assign and_dcpl_417 = (~ (cfg_proc_precision_1_sva_st_65[0])) & (~ cvt_unequal_tmp_20)
      & or_5189_cse;
  assign and_dcpl_420 = or_5189_cse & cvt_unequal_tmp_20;
  assign and_dcpl_424 = or_4862_cse & or_5189_cse;
  assign and_dcpl_425 = ((~ or_4862_cse) | (cfg_out_precision_1_sva_st_113[0])) &
      and_dcpl_420;
  assign and_dcpl_433 = (~ or_4862_cse) & (cfg_out_precision_1_sva_st_113==2'b01)
      & and_dcpl_408;
  assign or_dcpl_151 = ~(or_4862_cse & (~((cfg_proc_precision_1_sva_st_89==2'b10))));
  assign and_dcpl_444 = ~((cfg_out_precision_1_sva_st_113!=2'b00));
  assign and_dcpl_446 = or_4862_cse & and_dcpl_444 & and_dcpl_420;
  assign mux_1839_nl = MUX_s_1_2_2(nor_57_cse, nor_2099_cse, nor_50_cse);
  assign nor_1053_nl = ~(nor_1672_cse | (cfg_out_precision_1_sva_6!=2'b10));
  assign mux_1841_nl = MUX_s_1_2_2(or_1157_cse, (nor_1053_nl), cvt_unequal_tmp_21);
  assign not_tmp_2422 = MUX_s_1_2_2((mux_1841_nl), (mux_1839_nl), or_5189_cse);
  assign and_dcpl_458 = and_dcpl_444 & cvt_unequal_tmp_20;
  assign and_tmp_248 = or_5254_cse & mux_tmp_987;
  assign or_dcpl_160 = and_1021_cse | (cfg_out_precision_1_sva_st_113[0]);
  assign and_dcpl_473 = and_tmp_225 & or_5189_cse;
  assign and_dcpl_479 = (cfg_proc_precision_1_sva_st_89==2'b10);
  assign or_dcpl_163 = (~ or_4862_cse) | and_dcpl_479;
  assign and_dcpl_481 = and_dcpl_458 & or_5189_cse;
  assign nor_1025_nl = ~((cfg_proc_precision_1_sva_st_102[1]) | (~ and_tmp_165));
  assign mux_tmp_1899 = MUX_s_1_2_2((nor_1025_nl), and_tmp_165, cfg_proc_precision_1_sva_st_102[0]);
  assign and_dcpl_499 = mux_tmp_455 & or_5189_cse;
  assign or_dcpl_178 = ~(or_1159_cse & (~((cfg_proc_precision_1_sva_st_90==2'b10))));
  assign and_dcpl_535 = (cfg_proc_precision_1_sva_st_102==2'b10);
  assign or_dcpl_181 = or_dcpl_178 | and_dcpl_535;
  assign or_dcpl_184 = (~ and_tmp_165) | and_dcpl_535;
  assign and_1059_cse = (cfg_proc_precision_1_sva_st_108==2'b10);
  assign or_dcpl_188 = (~ and_tmp_165) | and_dcpl_535 | and_1059_cse;
  assign or_dcpl_195 = (~ mux_tmp_986) | and_dcpl_535;
  assign or_dcpl_197 = (~ mux_tmp_986) | and_dcpl_535 | and_1059_cse;
  assign or_dcpl_210 = or_dcpl_195 | and_1059_cse;
  assign mux_1966_itm = MUX_s_1_2_2(cvt_unequal_tmp_21, cvt_unequal_tmp_20, or_5189_cse);
  assign and_dcpl_617 = ((~ mux_tmp_455) | and_1021_cse | (~ main_stage_v_2)) & or_1159_cse
      & or_3538_cse & or_3542_cse & and_dcpl_103;
  assign and_dcpl_626 = or_400_cse_1 & main_stage_v_2;
  assign or_dcpl_243 = and_1021_cse | (~ main_stage_v_2);
  assign and_dcpl_631 = ((~ mux_tmp_455) | or_dcpl_243) & or_1159_cse & or_3538_cse
      & or_3542_cse & and_dcpl_103;
  assign and_dcpl_648 = ((~ and_tmp_225) | or_dcpl_243) & or_1159_cse & or_3538_cse
      & or_3542_cse & or_5254_cse & and_dcpl_103;
  assign or_tmp_3379 = nor_151_cse | nor_2219_cse | nor_50_cse | (~ main_stage_v_2)
      | (cfg_out_precision_1_sva_st_149!=2'b10);
  assign or_dcpl_277 = (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149[0]);
  assign or_dcpl_320 = (~ cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_itm_8_1) |
      cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_itm_7_1 | (~ cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_itm_8_1);
  assign or_dcpl_322 = (~ cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1) |
      cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 | (~ cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1);
  assign or_dcpl_324 = (~ cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1) |
      cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 | (~ cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1);
  assign or_dcpl_326 = (~ cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1) |
      cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1);
  assign or_dcpl_328 = (~ cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1) |
      cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 | (~ cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1);
  assign or_dcpl_330 = (~ cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1) |
      cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1);
  assign or_dcpl_332 = (~ cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1) |
      cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1);
  assign or_dcpl_334 = (~ cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1) | cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1
      | (~ cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1);
  assign or_dcpl_336 = (~ cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1) | cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1
      | (~ cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1);
  assign or_dcpl_338 = (~ cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1) | cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1
      | (~ cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1);
  assign or_dcpl_340 = (~ cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1) | cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1
      | (~ cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1);
  assign or_dcpl_342 = (~ cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1) | cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1
      | (~ cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1);
  assign or_dcpl_344 = (~ cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1) | cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1
      | (~ cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1);
  assign or_dcpl_346 = (~ cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1) | cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1
      | (~ cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1);
  assign or_dcpl_348 = (~ cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1) | cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1
      | (~ cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1);
  assign or_dcpl_350 = (~ cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_itm_8_1)
      | cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1 | (~ cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_itm_8_1);
  assign or_dcpl_353 = (~ and_tmp_50) | and_1021_cse;
  assign or_dcpl_386 = and_dcpl_3 | (~ main_stage_v_1);
  assign or_dcpl_389 = (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_113!=2'b10);
  assign and_dcpl_942 = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_16==5'b00000);
  assign or_dcpl_399 = and_dcpl_93 | (~ main_stage_v_2);
  assign and_dcpl_946 = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_17==5'b00000);
  assign and_dcpl_950 = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_18==5'b00000);
  assign or_dcpl_420 = nand_190_cse | FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_3
      | (cfg_out_precision_1_sva_st_149[0]);
  assign and_dcpl_954 = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_19==5'b00000);
  assign and_dcpl_958 = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_20==5'b00000);
  assign or_dcpl_439 = (~ main_stage_v_2) | FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_3
      | (cfg_out_precision_1_sva_st_149!=2'b10);
  assign and_dcpl_962 = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_21==5'b00000);
  assign or_dcpl_448 = nand_190_cse | FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_3
      | (cfg_out_precision_1_sva_st_149[0]);
  assign and_dcpl_966 = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_22==5'b00000);
  assign and_dcpl_970 = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_23==5'b00000);
  assign and_dcpl_974 = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_24==5'b00000);
  assign or_dcpl_480 = (~ main_stage_v_2) | FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_3;
  assign and_dcpl_978 = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_25==5'b00000);
  assign or_dcpl_490 = nand_190_cse | (cfg_out_precision_1_sva_st_149[0]) | FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_3;
  assign and_dcpl_982 = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_26==5'b00000);
  assign and_dcpl_987 = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_27==5'b00000);
  assign or_dcpl_511 = and_dcpl_93 | and_1021_cse;
  assign and_dcpl_991 = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_28==5'b00000);
  assign and_dcpl_995 = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_29==5'b00000);
  assign and_dcpl_999 = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_30==5'b00000);
  assign and_dcpl_1003 = (libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_31==5'b00000);
  assign or_dcpl_612 = (~ chn_in_rsci_bawt) | (~ (cfg_proc_precision_rsci_d[1]))
      | and_dcpl_93;
  assign or_tmp_3487 = or_5189_cse & chn_in_rsci_bawt & (fsm_output[1]);
  assign chn_in_rsci_ld_core_psct_mx0c0 = main_stage_en_1 | (fsm_output[0]);
  assign main_stage_v_1_mx0c1 = (~ chn_in_rsci_bawt) & main_stage_v_1 & or_5189_cse;
  assign IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1 = (~(cvt_cvt_nand_cse & chn_in_rsci_bawt))
      & or_4550_cse & or_183_cse_1 & and_dcpl_114;
  assign main_stage_v_2_mx0c1 = (~ main_stage_v_1) & main_stage_v_2 & or_5189_cse;
  assign main_stage_v_3_mx0c1 = (~ main_stage_v_2) & main_stage_v_3 & or_5189_cse;
  assign cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c0
      = ((~ cvt_2_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1) | (cfg_out_precision_1_sva_st_149!=2'b01)
      | (cfg_proc_precision_1_sva_st_65!=2'b10)) & and_dcpl_408;
  assign cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c1
      = (~((~ cvt_2_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1) | (cfg_out_precision_1_sva_st_149!=2'b01)))
      & (cfg_proc_precision_1_sva_st_65[1]) & and_dcpl_417;
  assign and_2158_nl = cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1 & nor_45_cse;
  assign mux_1836_nl = MUX_s_1_2_2((~ or_4862_cse), or_4862_cse, and_2158_nl);
  assign cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c0
      = (mux_1836_nl) & and_dcpl_408;
  assign cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c1
      = cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1 & (cfg_proc_precision_1_sva_st_65[1])
      & and_dcpl_417;
  assign and_2157_nl = cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1 & nor_45_cse;
  assign mux_1846_nl = MUX_s_1_2_2((~ or_4862_cse), or_4862_cse, and_2157_nl);
  assign cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0
      = (mux_1846_nl) & and_dcpl_408;
  assign cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1
      = cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1 & (cfg_proc_precision_1_sva_st_65[1])
      & and_dcpl_417;
  assign FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c1 = ((~ and_tmp_50)
      | and_1021_cse | (cfg_out_precision_1_sva_st_113[0])) & and_dcpl_420;
  assign FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c2 = mux_tmp_321 & (~
      (cfg_out_precision_1_sva_st_113[0])) & cvt_unequal_tmp_20 & or_5189_cse;
  assign cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1_mx0c0
      = ((~ cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_itm_11_1) | (cfg_out_precision_1_sva_st_149!=2'b01)
      | (cfg_proc_precision_1_sva_st_65!=2'b10)) & and_dcpl_408;
  assign cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1_mx0c1
      = (~((~ cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_itm_11_1) | (cfg_out_precision_1_sva_st_149!=2'b01)))
      & (cfg_proc_precision_1_sva_st_65[1]) & and_dcpl_417;
  assign and_2155_nl = cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1 & nor_45_cse;
  assign mux_1876_nl = MUX_s_1_2_2((~ or_4862_cse), or_4862_cse, and_2155_nl);
  assign cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0
      = (mux_1876_nl) & and_dcpl_408;
  assign cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1
      = cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1 & (cfg_proc_precision_1_sva_st_65[1])
      & and_dcpl_417;
  assign and_2152_nl = cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1 & nor_45_cse;
  assign mux_1903_nl = MUX_s_1_2_2((~ or_4862_cse), or_4862_cse, and_2152_nl);
  assign cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c0
      = (mux_1903_nl) & and_dcpl_408;
  assign cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c1
      = cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1 & (cfg_proc_precision_1_sva_st_65[1])
      & and_dcpl_417;
  assign and_2150_nl = cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1 & nor_45_cse;
  assign mux_1927_nl = MUX_s_1_2_2((~ or_4862_cse), or_4862_cse, and_2150_nl);
  assign cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0
      = (mux_1927_nl) & and_dcpl_408;
  assign cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1
      = cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1 & (cfg_proc_precision_1_sva_st_65[1])
      & and_dcpl_417;
  assign and_2148_nl = cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1 & nor_45_cse;
  assign mux_1940_nl = MUX_s_1_2_2((~ or_4862_cse), or_4862_cse, and_2148_nl);
  assign cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c0
      = (mux_1940_nl) & and_dcpl_408;
  assign cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c1
      = cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1 & (cfg_proc_precision_1_sva_st_65[1])
      & and_dcpl_417;
  assign and_2147_nl = cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1 & nor_45_cse;
  assign mux_1943_nl = MUX_s_1_2_2((~ or_4862_cse), or_4862_cse, and_2147_nl);
  assign cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c0
      = (mux_1943_nl) & and_dcpl_408;
  assign cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c1
      = cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1 & (cfg_proc_precision_1_sva_st_65[1])
      & and_dcpl_417;
  assign and_2146_nl = cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1 & nor_45_cse;
  assign mux_1953_nl = MUX_s_1_2_2((~ or_4862_cse), or_4862_cse, and_2146_nl);
  assign cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0
      = (mux_1953_nl) & and_dcpl_408;
  assign cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1
      = cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1 & (cfg_proc_precision_1_sva_st_65[1])
      & and_dcpl_417;
  assign and_2145_nl = cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1 & nor_45_cse;
  assign mux_1964_nl = MUX_s_1_2_2((~ or_4862_cse), or_4862_cse, and_2145_nl);
  assign cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0
      = (mux_1964_nl) & and_dcpl_408;
  assign cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1
      = cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1 & (cfg_proc_precision_1_sva_st_65[1])
      & and_dcpl_417;
  assign cvt_1_FpIntToFloat_17U_5U_10U_else_i_abs_conc_3_16 = cvt_1_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_itm_2
      & IntShiftRightSat_49U_6U_17U_o_16_1_sva_3;
  assign cvt_2_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16 = cvt_2_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2
      & IntShiftRightSat_49U_6U_17U_o_16_2_sva_2;
  assign cvt_3_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16 = cvt_3_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2
      & IntShiftRightSat_49U_6U_17U_o_16_3_sva_3;
  assign cvt_4_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16 = cvt_4_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2
      & IntShiftRightSat_49U_6U_17U_o_16_4_sva_2;
  assign cvt_5_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16 = cvt_5_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2
      & IntShiftRightSat_49U_6U_17U_o_16_5_sva_3;
  assign cvt_6_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16 = cvt_6_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2
      & IntShiftRightSat_49U_6U_17U_o_16_6_sva_2;
  assign cvt_7_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16 = cvt_7_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2
      & IntShiftRightSat_49U_6U_17U_o_16_7_sva_2;
  assign cvt_8_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16 = cvt_8_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2
      & IntShiftRightSat_49U_6U_17U_o_16_8_sva_2;
  assign cvt_9_FpIntToFloat_17U_5U_10U_else_i_abs_conc_4_16 = cvt_9_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2
      & IntShiftRightSat_49U_6U_17U_o_16_9_sva_3;
  assign cvt_10_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16 = cvt_10_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2
      & IntShiftRightSat_49U_6U_17U_o_16_10_sva_2;
  assign cvt_11_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16 = cvt_11_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2
      & IntShiftRightSat_49U_6U_17U_o_16_11_sva_2;
  assign cvt_12_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16 = cvt_12_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2
      & IntShiftRightSat_49U_6U_17U_o_16_12_sva_2;
  assign cvt_13_FpIntToFloat_17U_5U_10U_else_i_abs_conc_5_16 = cvt_13_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2
      & IntShiftRightSat_49U_6U_17U_o_16_13_sva_2;
  assign cvt_14_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16 = cvt_14_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2
      & IntShiftRightSat_49U_6U_17U_o_16_14_sva_2;
  assign cvt_15_FpIntToFloat_17U_5U_10U_else_i_abs_conc_6_16 = cvt_15_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2
      & IntShiftRightSat_49U_6U_17U_o_16_15_sva_2;
  assign cvt_16_FpIntToFloat_17U_5U_10U_else_i_abs_conc_7_16 = cvt_16_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_4_itm_2
      & IntShiftRightSat_49U_6U_17U_o_16_sva_2;
  assign or_tmp_3763 = nor_50_cse | nor_2219_cse | nor_151_cse | (cfg_out_precision_1_sva_st_149[0])
      | nand_190_cse;
  assign or_tmp_3768 = nor_50_cse | nor_2219_cse | (cfg_out_precision_1_sva_st_149!=2'b10);
  assign or_tmp_3826 = (cfg_proc_precision_1_sva_st_101[0]) | (fsm_output[1]);
  assign mux_2200_nl = MUX_s_1_2_2((fsm_output[1]), (~ or_5189_cse), cfg_proc_precision_1_sva_st_101[0]);
  assign mux_2201_nl = MUX_s_1_2_2(or_tmp_3826, (mux_2200_nl), main_stage_v_2);
  assign mux_2202_nl = MUX_s_1_2_2(or_tmp_3826, (~ or_5189_cse), main_stage_v_2);
  assign mux_2203_nl = MUX_s_1_2_2((mux_2202_nl), (mux_2201_nl), cfg_proc_precision_1_sva_st_101[1]);
  assign or_4667_nl = nor_151_cse | (cfg_out_precision_1_sva_st_149!=2'b10);
  assign mux_2204_nl = MUX_s_1_2_2((mux_2203_nl), or_tmp_3826, or_4667_nl);
  assign mux_2205_nl = MUX_s_1_2_2((mux_2204_nl), or_tmp_3826, nor_2219_cse);
  assign mux_tmp_2203 = MUX_s_1_2_2((mux_2205_nl), or_tmp_3826, nor_50_cse);
  assign or_tmp_3832 = (~((~ main_stage_v_2) | (cfg_proc_precision_1_sva_st_101[0])
      | (fsm_output[1]))) | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt;
  assign or_4675_nl = (~((~((cfg_out_precision_1_sva_st_149!=2'b10) | (cfg_proc_precision_1_sva_st_101[1])))
      | (~ main_stage_v_2) | (cfg_proc_precision_1_sva_st_101[0]) | (fsm_output[1])))
      | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt;
  assign mux_2207_nl = MUX_s_1_2_2((or_4675_nl), or_tmp_3832, nor_2219_cse);
  assign mux_2208_nl = MUX_s_1_2_2((mux_2207_nl), or_tmp_3832, nor_50_cse);
  assign mux_tmp_2206 = MUX_s_1_2_2((~ mux_tmp_2203), (mux_2208_nl), or_183_cse_1);
  assign or_tmp_3840 = nor_50_cse | nor_2219_cse | (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149[0])
      | (~((cfg_out_precision_1_sva_st_149[1]) & or_400_cse_1));
  assign or_tmp_3849 = nor_50_cse | nor_2219_cse | (cfg_out_precision_1_sva_st_149!=2'b10)
      | (~(main_stage_v_2 & or_400_cse_1));
  assign chn_in_rsci_oswt_unreg = or_tmp_3487;
  assign chn_out_rsci_oswt_unreg = and_dcpl_73;
  assign and_dcpl_1319 = main_stage_v_2 & core_wen;
  assign cvt_and_tmp_1 = (fsm_output[1]) & cvt_unequal_tmp_21;
  assign and_dcpl_1742 = main_stage_v_3 & core_wen;
  assign or_tmp = cvt_else_nor_dfs_2 | FpIntToFloat_17U_5U_10U_is_inf_2_lpi_1_dfm_6
      | cvt_else_equal_tmp_5;
  assign mux_2299_nl = MUX_s_1_2_2(and_2136_cse, (~ or_tmp), cfg_proc_precision_1_sva_st_90[1]);
  assign mux_tmp_2294 = MUX_s_1_2_2((mux_2299_nl), and_2136_cse, cfg_proc_precision_1_sva_st_90[0]);
  assign or_tmp_4080 = cvt_else_nor_dfs_10 | FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_7
      | cvt_else_equal_tmp_9;
  assign mux_2303_nl = MUX_s_1_2_2(and_2136_cse, (~ or_tmp_4080), cfg_proc_precision_1_sva_st_102[1]);
  assign mux_tmp_2298 = MUX_s_1_2_2((mux_2303_nl), and_2136_cse, cfg_proc_precision_1_sva_st_102[0]);
  assign mux_2305_nl = MUX_s_1_2_2(mux_tmp_2298, (~ or_tmp_4080), cfg_proc_precision_1_sva_st_90[1]);
  assign mux_tmp_2300 = MUX_s_1_2_2((mux_2305_nl), mux_tmp_2298, cfg_proc_precision_1_sva_st_90[0]);
  assign or_tmp_4081 = cvt_else_nor_dfs_10 | FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_7
      | cvt_else_equal_tmp_16;
  assign mux_2309_nl = MUX_s_1_2_2(and_2136_cse, (~ or_tmp_4081), cfg_proc_precision_1_sva_st_102[1]);
  assign mux_tmp_2304 = MUX_s_1_2_2((mux_2309_nl), and_2136_cse, cfg_proc_precision_1_sva_st_102[0]);
  assign mux_2311_nl = MUX_s_1_2_2(mux_tmp_2304, (~ or_tmp_4081), cfg_proc_precision_1_sva_st_66[1]);
  assign mux_tmp_2306 = MUX_s_1_2_2((mux_2311_nl), mux_tmp_2304, cfg_proc_precision_1_sva_st_66[0]);
  assign or_tmp_4082 = cvt_else_nor_dfs_10 | FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_7
      | FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_8;
  assign mux_2315_nl = MUX_s_1_2_2(and_2136_cse, (~ or_tmp_4082), cfg_proc_precision_1_sva_st_66[1]);
  assign mux_tmp_2310 = MUX_s_1_2_2((mux_2315_nl), and_2136_cse, cfg_proc_precision_1_sva_st_66[0]);
  assign mux_2317_nl = MUX_s_1_2_2(mux_tmp_2310, (~ or_tmp_4082), cfg_proc_precision_1_sva_st_90[1]);
  assign mux_tmp_2312 = MUX_s_1_2_2((mux_2317_nl), mux_tmp_2310, cfg_proc_precision_1_sva_st_90[0]);
  assign or_tmp_4084 = cvt_else_nor_dfs_11 | cvt_else_equal_tmp_33 | cvt_else_equal_tmp_34;
  assign mux_tmp_2315 = MUX_s_1_2_2((~ or_tmp_4084), and_2136_cse, or_5254_cse);
  assign mux_2322_nl = MUX_s_1_2_2(mux_tmp_2315, (~ or_tmp_4084), cfg_proc_precision_1_sva_st_102[1]);
  assign mux_tmp_2317 = MUX_s_1_2_2((mux_2322_nl), mux_tmp_2315, cfg_proc_precision_1_sva_st_102[0]);
  assign mux_2324_nl = MUX_s_1_2_2(mux_tmp_2317, (~ or_tmp_4084), cfg_proc_precision_1_sva_st_66[1]);
  assign mux_tmp_2319 = MUX_s_1_2_2((mux_2324_nl), mux_tmp_2317, cfg_proc_precision_1_sva_st_66[0]);
  assign or_tmp_4086 = reg_cvt_else_nor_dfs_9_cse | FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_7
      | cvt_else_equal_tmp_28;
  assign mux_tmp_2322 = MUX_s_1_2_2((~ or_tmp_4086), and_2136_cse, or_3542_cse);
  assign mux_2329_nl = MUX_s_1_2_2(mux_tmp_2322, (~ or_tmp_4086), cfg_proc_precision_1_sva_st_66[1]);
  assign mux_tmp_2324 = MUX_s_1_2_2((mux_2329_nl), mux_tmp_2322, cfg_proc_precision_1_sva_st_66[0]);
  assign or_tmp_4087 = cvt_else_nor_dfs_10 | FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_7
      | FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_8;
  assign mux_2333_nl = MUX_s_1_2_2(and_2136_cse, (~ or_tmp_4087), cfg_proc_precision_1_sva_st_66[1]);
  assign mux_tmp_2328 = MUX_s_1_2_2((mux_2333_nl), and_2136_cse, cfg_proc_precision_1_sva_st_66[0]);
  assign mux_2335_nl = MUX_s_1_2_2(mux_tmp_2328, (~ or_tmp_4087), cfg_proc_precision_1_sva_st_90[1]);
  assign mux_tmp_2330 = MUX_s_1_2_2((mux_2335_nl), mux_tmp_2328, cfg_proc_precision_1_sva_st_90[0]);
  assign mux_tmp_2334 = MUX_s_1_2_2((~ or_tmp_4084), mux_tmp_2315, or_3542_cse);
  assign mux_2341_nl = MUX_s_1_2_2(mux_tmp_2334, (~ or_tmp_4084), cfg_proc_precision_1_sva_st_66[1]);
  assign mux_tmp_2336 = MUX_s_1_2_2((mux_2341_nl), mux_tmp_2334, cfg_proc_precision_1_sva_st_66[0]);
  assign or_tmp_4092 = reg_cvt_else_nor_dfs_9_cse | FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_7
      | FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_8;
  assign mux_tmp_2339 = MUX_s_1_2_2((~ or_tmp_4092), and_2136_cse, or_3542_cse);
  assign mux_2346_nl = MUX_s_1_2_2(mux_tmp_2339, (~ or_tmp_4092), cfg_proc_precision_1_sva_st_66[1]);
  assign mux_tmp_2341 = MUX_s_1_2_2((mux_2346_nl), mux_tmp_2339, cfg_proc_precision_1_sva_st_66[0]);
  assign or_tmp_4095 = cvt_else_nor_dfs_15 | cvt_else_equal_tmp_45 | cvt_else_equal_tmp_46;
  assign mux_2350_nl = MUX_s_1_2_2((~ or_tmp_4095), and_2136_cse, or_5254_cse);
  assign mux_tmp_2345 = MUX_s_1_2_2((~ or_tmp_4095), (mux_2350_nl), or_3542_cse);
  assign mux_2352_nl = MUX_s_1_2_2(mux_tmp_2345, (~ or_tmp_4095), cfg_proc_precision_1_sva_st_66[1]);
  assign mux_tmp_2347 = MUX_s_1_2_2((mux_2352_nl), mux_tmp_2345, cfg_proc_precision_1_sva_st_66[0]);
  assign or_tmp_4097 = cvt_else_nor_dfs_15 | FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_8
      | FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_9;
  assign mux_2356_nl = MUX_s_1_2_2(and_2136_cse, (~ or_tmp_4097), cfg_proc_precision_1_sva_st_66[1]);
  assign mux_tmp_2351 = MUX_s_1_2_2((mux_2356_nl), and_2136_cse, cfg_proc_precision_1_sva_st_66[0]);
  assign mux_2358_nl = MUX_s_1_2_2(mux_tmp_2351, (~ or_tmp_4097), cfg_proc_precision_1_sva_st_90[1]);
  assign mux_tmp_2353 = MUX_s_1_2_2((mux_2358_nl), mux_tmp_2351, cfg_proc_precision_1_sva_st_90[0]);
  assign or_tmp_4102 = (cvt_asn_323 & (~ FpIntToFloat_17U_5U_10U_is_inf_1_lpi_1_dfm_6)
      & (~ IsNaN_5U_10U_land_2_lpi_1_dfm_4)) | cvt_asn_321;
  assign or_5174_tmp = (cvt_asn_329 & (~ FpIntToFloat_17U_5U_10U_is_inf_2_lpi_1_dfm_6)
      & (~ IsNaN_5U_10U_land_3_lpi_1_dfm_5)) | cvt_asn_321;
  assign or_5175_tmp = (cvt_asn_323 & (~ FpIntToFloat_17U_5U_10U_is_inf_3_lpi_1_dfm_7)
      & (~ IsNaN_5U_10U_land_4_lpi_1_dfm_5)) | cvt_asn_321;
  assign or_5176_tmp = (cvt_asn_335 & (~ FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_7)
      & (~ IsNaN_5U_10U_land_5_lpi_1_dfm_5)) | cvt_asn_321;
  assign or_5177_tmp = (cvt_asn_323 & (~ FpIntToFloat_17U_5U_10U_is_inf_5_lpi_1_dfm_7)
      & (~ IsNaN_5U_10U_land_6_lpi_1_dfm_5)) | cvt_asn_321;
  assign or_5178_tmp = (cvt_asn_353 & (~ FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_7)
      & (~ IsNaN_5U_10U_land_7_lpi_1_dfm_6)) | cvt_asn_321;
  assign or_5179_tmp = (cvt_asn_365 & (~ FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_7)
      & (~ IsNaN_5U_10U_land_8_lpi_1_dfm_5)) | cvt_asn_321;
  assign or_5180_tmp = (cvt_asn_377 & (~ FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_8)
      & (~ IsNaN_5U_10U_land_9_lpi_1_dfm_5)) | cvt_asn_321;
  assign or_5181_tmp = (cvt_asn_323 & (~ FpIntToFloat_17U_5U_10U_is_inf_9_lpi_1_dfm_7)
      & (~ IsNaN_5U_10U_land_lpi_1_dfm_5)) | cvt_asn_321;
  assign or_5182_tmp = (cvt_asn_371 & (~ FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_7)
      & (~ IsNaN_5U_10U_land_1_lpi_1_dfm_3)) | cvt_asn_321;
  assign or_5183_tmp = (cvt_asn_389 & (~ FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_7)
      & (~ IsNaN_5U_10U_land_10_lpi_1_dfm_5)) | cvt_asn_321;
  assign or_5184_tmp = (cvt_asn_383 & (~ FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_8)
      & (~ IsNaN_5U_10U_land_11_lpi_1_dfm_5)) | cvt_asn_321;
  assign or_5185_tmp = (cvt_asn_371 & (~ FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_7)
      & (~ IsNaN_5U_10U_land_12_lpi_1_dfm_5)) | cvt_asn_321;
  assign or_5186_tmp = (cvt_asn_359 & (~ FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_8)
      & (~ IsNaN_5U_10U_land_13_lpi_1_dfm_5)) | cvt_asn_321;
  assign or_5187_tmp = (cvt_asn_347 & (~ FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_8)
      & (~ IsNaN_5U_10U_land_14_lpi_1_dfm_6)) | cvt_asn_321;
  assign or_5188_tmp = (cvt_asn_341 & (~ FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_9)
      & (~ IsNaN_5U_10U_land_15_lpi_1_dfm_3)) | cvt_asn_321;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_in_rsci_iswt0 <= 1'b0;
      chn_out_rsci_iswt0 <= 1'b0;
    end
    else if ( core_wen ) begin
      chn_in_rsci_iswt0 <= ~((~ main_stage_en_1) & (fsm_output[1]));
      chn_out_rsci_iswt0 <= and_dcpl_103;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_in_rsci_ld_core_psct <= 1'b0;
    end
    else if ( core_wen & chn_in_rsci_ld_core_psct_mx0c0 ) begin
      chn_in_rsci_ld_core_psct <= chn_in_rsci_ld_core_psct_mx0c0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_out_rsci_d_13_10 <= 4'b0;
      chn_out_rsci_d_45_42 <= 4'b0;
      chn_out_rsci_d_77_74 <= 4'b0;
      chn_out_rsci_d_141_138 <= 4'b0;
    end
    else if ( and_3024_cse ) begin
      chn_out_rsci_d_13_10 <= MUX1HOT_v_4_6_2(({(reg_chn_idata_data_sva_3_15_0_1_reg[2:0])
          , (reg_chn_idata_data_sva_3_15_0_2_reg[9])}), (reg_chn_idata_data_sva_3_15_0_1_reg[3:0]),
          (signext_4_1(~ IsNaN_5U_10U_land_2_lpi_1_dfm_4)), 4'b1110, (signext_4_1(IntSaturation_17U_8U_o_7_1_1_lpi_1_dfm_1[6])),
          reg_FpIntToFloat_17U_5U_10U_o_expo_1_lpi_1_dfm_7_1_itm, {cvt_or_cse , cfg_mode_eql_1_sva_6
          , (cvt_and_261_nl) , (cvt_and_262_nl) , cvt_asn_327 , or_tmp_4102});
      chn_out_rsci_d_45_42 <= MUX1HOT_v_4_6_2(({(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_reg[2:0])
          , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_1_reg[9])}), (chn_idata_data_sva_3_79_63_1[14:11]),
          (signext_4_1(~ IsNaN_5U_10U_land_4_lpi_1_dfm_5)), 4'b1110, (signext_4_1(IntSaturation_17U_8U_o_7_1_3_lpi_1_dfm_1[6])),
          reg_FpIntToFloat_17U_5U_10U_o_expo_3_lpi_1_dfm_8_1_itm, {cvt_or_cse , cfg_mode_eql_1_sva_6
          , (cvt_and_257_nl) , (cvt_and_258_nl) , cvt_asn_327 , or_5175_tmp});
      chn_out_rsci_d_77_74 <= MUX1HOT_v_4_6_2(({(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_reg[2:0])
          , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_1_reg[9])}), (chn_idata_data_sva_3_143_127_1[14:11]),
          (signext_4_1(~ IsNaN_5U_10U_land_6_lpi_1_dfm_5)), 4'b1110, (signext_4_1(IntSaturation_17U_8U_o_7_1_5_lpi_1_dfm_1[6])),
          reg_FpIntToFloat_17U_5U_10U_o_expo_5_lpi_1_dfm_8_1_itm, {cvt_or_cse , cfg_mode_eql_1_sva_6
          , (cvt_and_253_nl) , (cvt_and_254_nl) , cvt_asn_327 , or_5177_tmp});
      chn_out_rsci_d_141_138 <= MUX1HOT_v_4_6_2(({(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_reg[2:0])
          , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_1_reg[9])}), (chn_idata_data_sva_3_271_255_1[14:11]),
          (signext_4_1(~ IsNaN_5U_10U_land_lpi_1_dfm_5)), 4'b1110, (signext_4_1(IntSaturation_17U_8U_o_7_1_9_lpi_1_dfm_1[6])),
          reg_FpIntToFloat_17U_5U_10U_o_expo_9_lpi_1_dfm_8_1_itm, {cvt_or_cse , cfg_mode_eql_1_sva_6
          , (cvt_and_245_nl) , (cvt_and_246_nl) , cvt_asn_327 , or_5181_tmp});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_out_rsci_d_14 <= 1'b0;
      chn_out_rsci_d_30 <= 1'b0;
      chn_out_rsci_d_46 <= 1'b0;
      chn_out_rsci_d_62 <= 1'b0;
      chn_out_rsci_d_78 <= 1'b0;
      chn_out_rsci_d_94 <= 1'b0;
      chn_out_rsci_d_110 <= 1'b0;
      chn_out_rsci_d_126 <= 1'b0;
      chn_out_rsci_d_142 <= 1'b0;
      chn_out_rsci_d_158 <= 1'b0;
      chn_out_rsci_d_174 <= 1'b0;
      chn_out_rsci_d_190 <= 1'b0;
      chn_out_rsci_d_206 <= 1'b0;
      chn_out_rsci_d_222 <= 1'b0;
      chn_out_rsci_d_238 <= 1'b0;
      chn_out_rsci_d_254 <= 1'b0;
      chn_out_rsci_d_9_1 <= 9'b0;
      chn_out_rsci_d_25_17 <= 9'b0;
      chn_out_rsci_d_41_33 <= 9'b0;
      chn_out_rsci_d_57_49 <= 9'b0;
      chn_out_rsci_d_73_65 <= 9'b0;
      chn_out_rsci_d_89_81 <= 9'b0;
      chn_out_rsci_d_105_97 <= 9'b0;
      chn_out_rsci_d_121_113 <= 9'b0;
      chn_out_rsci_d_137_129 <= 9'b0;
      chn_out_rsci_d_153_145 <= 9'b0;
      chn_out_rsci_d_169_161 <= 9'b0;
      chn_out_rsci_d_185_177 <= 9'b0;
      chn_out_rsci_d_201_193 <= 9'b0;
      chn_out_rsci_d_217_209 <= 9'b0;
      chn_out_rsci_d_233_225 <= 9'b0;
      chn_out_rsci_d_249_241 <= 9'b0;
      chn_out_rsci_d_256 <= 1'b0;
      chn_out_rsci_d_257 <= 1'b0;
      chn_out_rsci_d_258 <= 1'b0;
      chn_out_rsci_d_259 <= 1'b0;
      chn_out_rsci_d_260 <= 1'b0;
      chn_out_rsci_d_261 <= 1'b0;
      chn_out_rsci_d_262 <= 1'b0;
      chn_out_rsci_d_263 <= 1'b0;
      chn_out_rsci_d_264 <= 1'b0;
      chn_out_rsci_d_265 <= 1'b0;
      chn_out_rsci_d_266 <= 1'b0;
      chn_out_rsci_d_267 <= 1'b0;
      chn_out_rsci_d_268 <= 1'b0;
      chn_out_rsci_d_269 <= 1'b0;
      chn_out_rsci_d_270 <= 1'b0;
      chn_out_rsci_d_271 <= 1'b0;
    end
    else if ( chn_out_and_cse ) begin
      chn_out_rsci_d_14 <= MUX1HOT_s_1_5_2((reg_chn_idata_data_sva_3_15_0_1_reg[3]),
          FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_2, (reg_chn_idata_data_sva_3_15_0_1_reg[4]),
          (SetToInf_5U_10U_SetToInf_5U_10U_or_nl), (IntSaturation_17U_8U_o_7_1_1_lpi_1_dfm_1[6]),
          {cvt_or_cse , cvt_asn_321 , cfg_mode_eql_1_sva_6 , cvt_asn_323 , cvt_asn_327});
      chn_out_rsci_d_30 <= MUX1HOT_s_1_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_reg[3]),
          FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_2, (chn_idata_data_sva_3_47_31_1[15]),
          (SetToInf_5U_10U_SetToInf_5U_10U_or_1_nl), (IntSaturation_17U_8U_o_7_1_2_lpi_1_dfm_1[6]),
          {cvt_or_2_cse , cvt_asn_321 , cfg_mode_eql_1_sva_6 , cvt_asn_329 , cvt_asn_333});
      chn_out_rsci_d_46 <= MUX1HOT_s_1_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_reg[3]),
          FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_2, (chn_idata_data_sva_3_79_63_1[15]),
          (SetToInf_5U_10U_SetToInf_5U_10U_or_2_nl), (IntSaturation_17U_8U_o_7_1_3_lpi_1_dfm_1[6]),
          {cvt_or_cse , cvt_asn_321 , cfg_mode_eql_1_sva_6 , cvt_asn_323 , cvt_asn_327});
      chn_out_rsci_d_62 <= MUX1HOT_s_1_5_2((FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5[13]),
          FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_2, (chn_idata_data_sva_3_111_95_1[15]),
          (SetToInf_5U_10U_SetToInf_5U_10U_or_3_nl), (IntSaturation_17U_8U_o_7_1_4_lpi_1_dfm_1[6]),
          {cvt_or_6_cse , cvt_asn_321 , cfg_mode_eql_1_sva_6 , cvt_asn_335 , cvt_asn_339});
      chn_out_rsci_d_78 <= MUX1HOT_s_1_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_reg[3]),
          FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_2, (chn_idata_data_sva_3_143_127_1[15]),
          (SetToInf_5U_10U_SetToInf_5U_10U_or_4_nl), (IntSaturation_17U_8U_o_7_1_5_lpi_1_dfm_1[6]),
          {cvt_or_cse , cvt_asn_321 , cfg_mode_eql_1_sva_6 , cvt_asn_323 , cvt_asn_327});
      chn_out_rsci_d_94 <= MUX1HOT_s_1_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_reg[3]),
          FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_2, (chn_idata_data_sva_3_175_159_1[15]),
          (SetToInf_5U_10U_SetToInf_5U_10U_or_5_nl), (IntSaturation_17U_8U_o_7_1_6_lpi_1_dfm_1[6]),
          {cvt_or_10_cse , cvt_asn_321 , cfg_mode_eql_1_sva_6 , cvt_asn_353 , cvt_asn_357});
      chn_out_rsci_d_110 <= MUX1HOT_s_1_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_reg[3]),
          FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_2, (chn_idata_data_sva_3_207_191_1[15]),
          (SetToInf_5U_10U_SetToInf_5U_10U_or_6_nl), (IntSaturation_17U_8U_o_7_1_7_lpi_1_dfm_1[6]),
          {cvt_or_12_cse , cvt_asn_321 , cfg_mode_eql_1_sva_6 , cvt_asn_365 , cvt_asn_369});
      chn_out_rsci_d_126 <= MUX1HOT_s_1_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_reg[3]),
          FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_2, (chn_idata_data_sva_3_239_223_1[15]),
          (SetToInf_5U_10U_SetToInf_5U_10U_or_7_nl), (IntSaturation_17U_8U_o_7_1_8_lpi_1_dfm_1[6]),
          {cvt_or_14_cse , cvt_asn_321 , cfg_mode_eql_1_sva_6 , cvt_asn_377 , cvt_asn_381});
      chn_out_rsci_d_142 <= MUX1HOT_s_1_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_reg[3]),
          FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_2, (chn_idata_data_sva_3_271_255_1[15]),
          (SetToInf_5U_10U_SetToInf_5U_10U_or_8_nl), (IntSaturation_17U_8U_o_7_1_9_lpi_1_dfm_1[6]),
          {cvt_or_cse , cvt_asn_321 , cfg_mode_eql_1_sva_6 , cvt_asn_323 , cvt_asn_327});
      chn_out_rsci_d_158 <= MUX1HOT_s_1_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_reg[3]),
          FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_2, (chn_idata_data_sva_3_303_287_1[15]),
          (SetToInf_5U_10U_SetToInf_5U_10U_or_9_nl), (IntSaturation_17U_8U_o_7_1_10_lpi_1_dfm_1[6]),
          {cvt_or_18_cse , cvt_asn_321 , cfg_mode_eql_1_sva_6 , cvt_asn_371 , cvt_asn_399});
      chn_out_rsci_d_174 <= MUX1HOT_s_1_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_reg[3]),
          FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_2, (chn_idata_data_sva_3_335_319_1[15]),
          (SetToInf_5U_10U_SetToInf_5U_10U_or_10_nl), (IntSaturation_17U_8U_o_7_1_11_lpi_1_dfm_1[6]),
          {cvt_or_20_cse , cvt_asn_321 , cfg_mode_eql_1_sva_6 , cvt_asn_389 , cvt_asn_393});
      chn_out_rsci_d_190 <= MUX1HOT_s_1_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_reg[3]),
          FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_2, (chn_idata_data_sva_3_367_351_1[15]),
          (SetToInf_5U_10U_SetToInf_5U_10U_or_11_nl), (IntSaturation_17U_8U_o_7_1_12_lpi_1_dfm_1[6]),
          {cvt_or_22_cse , cvt_asn_321 , cfg_mode_eql_1_sva_6 , cvt_asn_383 , cvt_asn_387});
      chn_out_rsci_d_206 <= MUX1HOT_s_1_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_reg[3]),
          FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_2, (chn_idata_data_sva_3_399_383_1[15]),
          (SetToInf_5U_10U_SetToInf_5U_10U_or_12_nl), (IntSaturation_17U_8U_o_7_1_13_lpi_1_dfm_1[6]),
          {cvt_or_24_cse , cvt_asn_321 , cfg_mode_eql_1_sva_6 , cvt_asn_371 , cvt_asn_375});
      chn_out_rsci_d_222 <= MUX1HOT_s_1_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_reg[3]),
          FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_2, (chn_idata_data_sva_3_431_415_1[15]),
          (SetToInf_5U_10U_SetToInf_5U_10U_or_13_nl), (IntSaturation_17U_8U_o_7_1_14_lpi_1_dfm_1[6]),
          {cvt_or_26_cse , cvt_asn_321 , cfg_mode_eql_1_sva_6 , cvt_asn_359 , cvt_asn_363});
      chn_out_rsci_d_238 <= MUX1HOT_s_1_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_reg[3]),
          FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_2, (chn_idata_data_sva_3_463_447_1[15]),
          (SetToInf_5U_10U_SetToInf_5U_10U_or_14_nl), (IntSaturation_17U_8U_o_7_1_15_lpi_1_dfm_1[6]),
          {cvt_or_28_cse , cvt_asn_321 , cfg_mode_eql_1_sva_6 , cvt_asn_347 , cvt_asn_351});
      chn_out_rsci_d_254 <= MUX1HOT_s_1_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_reg[3]),
          FpFloatToInt_16U_5U_10U_internal_int_0_sva_3, (SetToInf_5U_10U_SetToInf_5U_10U_or_15_nl),
          (IntSaturation_17U_8U_o_7_1_lpi_1_dfm_1[6]), (chn_idata_data_sva_3_495_479_1[15]),
          {cvt_or_30_cse , cvt_asn_321 , cvt_asn_341 , cvt_asn_345 , cfg_mode_eql_1_sva_6});
      chn_out_rsci_d_9_1 <= MUX1HOT_v_9_4_2((reg_chn_idata_data_sva_3_15_0_2_reg[8:0]),
          (reg_chn_idata_data_sva_3_15_0_2_reg[9:1]), (FpIntToFloat_17U_5U_10U_o_mant_1_lpi_1_dfm_1[9:1]),
          ({{2{IntSaturation_17U_8U_o_7_1_1_lpi_1_dfm_1[6]}}, IntSaturation_17U_8U_o_7_1_1_lpi_1_dfm_1}),
          {cvt_or_cse , (cvt_or_48_nl) , cvt_asn_323 , cvt_asn_327});
      chn_out_rsci_d_25_17 <= MUX1HOT_v_9_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_1_reg[8:0]),
          (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_1_reg[9:1]), (chn_idata_data_sva_3_47_31_1[10:2]),
          (FpIntToFloat_17U_5U_10U_o_mant_2_lpi_1_dfm_1[9:1]), ({{2{IntSaturation_17U_8U_o_7_1_2_lpi_1_dfm_1[6]}},
          IntSaturation_17U_8U_o_7_1_2_lpi_1_dfm_1}), {cvt_or_2_cse , cvt_asn_321
          , cfg_mode_eql_1_sva_6 , cvt_asn_329 , cvt_asn_333});
      chn_out_rsci_d_41_33 <= MUX1HOT_v_9_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_1_reg[8:0]),
          (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_1_reg[9:1]), (chn_idata_data_sva_3_79_63_1[10:2]),
          (FpIntToFloat_17U_5U_10U_o_mant_3_lpi_1_dfm_1[9:1]), ({{2{IntSaturation_17U_8U_o_7_1_3_lpi_1_dfm_1[6]}},
          IntSaturation_17U_8U_o_7_1_3_lpi_1_dfm_1}), {cvt_or_cse , cvt_asn_321 ,
          cfg_mode_eql_1_sva_6 , cvt_asn_323 , cvt_asn_327});
      chn_out_rsci_d_57_49 <= MUX1HOT_v_9_5_2((FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5[8:0]),
          (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_1_reg[9:1]), (chn_idata_data_sva_3_111_95_1[10:2]),
          (FpIntToFloat_17U_5U_10U_o_mant_4_lpi_1_dfm_1[9:1]), ({{2{IntSaturation_17U_8U_o_7_1_4_lpi_1_dfm_1[6]}},
          IntSaturation_17U_8U_o_7_1_4_lpi_1_dfm_1}), {cvt_or_6_cse , cvt_asn_321
          , cfg_mode_eql_1_sva_6 , cvt_asn_335 , cvt_asn_339});
      chn_out_rsci_d_73_65 <= MUX1HOT_v_9_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_1_reg[8:0]),
          (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_1_reg[9:1]), (chn_idata_data_sva_3_143_127_1[10:2]),
          (FpIntToFloat_17U_5U_10U_o_mant_5_lpi_1_dfm_1[9:1]), ({{2{IntSaturation_17U_8U_o_7_1_5_lpi_1_dfm_1[6]}},
          IntSaturation_17U_8U_o_7_1_5_lpi_1_dfm_1}), {cvt_or_cse , cvt_asn_321 ,
          cfg_mode_eql_1_sva_6 , cvt_asn_323 , cvt_asn_327});
      chn_out_rsci_d_89_81 <= MUX1HOT_v_9_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_1_reg[8:0]),
          (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_1_reg[9:1]), (chn_idata_data_sva_3_175_159_1[10:2]),
          (FpIntToFloat_17U_5U_10U_o_mant_6_lpi_1_dfm_1[9:1]), ({{2{IntSaturation_17U_8U_o_7_1_6_lpi_1_dfm_1[6]}},
          IntSaturation_17U_8U_o_7_1_6_lpi_1_dfm_1}), {cvt_or_10_cse , cvt_asn_321
          , cfg_mode_eql_1_sva_6 , cvt_asn_353 , cvt_asn_357});
      chn_out_rsci_d_105_97 <= MUX1HOT_v_9_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_1_reg[8:0]),
          (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_1_reg[9:1]), (chn_idata_data_sva_3_207_191_1[10:2]),
          (FpIntToFloat_17U_5U_10U_o_mant_7_lpi_1_dfm_1[9:1]), ({{2{IntSaturation_17U_8U_o_7_1_7_lpi_1_dfm_1[6]}},
          IntSaturation_17U_8U_o_7_1_7_lpi_1_dfm_1}), {cvt_or_12_cse , cvt_asn_321
          , cfg_mode_eql_1_sva_6 , cvt_asn_365 , cvt_asn_369});
      chn_out_rsci_d_121_113 <= MUX1HOT_v_9_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_1_reg[8:0]),
          (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_1_reg[9:1]), (chn_idata_data_sva_3_239_223_1[10:2]),
          (FpIntToFloat_17U_5U_10U_o_mant_8_lpi_1_dfm_1[9:1]), ({{2{IntSaturation_17U_8U_o_7_1_8_lpi_1_dfm_1[6]}},
          IntSaturation_17U_8U_o_7_1_8_lpi_1_dfm_1}), {cvt_or_14_cse , cvt_asn_321
          , cfg_mode_eql_1_sva_6 , cvt_asn_377 , cvt_asn_381});
      chn_out_rsci_d_137_129 <= MUX1HOT_v_9_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_1_reg[8:0]),
          (FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_7_itm_1[9:1]), (chn_idata_data_sva_3_271_255_1[10:2]),
          (FpIntToFloat_17U_5U_10U_o_mant_9_lpi_1_dfm_1[9:1]), ({{2{IntSaturation_17U_8U_o_7_1_9_lpi_1_dfm_1[6]}},
          IntSaturation_17U_8U_o_7_1_9_lpi_1_dfm_1}), {cvt_or_cse , cvt_asn_321 ,
          cfg_mode_eql_1_sva_6 , cvt_asn_323 , cvt_asn_327});
      chn_out_rsci_d_153_145 <= MUX1HOT_v_9_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_1_reg[8:0]),
          (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_1_reg[9:1]), (chn_idata_data_sva_3_303_287_1[10:2]),
          (FpIntToFloat_17U_5U_10U_o_mant_10_lpi_1_dfm_1[9:1]), ({{2{IntSaturation_17U_8U_o_7_1_10_lpi_1_dfm_1[6]}},
          IntSaturation_17U_8U_o_7_1_10_lpi_1_dfm_1}), {cvt_or_18_cse , cvt_asn_321
          , cfg_mode_eql_1_sva_6 , cvt_asn_371 , cvt_asn_399});
      chn_out_rsci_d_169_161 <= MUX1HOT_v_9_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_1_reg[8:0]),
          (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_1_reg[9:1]), (chn_idata_data_sva_3_335_319_1[10:2]),
          (FpIntToFloat_17U_5U_10U_o_mant_11_lpi_1_dfm_1[9:1]), ({{2{IntSaturation_17U_8U_o_7_1_11_lpi_1_dfm_1[6]}},
          IntSaturation_17U_8U_o_7_1_11_lpi_1_dfm_1}), {cvt_or_20_cse , cvt_asn_321
          , cfg_mode_eql_1_sva_6 , cvt_asn_389 , cvt_asn_393});
      chn_out_rsci_d_185_177 <= MUX1HOT_v_9_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_1_reg[8:0]),
          (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_1_reg[9:1]), (chn_idata_data_sva_3_367_351_1[10:2]),
          (FpIntToFloat_17U_5U_10U_o_mant_12_lpi_1_dfm_1[9:1]), ({{2{IntSaturation_17U_8U_o_7_1_12_lpi_1_dfm_1[6]}},
          IntSaturation_17U_8U_o_7_1_12_lpi_1_dfm_1}), {cvt_or_22_cse , cvt_asn_321
          , cfg_mode_eql_1_sva_6 , cvt_asn_383 , cvt_asn_387});
      chn_out_rsci_d_201_193 <= MUX1HOT_v_9_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_1_reg[8:0]),
          (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_1_reg[9:1]), (chn_idata_data_sva_3_399_383_1[10:2]),
          (FpIntToFloat_17U_5U_10U_o_mant_13_lpi_1_dfm_1[9:1]), ({{2{IntSaturation_17U_8U_o_7_1_13_lpi_1_dfm_1[6]}},
          IntSaturation_17U_8U_o_7_1_13_lpi_1_dfm_1}), {cvt_or_24_cse , cvt_asn_321
          , cfg_mode_eql_1_sva_6 , cvt_asn_371 , cvt_asn_375});
      chn_out_rsci_d_217_209 <= MUX1HOT_v_9_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_1_reg[8:0]),
          (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_1_reg[9:1]), (chn_idata_data_sva_3_431_415_1[10:2]),
          (FpIntToFloat_17U_5U_10U_o_mant_14_lpi_1_dfm_1[9:1]), ({{2{IntSaturation_17U_8U_o_7_1_14_lpi_1_dfm_1[6]}},
          IntSaturation_17U_8U_o_7_1_14_lpi_1_dfm_1}), {cvt_or_26_cse , cvt_asn_321
          , cfg_mode_eql_1_sva_6 , cvt_asn_359 , cvt_asn_363});
      chn_out_rsci_d_233_225 <= MUX1HOT_v_9_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_1_reg[8:0]),
          (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_1_reg[9:1]), (chn_idata_data_sva_3_463_447_1[10:2]),
          (FpIntToFloat_17U_5U_10U_o_mant_15_lpi_1_dfm_1[9:1]), ({{2{IntSaturation_17U_8U_o_7_1_15_lpi_1_dfm_1[6]}},
          IntSaturation_17U_8U_o_7_1_15_lpi_1_dfm_1}), {cvt_or_28_cse , cvt_asn_321
          , cfg_mode_eql_1_sva_6 , cvt_asn_347 , cvt_asn_351});
      chn_out_rsci_d_249_241 <= MUX1HOT_v_9_5_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_1_reg[8:0]),
          (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_1_reg[9:1]), (FpIntToFloat_17U_5U_10U_o_mant_lpi_1_dfm_1[9:1]),
          ({{2{IntSaturation_17U_8U_o_7_1_lpi_1_dfm_1[6]}}, IntSaturation_17U_8U_o_7_1_lpi_1_dfm_1}),
          (chn_idata_data_sva_3_495_479_1[10:2]), {cvt_or_30_cse , cvt_asn_321 ,
          cvt_asn_341 , cvt_asn_345 , cfg_mode_eql_1_sva_6});
      chn_out_rsci_d_256 <= cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          & cvt_unequal_tmp_21;
      chn_out_rsci_d_257 <= cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          & cvt_unequal_tmp_21;
      chn_out_rsci_d_258 <= cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          & cvt_unequal_tmp_21;
      chn_out_rsci_d_259 <= cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          & cvt_unequal_tmp_21;
      chn_out_rsci_d_260 <= cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          & cvt_unequal_tmp_21;
      chn_out_rsci_d_261 <= cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          & cvt_unequal_tmp_21;
      chn_out_rsci_d_262 <= cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          & cvt_unequal_tmp_21;
      chn_out_rsci_d_263 <= cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          & cvt_unequal_tmp_21;
      chn_out_rsci_d_264 <= cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          & cvt_unequal_tmp_21;
      chn_out_rsci_d_265 <= cvt_10_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          & cvt_unequal_tmp_21;
      chn_out_rsci_d_266 <= cvt_11_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          & cvt_unequal_tmp_21;
      chn_out_rsci_d_267 <= cvt_12_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          & cvt_unequal_tmp_21;
      chn_out_rsci_d_268 <= cvt_13_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          & cvt_unequal_tmp_21;
      chn_out_rsci_d_269 <= cvt_14_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          & cvt_unequal_tmp_21;
      chn_out_rsci_d_270 <= cvt_15_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          & cvt_unequal_tmp_21;
      chn_out_rsci_d_271 <= cvt_16_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          & cvt_unequal_tmp_21;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_out_rsci_d_29_26 <= 4'b0;
    end
    else if ( ((~ (mux_2302_nl)) | (~ cvt_unequal_tmp_21) | cfg_mode_eql_1_sva_6)
        & or_5189_cse & and_dcpl_1742 ) begin
      chn_out_rsci_d_29_26 <= MUX1HOT_v_4_6_2(({(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_reg[2:0])
          , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_1_reg[9])}), (chn_idata_data_sva_3_47_31_1[14:11]),
          (signext_4_1(~ IsNaN_5U_10U_land_3_lpi_1_dfm_5)), 4'b1110, (signext_4_1(IntSaturation_17U_8U_o_7_1_2_lpi_1_dfm_1[6])),
          reg_FpIntToFloat_17U_5U_10U_o_expo_2_lpi_1_dfm_8_1_itm, {cvt_or_2_cse ,
          cfg_mode_eql_1_sva_6 , (cvt_and_259_nl) , (cvt_and_260_nl) , (and_3148_nl)
          , or_5174_tmp});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_out_rsci_d_61_58 <= 4'b0;
    end
    else if ( ((~ (mux_2308_nl)) | (~ cvt_unequal_tmp_21) | cfg_mode_eql_1_sva_6)
        & or_5189_cse & and_dcpl_1742 ) begin
      chn_out_rsci_d_61_58 <= MUX1HOT_v_4_6_2((FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5[12:9]),
          (chn_idata_data_sva_3_111_95_1[14:11]), (signext_4_1(~ IsNaN_5U_10U_land_5_lpi_1_dfm_5)),
          4'b1110, (signext_4_1(IntSaturation_17U_8U_o_7_1_4_lpi_1_dfm_1[6])), reg_FpIntToFloat_17U_5U_10U_o_expo_4_lpi_1_dfm_9_1_itm,
          {(and_3140_nl) , cfg_mode_eql_1_sva_6 , (cvt_and_255_nl) , (cvt_and_256_nl)
          , cvt_asn_339 , or_5176_tmp});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_out_rsci_d_93_90 <= 4'b0;
    end
    else if ( ((~ (mux_2314_nl)) | (~ cvt_unequal_tmp_21) | cfg_mode_eql_1_sva_6)
        & or_5189_cse & and_dcpl_1742 ) begin
      chn_out_rsci_d_93_90 <= MUX1HOT_v_4_6_2(({(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_reg[2:0])
          , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_1_reg[9])}), (chn_idata_data_sva_3_175_159_1[14:11]),
          (signext_4_1(~ IsNaN_5U_10U_land_7_lpi_1_dfm_6)), 4'b1110, (signext_4_1(IntSaturation_17U_8U_o_7_1_6_lpi_1_dfm_1[6])),
          reg_FpIntToFloat_17U_5U_10U_o_expo_6_lpi_1_dfm_9_1_itm, {cvt_or_10_cse
          , cfg_mode_eql_1_sva_6 , (cvt_and_251_nl) , (cvt_and_252_nl) , (and_3136_nl)
          , or_5178_tmp});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_out_rsci_d_109_106 <= 4'b0;
    end
    else if ( ((~ (mux_2320_nl)) | (~ cvt_unequal_tmp_21) | cfg_mode_eql_1_sva_6)
        & or_5189_cse & and_dcpl_1742 ) begin
      chn_out_rsci_d_109_106 <= MUX1HOT_v_4_6_2(({(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_reg[2:0])
          , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_1_reg[9])}), (chn_idata_data_sva_3_207_191_1[14:11]),
          (signext_4_1(~ IsNaN_5U_10U_land_8_lpi_1_dfm_5)), 4'b1110, (signext_4_1(IntSaturation_17U_8U_o_7_1_7_lpi_1_dfm_1[6])),
          reg_FpIntToFloat_17U_5U_10U_o_expo_7_lpi_1_dfm_9_1_itm, {cvt_or_12_cse
          , cfg_mode_eql_1_sva_6 , (cvt_and_249_nl) , (cvt_and_250_nl) , (and_3133_nl)
          , or_5179_tmp});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_out_rsci_d_125_122 <= 4'b0;
    end
    else if ( ((~ (mux_2327_nl)) | (~ cvt_unequal_tmp_21) | cfg_mode_eql_1_sva_6)
        & or_5189_cse & and_dcpl_1742 ) begin
      chn_out_rsci_d_125_122 <= MUX1HOT_v_4_6_2(({(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_reg[2:0])
          , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_1_reg[9])}), (chn_idata_data_sva_3_239_223_1[14:11]),
          (signext_4_1(~ IsNaN_5U_10U_land_9_lpi_1_dfm_5)), 4'b1110, (signext_4_1(IntSaturation_17U_8U_o_7_1_8_lpi_1_dfm_1[6])),
          reg_FpIntToFloat_17U_5U_10U_o_expo_8_lpi_1_dfm_10_1_itm, {(and_3128_nl)
          , cfg_mode_eql_1_sva_6 , (cvt_and_247_nl) , (cvt_and_248_nl) , (and_3130_nl)
          , or_5180_tmp});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_out_rsci_d_157_154 <= 4'b0;
    end
    else if ( ((~ (mux_2332_nl)) | (~ cvt_unequal_tmp_21) | cfg_mode_eql_1_sva_6)
        & or_5189_cse & and_dcpl_1742 ) begin
      chn_out_rsci_d_157_154 <= MUX1HOT_v_4_6_2(({(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_reg[2:0])
          , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_1_reg[9])}), (chn_idata_data_sva_3_303_287_1[14:11]),
          (signext_4_1(~ IsNaN_5U_10U_land_1_lpi_1_dfm_3)), 4'b1110, (signext_4_1(IntSaturation_17U_8U_o_7_1_10_lpi_1_dfm_1[6])),
          reg_FpIntToFloat_17U_5U_10U_o_expo_10_lpi_1_dfm_9_1_itm, {cvt_or_18_cse
          , cfg_mode_eql_1_sva_6 , (cvt_and_243_nl) , (cvt_and_244_nl) , (and_3124_nl)
          , or_5182_tmp});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_out_rsci_d_173_170 <= 4'b0;
    end
    else if ( ((~ (mux_2338_nl)) | (~ cvt_unequal_tmp_21) | cfg_mode_eql_1_sva_6)
        & or_5189_cse & and_dcpl_1742 ) begin
      chn_out_rsci_d_173_170 <= MUX1HOT_v_4_6_2(({(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_reg[2:0])
          , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_1_reg[9])}), (chn_idata_data_sva_3_335_319_1[14:11]),
          (signext_4_1(~ IsNaN_5U_10U_land_10_lpi_1_dfm_5)), 4'b1110, (signext_4_1(IntSaturation_17U_8U_o_7_1_11_lpi_1_dfm_1[6])),
          reg_FpIntToFloat_17U_5U_10U_o_expo_11_lpi_1_dfm_9_1_itm, {cvt_or_20_cse
          , cfg_mode_eql_1_sva_6 , (cvt_and_241_nl) , (cvt_and_242_nl) , (and_3121_nl)
          , or_5183_tmp});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_out_rsci_d_189_186 <= 4'b0;
    end
    else if ( ((~ (mux_2344_nl)) | (~ cvt_unequal_tmp_21) | cfg_mode_eql_1_sva_6)
        & or_5189_cse & and_dcpl_1742 ) begin
      chn_out_rsci_d_189_186 <= MUX1HOT_v_4_6_2(({(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_reg[2:0])
          , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_1_reg[9])}), (chn_idata_data_sva_3_367_351_1[14:11]),
          (signext_4_1(~ IsNaN_5U_10U_land_11_lpi_1_dfm_5)), 4'b1110, (signext_4_1(IntSaturation_17U_8U_o_7_1_12_lpi_1_dfm_1[6])),
          reg_FpIntToFloat_17U_5U_10U_o_expo_12_lpi_1_dfm_10_1_itm, {(and_3116_nl)
          , cfg_mode_eql_1_sva_6 , (cvt_and_239_nl) , (cvt_and_240_nl) , (and_3118_nl)
          , or_5184_tmp});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_out_rsci_d_205_202 <= 4'b0;
    end
    else if ( ((~ (mux_2349_nl)) | (~ cvt_unequal_tmp_21) | cfg_mode_eql_1_sva_6)
        & or_5189_cse & and_dcpl_1742 ) begin
      chn_out_rsci_d_205_202 <= MUX1HOT_v_4_6_2(({(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_reg[2:0])
          , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_1_reg[9])}), (chn_idata_data_sva_3_399_383_1[14:11]),
          (signext_4_1(~ IsNaN_5U_10U_land_12_lpi_1_dfm_5)), 4'b1110, (signext_4_1(IntSaturation_17U_8U_o_7_1_13_lpi_1_dfm_1[6])),
          reg_FpIntToFloat_17U_5U_10U_o_expo_13_lpi_1_dfm_9_1_itm, {cvt_or_24_cse
          , cfg_mode_eql_1_sva_6 , (cvt_and_237_nl) , (cvt_and_238_nl) , (and_3115_nl)
          , or_5185_tmp});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_out_rsci_d_221_218 <= 4'b0;
      chn_out_rsci_d_253_250 <= 4'b0;
    end
    else if ( and_3063_cse ) begin
      chn_out_rsci_d_221_218 <= MUX1HOT_v_4_6_2(({(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_reg[2:0])
          , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_1_reg[9])}), (chn_idata_data_sva_3_431_415_1[14:11]),
          (signext_4_1(~ IsNaN_5U_10U_land_13_lpi_1_dfm_5)), 4'b1110, (signext_4_1(IntSaturation_17U_8U_o_7_1_14_lpi_1_dfm_1[6])),
          reg_FpIntToFloat_17U_5U_10U_o_expo_14_lpi_1_dfm_10_1_itm, {(and_3110_nl)
          , cfg_mode_eql_1_sva_6 , (cvt_and_235_nl) , (cvt_and_236_nl) , (and_3112_nl)
          , or_5186_tmp});
      chn_out_rsci_d_253_250 <= MUX1HOT_v_4_6_2(({(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_reg[2:0])
          , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_1_reg[9])}), (signext_4_1(~
          IsNaN_5U_10U_land_15_lpi_1_dfm_3)), 4'b1110, (signext_4_1(IntSaturation_17U_8U_o_7_1_lpi_1_dfm_1[6])),
          (chn_idata_data_sva_3_495_479_1[14:11]), reg_FpIntToFloat_17U_5U_10U_o_expo_lpi_1_dfm_11_1_itm,
          {(and_3104_nl) , (cvt_and_231_nl) , (cvt_and_232_nl) , (and_3105_nl) ,
          cfg_mode_eql_1_sva_6 , or_5188_tmp});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_out_rsci_d_237_234 <= 4'b0;
    end
    else if ( ((mux_2362_nl) | (~ cvt_unequal_tmp_21) | cfg_mode_eql_1_sva_6) & or_5189_cse
        & and_dcpl_1742 ) begin
      chn_out_rsci_d_237_234 <= MUX1HOT_v_4_6_2(({(reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_reg[2:0])
          , (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_1_reg[9])}), (chn_idata_data_sva_3_463_447_1[14:11]),
          (signext_4_1(~ IsNaN_5U_10U_land_14_lpi_1_dfm_6)), 4'b1110, (signext_4_1(IntSaturation_17U_8U_o_7_1_15_lpi_1_dfm_1[6])),
          reg_FpIntToFloat_17U_5U_10U_o_expo_15_lpi_1_dfm_10_1_itm, {cvt_or_28_cse
          , cfg_mode_eql_1_sva_6 , (cvt_and_233_nl) , (cvt_and_234_nl) , (and_3109_nl)
          , or_5187_tmp});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_out_rsci_d_0 <= 1'b0;
      chn_out_rsci_d_15 <= 1'b0;
      chn_out_rsci_d_16 <= 1'b0;
      chn_out_rsci_d_31 <= 1'b0;
      chn_out_rsci_d_32 <= 1'b0;
      chn_out_rsci_d_47 <= 1'b0;
      chn_out_rsci_d_48 <= 1'b0;
      chn_out_rsci_d_63 <= 1'b0;
      chn_out_rsci_d_64 <= 1'b0;
      chn_out_rsci_d_79 <= 1'b0;
      chn_out_rsci_d_80 <= 1'b0;
      chn_out_rsci_d_95 <= 1'b0;
      chn_out_rsci_d_96 <= 1'b0;
      chn_out_rsci_d_111 <= 1'b0;
      chn_out_rsci_d_112 <= 1'b0;
      chn_out_rsci_d_127 <= 1'b0;
      chn_out_rsci_d_128 <= 1'b0;
      chn_out_rsci_d_143 <= 1'b0;
      chn_out_rsci_d_144 <= 1'b0;
      chn_out_rsci_d_159 <= 1'b0;
      chn_out_rsci_d_160 <= 1'b0;
      chn_out_rsci_d_175 <= 1'b0;
      chn_out_rsci_d_176 <= 1'b0;
      chn_out_rsci_d_191 <= 1'b0;
      chn_out_rsci_d_192 <= 1'b0;
      chn_out_rsci_d_207 <= 1'b0;
      chn_out_rsci_d_208 <= 1'b0;
      chn_out_rsci_d_223 <= 1'b0;
      chn_out_rsci_d_224 <= 1'b0;
      chn_out_rsci_d_239 <= 1'b0;
    end
    else if ( chn_out_and_32_cse ) begin
      chn_out_rsci_d_0 <= MUX_s_1_2_2((cvt_mux_2280_nl), (cvt_mux_2281_nl), and_dcpl_98);
      chn_out_rsci_d_15 <= MUX_s_1_2_2((cvt_mux_2373_nl), reg_chn_idata_data_sva_3_15_0_reg,
          cfg_mode_eql_1_sva_6);
      chn_out_rsci_d_16 <= MUX_s_1_2_2((cvt_mux_2284_nl), (cvt_mux_2285_nl), and_dcpl_98);
      chn_out_rsci_d_31 <= MUX_s_1_2_2((cvt_mux_2346_nl), (chn_idata_data_sva_3_47_31_1[16]),
          cfg_mode_eql_1_sva_6);
      chn_out_rsci_d_32 <= MUX_s_1_2_2((cvt_mux_2288_nl), (cvt_mux_2289_nl), and_dcpl_98);
      chn_out_rsci_d_47 <= MUX_s_1_2_2((cvt_mux_2348_nl), (chn_idata_data_sva_3_79_63_1[16]),
          cfg_mode_eql_1_sva_6);
      chn_out_rsci_d_48 <= MUX_s_1_2_2((cvt_mux_2292_nl), (cvt_mux_2293_nl), and_dcpl_98);
      chn_out_rsci_d_63 <= MUX_s_1_2_2((cvt_mux_2350_nl), (chn_idata_data_sva_3_111_95_1[16]),
          cfg_mode_eql_1_sva_6);
      chn_out_rsci_d_64 <= MUX_s_1_2_2((cvt_mux_2296_nl), (cvt_mux_2297_nl), and_dcpl_98);
      chn_out_rsci_d_79 <= MUX_s_1_2_2((cvt_mux_2352_nl), (chn_idata_data_sva_3_143_127_1[16]),
          cfg_mode_eql_1_sva_6);
      chn_out_rsci_d_80 <= MUX_s_1_2_2((cvt_mux_2300_nl), (cvt_mux_2301_nl), and_dcpl_98);
      chn_out_rsci_d_95 <= MUX_s_1_2_2((cvt_mux_2354_nl), (chn_idata_data_sva_3_175_159_1[16]),
          cfg_mode_eql_1_sva_6);
      chn_out_rsci_d_96 <= MUX_s_1_2_2((cvt_mux_2304_nl), (cvt_mux_2305_nl), and_dcpl_98);
      chn_out_rsci_d_111 <= MUX_s_1_2_2((cvt_mux_2358_nl), (chn_idata_data_sva_3_207_191_1[16]),
          cfg_mode_eql_1_sva_6);
      chn_out_rsci_d_112 <= MUX_s_1_2_2((cvt_mux_2308_nl), (cvt_mux_2309_nl), and_dcpl_98);
      chn_out_rsci_d_127 <= MUX_s_1_2_2((cvt_mux_2360_nl), (chn_idata_data_sva_3_239_223_1[16]),
          cfg_mode_eql_1_sva_6);
      chn_out_rsci_d_128 <= MUX_s_1_2_2((cvt_mux_2312_nl), (cvt_mux_2313_nl), and_dcpl_98);
      chn_out_rsci_d_143 <= MUX_s_1_2_2((cvt_mux_2362_nl), (chn_idata_data_sva_3_271_255_1[16]),
          cfg_mode_eql_1_sva_6);
      chn_out_rsci_d_144 <= MUX_s_1_2_2((cvt_mux_2316_nl), (cvt_mux_2317_nl), and_dcpl_98);
      chn_out_rsci_d_159 <= MUX_s_1_2_2((cvt_mux_2364_nl), (chn_idata_data_sva_3_303_287_1[16]),
          cfg_mode_eql_1_sva_6);
      chn_out_rsci_d_160 <= MUX_s_1_2_2((cvt_mux_2320_nl), (cvt_mux_2321_nl), and_dcpl_98);
      chn_out_rsci_d_175 <= MUX_s_1_2_2((cvt_mux_2366_nl), (chn_idata_data_sva_3_335_319_1[16]),
          cfg_mode_eql_1_sva_6);
      chn_out_rsci_d_176 <= MUX_s_1_2_2((cvt_mux_2324_nl), (cvt_mux_2325_nl), and_dcpl_98);
      chn_out_rsci_d_191 <= MUX_s_1_2_2((cvt_mux_2370_nl), (chn_idata_data_sva_3_367_351_1[16]),
          cfg_mode_eql_1_sva_6);
      chn_out_rsci_d_192 <= MUX_s_1_2_2((cvt_mux_2328_nl), (cvt_mux_2329_nl), and_dcpl_98);
      chn_out_rsci_d_207 <= MUX_s_1_2_2((cvt_mux_2372_nl), (chn_idata_data_sva_3_399_383_1[16]),
          cfg_mode_eql_1_sva_6);
      chn_out_rsci_d_208 <= MUX_s_1_2_2((cvt_mux_2332_nl), (cvt_mux_2333_nl), and_dcpl_98);
      chn_out_rsci_d_223 <= MUX_s_1_2_2((cvt_mux_2368_nl), (chn_idata_data_sva_3_431_415_1[16]),
          cfg_mode_eql_1_sva_6);
      chn_out_rsci_d_224 <= MUX_s_1_2_2((cvt_mux_2336_nl), (cvt_mux_2337_nl), and_dcpl_98);
      chn_out_rsci_d_239 <= MUX_s_1_2_2((cvt_mux_2356_nl), (chn_idata_data_sva_3_463_447_1[16]),
          cfg_mode_eql_1_sva_6);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_out_rsci_d_240 <= 1'b0;
      chn_out_rsci_d_255 <= 1'b0;
    end
    else if ( chn_out_and_77_cse ) begin
      chn_out_rsci_d_240 <= MUX_s_1_2_2((chn_idata_data_sva_3_495_479_1[1]), (cvt_mux_2340_nl),
          and_dcpl_102);
      chn_out_rsci_d_255 <= MUX_s_1_2_2((chn_idata_data_sva_3_495_479_1[16]), (cvt_mux_2341_nl),
          and_dcpl_102);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_out_rsci_ld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_103 | and_dcpl_105) ) begin
      reg_chn_out_rsci_ld_core_psct_cse <= ~ and_dcpl_105;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_1 <= 1'b0;
    end
    else if ( core_wen & (or_tmp_3487 | main_stage_v_1_mx0c1) ) begin
      main_stage_v_1 <= ~ main_stage_v_1_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_2_sva_2 <= 3'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_nl) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_2_sva_2 <= FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_2_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_idata_data_sva_1_27_0_1 <= 28'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_5_nl) ) begin
      chn_idata_data_sva_1_27_0_1 <= chn_in_rsci_d_mxwt[27:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_8_nl)) ) begin
      cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_2
          <= cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_10_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_st_2
          <= cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_3_sva_2 <= 3'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_11_nl) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_3_sva_2 <= FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_3_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_idata_data_sva_1_59_31_1 <= 29'b0;
      chn_idata_data_sva_1_91_63_1 <= 29'b0;
      chn_idata_data_sva_1_123_95_1 <= 29'b0;
      chn_idata_data_sva_1_155_127_1 <= 29'b0;
      chn_idata_data_sva_1_187_159_1 <= 29'b0;
      chn_idata_data_sva_1_219_191_1 <= 29'b0;
      chn_idata_data_sva_1_251_223_1 <= 29'b0;
      chn_idata_data_sva_1_283_255_1 <= 29'b0;
      chn_idata_data_sva_1_315_287_1 <= 29'b0;
      chn_idata_data_sva_1_347_319_1 <= 29'b0;
      chn_idata_data_sva_1_379_351_1 <= 29'b0;
      chn_idata_data_sva_1_411_383_1 <= 29'b0;
      chn_idata_data_sva_1_443_415_1 <= 29'b0;
      chn_idata_data_sva_1_475_447_1 <= 29'b0;
      chn_idata_data_sva_1_507_479_1 <= 29'b0;
      cfg_truncate_1_sva_2 <= 6'b0;
      cfg_proc_precision_1_sva_st_64 <= 2'b0;
      cfg_mode_eql_1_sva_4 <= 1'b0;
      cvt_unequal_tmp_19 <= 1'b0;
    end
    else if ( chn_idata_data_and_1_cse ) begin
      chn_idata_data_sva_1_59_31_1 <= chn_in_rsci_d_mxwt[59:31];
      chn_idata_data_sva_1_91_63_1 <= chn_in_rsci_d_mxwt[91:63];
      chn_idata_data_sva_1_123_95_1 <= chn_in_rsci_d_mxwt[123:95];
      chn_idata_data_sva_1_155_127_1 <= chn_in_rsci_d_mxwt[155:127];
      chn_idata_data_sva_1_187_159_1 <= chn_in_rsci_d_mxwt[187:159];
      chn_idata_data_sva_1_219_191_1 <= chn_in_rsci_d_mxwt[219:191];
      chn_idata_data_sva_1_251_223_1 <= chn_in_rsci_d_mxwt[251:223];
      chn_idata_data_sva_1_283_255_1 <= chn_in_rsci_d_mxwt[283:255];
      chn_idata_data_sva_1_315_287_1 <= chn_in_rsci_d_mxwt[315:287];
      chn_idata_data_sva_1_347_319_1 <= chn_in_rsci_d_mxwt[347:319];
      chn_idata_data_sva_1_379_351_1 <= chn_in_rsci_d_mxwt[379:351];
      chn_idata_data_sva_1_411_383_1 <= chn_in_rsci_d_mxwt[411:383];
      chn_idata_data_sva_1_443_415_1 <= chn_in_rsci_d_mxwt[443:415];
      chn_idata_data_sva_1_475_447_1 <= chn_in_rsci_d_mxwt[475:447];
      chn_idata_data_sva_1_507_479_1 <= chn_in_rsci_d_mxwt[507:479];
      cfg_truncate_1_sva_2 <= cfg_truncate_rsci_d;
      cfg_proc_precision_1_sva_st_64 <= cfg_proc_precision_rsci_d;
      cfg_mode_eql_1_sva_4 <= cfg_mode_eql_rsci_d;
      cvt_unequal_tmp_19 <= cvt_cvt_nand_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_14_nl)) ) begin
      cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2
          <= cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_16_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_st_2
          <= cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_4_sva_2 <= 3'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_17_nl) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_4_sva_2 <= FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_4_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_19_nl)) ) begin
      cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2
          <= cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_21_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_st_2
          <= cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_5_sva_2 <= 3'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_22_nl) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_5_sva_2 <= FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_5_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_24_nl)) ) begin
      cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2
          <= cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_26_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_st_2
          <= cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_6_sva_2 <= 3'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_28_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_6_sva_2 <= FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_6_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_30_nl)) ) begin
      cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2
          <= cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_32_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_st_2
          <= cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_7_sva_2 <= 3'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_34_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_7_sva_2 <= FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_7_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_36_nl)) ) begin
      cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2
          <= cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_38_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_st_2
          <= cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_8_sva_2 <= 3'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_41_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_8_sva_2 <= FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_8_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_42_nl)) ) begin
      cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2
          <= cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_44_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_st_2
          <= cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_9_sva_2 <= 3'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_45_nl) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_9_sva_2 <= FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_9_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_47_nl)) ) begin
      cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2
          <= cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_49_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_st_2
          <= cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_10_sva_2 <= 3'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_50_nl) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_10_sva_2 <= FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_10_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_52_nl)) ) begin
      cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2
          <= cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_54_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_st_2
          <= cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_11_sva_2 <= 3'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_56_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_11_sva_2 <= FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_11_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_58_nl)) ) begin
      cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2
          <= cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_60_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_st_2
          <= cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_12_sva_2 <= 3'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_61_nl) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_12_sva_2 <= FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_12_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_63_nl)) ) begin
      cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2
          <= cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_65_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_st_2
          <= cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_13_sva_2 <= 3'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_66_nl) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_13_sva_2 <= FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_13_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_68_nl)) ) begin
      cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2
          <= cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_70_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_st_2
          <= cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_14_sva_2 <= 3'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_72_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_14_sva_2 <= FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_14_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_74_nl)) ) begin
      cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2
          <= cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_76_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_st_2
          <= cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_15_sva_2 <= 3'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_77_nl) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_15_sva_2 <= FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_15_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_79_nl)) ) begin
      cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2
          <= cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_81_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_st_2
          <= cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_16_sva_2 <= 3'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_82_nl) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_16_sva_2 <= FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_16_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_84_nl)) ) begin
      cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2
          <= cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_86_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_st_2
          <= cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_2 <= 3'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_87_nl) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_2 <= FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_89_nl)) ) begin
      cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_st_2
          <= cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_itm_8_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_91_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_2
          <= cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_itm_7_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_4_svs_st_2
          <= 1'b0;
      cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2
          <= 1'b0;
      cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2
          <= 1'b0;
      cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
          <= 1'b0;
      cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2
          <= 1'b0;
      cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
          <= 1'b0;
      cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
          <= 1'b0;
      cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2
          <= 1'b0;
      cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2
          <= 1'b0;
      cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
          <= 1'b0;
      cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
          <= 1'b0;
      cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2
          <= 1'b0;
      cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
          <= 1'b0;
      cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2
          <= 1'b0;
      cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2
          <= 1'b0;
      cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_2
          <= 1'b0;
      cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_2
          <= 1'b0;
      IsNaN_8U_23U_land_lpi_1_dfm_3 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_2
          <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_15_itm_2 <= 1'b0;
      cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2
          <= 1'b0;
      IsNaN_8U_23U_land_15_lpi_1_dfm_3 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_2
          <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_14_itm_2 <= 1'b0;
      cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2
          <= 1'b0;
      IsNaN_8U_23U_land_14_lpi_1_dfm_3 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_2
          <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_13_itm_2 <= 1'b0;
      cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2
          <= 1'b0;
      IsNaN_8U_23U_land_13_lpi_1_dfm_3 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_2
          <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_12_itm_2 <= 1'b0;
      cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2
          <= 1'b0;
      IsNaN_8U_23U_land_12_lpi_1_dfm_3 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_2
          <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_11_itm_2 <= 1'b0;
      cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2
          <= 1'b0;
      IsNaN_8U_23U_land_11_lpi_1_dfm_3 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_2
          <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_10_itm_2 <= 1'b0;
      cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2
          <= 1'b0;
      IsNaN_8U_23U_land_10_lpi_1_dfm_3 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_2
          <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_9_itm_2 <= 1'b0;
      cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2
          <= 1'b0;
      IsNaN_8U_23U_land_9_lpi_1_dfm_3 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_2
          <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_8_itm_2 <= 1'b0;
      cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2
          <= 1'b0;
      IsNaN_8U_23U_land_8_lpi_1_dfm_3 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_2
          <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_7_itm_2 <= 1'b0;
      cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2
          <= 1'b0;
      IsNaN_8U_23U_land_7_lpi_1_dfm_3 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_2
          <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_6_itm_2 <= 1'b0;
      cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2
          <= 1'b0;
      IsNaN_8U_23U_land_6_lpi_1_dfm_3 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_2
          <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_5_itm_2 <= 1'b0;
      cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2
          <= 1'b0;
      IsNaN_8U_23U_nor_4_itm_2 <= 1'b0;
      IsNaN_8U_23U_IsNaN_8U_23U_nand_4_itm_2 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_2
          <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_4_itm_2 <= 1'b0;
      cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2
          <= 1'b0;
      IsNaN_8U_23U_land_4_lpi_1_dfm_3 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_2
          <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_3_itm_2 <= 1'b0;
      cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2
          <= 1'b0;
      IsNaN_8U_23U_land_3_lpi_1_dfm_3 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_2
          <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_2_itm_2 <= 1'b0;
      cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2
          <= 1'b0;
      IsNaN_8U_23U_land_2_lpi_1_dfm_3 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_2
          <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_1_itm_2 <= 1'b0;
      cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_2
          <= 1'b0;
      IsNaN_8U_23U_land_1_lpi_1_dfm_3 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_2
          <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_itm_2 <= 1'b0;
    end
    else if ( FpWidthDec_8U_23U_5U_10U_1U_1U_if_and_cse ) begin
      cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_4_svs_st_2
          <= cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_itm_8_1;
      cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2
          <= cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1;
      cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2
          <= cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1;
      cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
          <= cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1;
      cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2
          <= cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1;
      cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
          <= cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1;
      cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
          <= cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1;
      cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2
          <= cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1;
      cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2
          <= cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1;
      cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
          <= cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1;
      cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
          <= cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1;
      cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2
          <= cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1;
      cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
          <= cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1;
      cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2
          <= cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1;
      cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2
          <= cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1;
      cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_2
          <= cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_itm_8_1;
      cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_2
          <= cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_itm_8_1;
      IsNaN_8U_23U_land_lpi_1_dfm_3 <= IsNaN_8U_23U_IsNaN_8U_23U_nor_15_tmp;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_2
          <= cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_itm_7_1;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_15_itm_2 <= ~((cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_4_tmp==5'b11111)
          & (FpMantRNE_24U_11U_else_mux_31_nl) & cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_itm_8_1
          & (~ cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_itm_7_1));
      cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2
          <= cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1;
      IsNaN_8U_23U_land_15_lpi_1_dfm_3 <= IsNaN_8U_23U_IsNaN_8U_23U_nor_14_tmp;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_2
          <= cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_14_itm_2 <= ~((cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp==5'b11111)
          & (FpMantRNE_24U_11U_else_mux_29_nl) & cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1
          & (~ cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1));
      cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2
          <= cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1;
      IsNaN_8U_23U_land_14_lpi_1_dfm_3 <= IsNaN_8U_23U_IsNaN_8U_23U_nor_13_tmp;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_2
          <= cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_13_itm_2 <= ~((cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp==5'b11111)
          & (FpMantRNE_24U_11U_else_mux_27_nl) & cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1
          & (~ cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1));
      cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2
          <= cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1;
      IsNaN_8U_23U_land_13_lpi_1_dfm_3 <= IsNaN_8U_23U_IsNaN_8U_23U_nor_12_tmp;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_2
          <= cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_12_itm_2 <= ~((cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp==5'b11111)
          & (FpMantRNE_24U_11U_else_mux_25_nl) & cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1
          & (~ cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1));
      cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2
          <= cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1;
      IsNaN_8U_23U_land_12_lpi_1_dfm_3 <= IsNaN_8U_23U_IsNaN_8U_23U_nor_11_tmp;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_2
          <= cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_11_itm_2 <= ~((cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp==5'b11111)
          & (FpMantRNE_24U_11U_else_mux_23_nl) & cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1
          & (~ cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1));
      cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2
          <= cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1;
      IsNaN_8U_23U_land_11_lpi_1_dfm_3 <= IsNaN_8U_23U_IsNaN_8U_23U_nor_10_tmp;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_2
          <= cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_10_itm_2 <= ~((cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp==5'b11111)
          & (FpMantRNE_24U_11U_else_mux_21_nl) & cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1
          & (~ cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1));
      cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2
          <= cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1;
      IsNaN_8U_23U_land_10_lpi_1_dfm_3 <= IsNaN_8U_23U_IsNaN_8U_23U_nor_9_tmp;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_2
          <= cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_9_itm_2 <= ~((cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp==5'b11111)
          & (FpMantRNE_24U_11U_else_mux_19_nl) & cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1
          & (~ cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1));
      cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2
          <= cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1;
      IsNaN_8U_23U_land_9_lpi_1_dfm_3 <= IsNaN_8U_23U_IsNaN_8U_23U_nor_8_tmp;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_2
          <= cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_8_itm_2 <= ~((cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp==5'b11111)
          & (FpMantRNE_24U_11U_else_mux_17_nl) & cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1
          & (~ cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1));
      cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2
          <= cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1;
      IsNaN_8U_23U_land_8_lpi_1_dfm_3 <= IsNaN_8U_23U_IsNaN_8U_23U_nor_7_tmp;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_2
          <= cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_7_itm_2 <= ~((cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp==5'b11111)
          & (FpMantRNE_24U_11U_else_mux_15_nl) & cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1
          & (~ cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1));
      cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2
          <= cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1;
      IsNaN_8U_23U_land_7_lpi_1_dfm_3 <= IsNaN_8U_23U_IsNaN_8U_23U_nor_6_tmp;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_2
          <= cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_6_itm_2 <= ~((cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp==5'b11111)
          & (FpMantRNE_24U_11U_else_mux_13_nl) & cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1
          & (~ cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1));
      cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2
          <= cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1;
      IsNaN_8U_23U_land_6_lpi_1_dfm_3 <= IsNaN_8U_23U_IsNaN_8U_23U_nor_5_tmp;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_2
          <= cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_5_itm_2 <= ~((cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp==5'b11111)
          & (FpMantRNE_24U_11U_else_mux_11_nl) & cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1
          & (~ cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1));
      cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2
          <= cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1;
      IsNaN_8U_23U_nor_4_itm_2 <= IsNaN_8U_23U_nor_4_tmp;
      IsNaN_8U_23U_IsNaN_8U_23U_nand_4_itm_2 <= IsNaN_8U_23U_IsNaN_8U_23U_nand_4_tmp;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_2
          <= cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_4_itm_2 <= ~((cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp==5'b11111)
          & (FpMantRNE_24U_11U_else_mux_9_nl) & cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1
          & (~ cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1));
      cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2
          <= cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1;
      IsNaN_8U_23U_land_4_lpi_1_dfm_3 <= IsNaN_8U_23U_IsNaN_8U_23U_nor_3_tmp;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_2
          <= cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_3_itm_2 <= ~((cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp==5'b11111)
          & (FpMantRNE_24U_11U_else_mux_7_nl) & cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1
          & (~ cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1));
      cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2
          <= cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1;
      IsNaN_8U_23U_land_3_lpi_1_dfm_3 <= IsNaN_8U_23U_IsNaN_8U_23U_nor_2_tmp;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_2
          <= cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_2_itm_2 <= ~((cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp==5'b11111)
          & (FpMantRNE_24U_11U_else_mux_5_nl) & cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1
          & (~ cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1));
      cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2
          <= cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1;
      IsNaN_8U_23U_land_2_lpi_1_dfm_3 <= IsNaN_8U_23U_IsNaN_8U_23U_nor_1_tmp;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_2
          <= cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_1_itm_2 <= ~((cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp==5'b11111)
          & (FpMantRNE_24U_11U_else_mux_3_nl) & cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1
          & (~ cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1));
      cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_2
          <= cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_itm_8_1;
      IsNaN_8U_23U_land_1_lpi_1_dfm_3 <= IsNaN_8U_23U_IsNaN_8U_23U_nor_tmp;
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_2
          <= cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1;
      FpWidthDec_8U_23U_5U_10U_1U_1U_nand_itm_2 <= ~((cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_tmp==5'b11111)
          & (FpMantRNE_24U_11U_else_mux_1_nl) & cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_itm_8_1
          & (~ cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntMulExt_33U_16U_49U_return_2_sva_2 <= 49'b0;
      IntMulExt_33U_16U_49U_return_3_sva_2 <= 49'b0;
      IntMulExt_33U_16U_49U_return_9_sva_2 <= 49'b0;
    end
    else if ( IntMulExt_33U_16U_49U_and_11_cse ) begin
      IntMulExt_33U_16U_49U_return_2_sva_2 <= conv_s2u_49_49($signed((cvt_2_IntSubExt_32U_32U_33U_o_acc_1_nl))
          * $signed((cfg_scale_rsci_d)));
      IntMulExt_33U_16U_49U_return_3_sva_2 <= conv_s2u_49_49($signed((cvt_3_IntSubExt_32U_32U_33U_o_acc_1_nl))
          * $signed((cfg_scale_rsci_d)));
      IntMulExt_33U_16U_49U_return_9_sva_2 <= conv_s2u_49_49($signed((cvt_9_IntSubExt_32U_32U_33U_o_acc_1_nl))
          * $signed((cfg_scale_rsci_d)));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntMulExt_33U_16U_49U_return_4_sva_1 <= 49'b0;
    end
    else if ( core_wen & (and_550_cse | (and_2186_cse & and_dcpl_73) | IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1)
        ) begin
      IntMulExt_33U_16U_49U_return_4_sva_1 <= MUX_v_49_2_2((cvt_4_IntMulExt_33U_16U_49U_o_mul_2_nl),
          IntShiftRightSat_49U_6U_17U_i_4_sva_mx0w1, IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntMulExt_33U_16U_49U_return_6_sva_1 <= 49'b0;
      IntMulExt_33U_16U_49U_return_8_sva_1 <= 49'b0;
      IntMulExt_33U_16U_49U_return_7_sva_1 <= 49'b0;
      IntMulExt_33U_16U_49U_return_10_sva_1 <= 49'b0;
      IntMulExt_33U_16U_49U_return_12_sva_1 <= 49'b0;
      IntMulExt_33U_16U_49U_return_11_sva_1 <= 49'b0;
      IntMulExt_33U_16U_49U_return_14_sva_1 <= 49'b0;
      IntMulExt_33U_16U_49U_return_sva_1 <= 49'b0;
      IntMulExt_33U_16U_49U_return_15_sva_1 <= 49'b0;
      IntMulExt_33U_16U_49U_return_13_sva_1 <= 49'b0;
    end
    else if ( IntMulExt_33U_16U_49U_and_1_cse ) begin
      IntMulExt_33U_16U_49U_return_6_sva_1 <= MUX_v_49_2_2((cvt_6_IntMulExt_33U_16U_49U_o_mul_2_nl),
          IntShiftRightSat_49U_6U_17U_i_6_sva_mx0w1, IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1);
      IntMulExt_33U_16U_49U_return_8_sva_1 <= MUX_v_49_2_2((cvt_8_IntMulExt_33U_16U_49U_o_mul_3_nl),
          IntShiftRightSat_49U_6U_17U_i_8_sva_mx0w1, IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1);
      IntMulExt_33U_16U_49U_return_7_sva_1 <= MUX_v_49_2_2((cvt_7_IntMulExt_33U_16U_49U_o_mul_2_nl),
          IntShiftRightSat_49U_6U_17U_i_7_sva_mx0w1, IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1);
      IntMulExt_33U_16U_49U_return_10_sva_1 <= MUX_v_49_2_2((cvt_10_IntMulExt_33U_16U_49U_o_mul_2_nl),
          IntShiftRightSat_49U_6U_17U_i_10_sva_mx0w1, IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1);
      IntMulExt_33U_16U_49U_return_12_sva_1 <= MUX_v_49_2_2((cvt_12_IntMulExt_33U_16U_49U_o_mul_3_nl),
          IntShiftRightSat_49U_6U_17U_i_12_sva_mx0w1, IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1);
      IntMulExt_33U_16U_49U_return_11_sva_1 <= MUX_v_49_2_2((cvt_11_IntMulExt_33U_16U_49U_o_mul_2_nl),
          IntShiftRightSat_49U_6U_17U_i_11_sva_mx0w1, IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1);
      IntMulExt_33U_16U_49U_return_14_sva_1 <= MUX_v_49_2_2((cvt_14_IntMulExt_33U_16U_49U_o_mul_3_nl),
          IntShiftRightSat_49U_6U_17U_i_14_sva_mx0w1, IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1);
      IntMulExt_33U_16U_49U_return_sva_1 <= MUX_v_49_2_2((cvt_16_IntMulExt_33U_16U_49U_o_mul_4_nl),
          IntShiftRightSat_49U_6U_17U_i_sva_mx0w1, IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1);
      IntMulExt_33U_16U_49U_return_15_sva_1 <= MUX_v_49_2_2((cvt_15_IntMulExt_33U_16U_49U_o_mul_3_nl),
          IntShiftRightSat_49U_6U_17U_i_15_sva_mx0w1, IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1);
      IntMulExt_33U_16U_49U_return_13_sva_1 <= MUX_v_49_2_2((cvt_13_IntMulExt_33U_16U_49U_o_mul_2_nl),
          IntShiftRightSat_49U_6U_17U_i_13_sva_mx0w1, IntMulExt_33U_16U_49U_return_4_sva_1_mx0c1);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntMulExt_33U_16U_49U_return_5_sva_2 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & mux_tmp_122 ) begin
      IntMulExt_33U_16U_49U_return_5_sva_2 <= conv_s2u_49_49($signed((cvt_5_IntSubExt_32U_32U_33U_o_acc_1_nl))
          * $signed((cfg_scale_rsci_d)));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_out_precision_1_sva_st_154 <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_159_nl) ) begin
      cfg_out_precision_1_sva_st_154 <= cfg_out_precision_rsci_d;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_cfg_proc_precision_1_sva_st_40_cse <= 2'b0;
      IntMulExt_33U_16U_49U_return_1_sva_2 <= 49'b0;
    end
    else if ( cfg_proc_precision_and_11_cse ) begin
      reg_cfg_proc_precision_1_sva_st_40_cse <= cfg_proc_precision_rsci_d;
      IntMulExt_33U_16U_49U_return_1_sva_2 <= conv_s2u_49_49($signed((cvt_1_IntSubExt_32U_32U_33U_o_acc_nl))
          * $signed((cfg_scale_rsci_d)));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_2 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_114 | main_stage_v_2_mx0c1) ) begin
      main_stage_v_2 <= ~ main_stage_v_2_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_idata_data_sva_2_47_31_1 <= 17'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_9_3_0_1 <= 4'b0;
      chn_idata_data_sva_2_79_63_1 <= 17'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_9_3_0_1 <= 4'b0;
      chn_idata_data_sva_2_111_95_1 <= 17'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_9_3_0_1 <= 4'b0;
      chn_idata_data_sva_2_143_127_1 <= 17'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_9_3_0_1 <= 4'b0;
      chn_idata_data_sva_2_175_159_1 <= 17'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_9_3_0_1 <= 4'b0;
      chn_idata_data_sva_2_207_191_1 <= 17'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_9_3_0_1 <= 4'b0;
      chn_idata_data_sva_2_239_223_1 <= 17'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_9_3_0_1 <= 4'b0;
      chn_idata_data_sva_2_271_255_1 <= 17'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_9_3_0_1 <= 4'b0;
      chn_idata_data_sva_2_303_287_1 <= 17'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_9_3_0_1 <= 4'b0;
      chn_idata_data_sva_2_335_319_1 <= 17'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_9_3_0_1 <= 4'b0;
      chn_idata_data_sva_2_367_351_1 <= 17'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_9_3_0_1 <= 4'b0;
      chn_idata_data_sva_2_399_383_1 <= 17'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_9_3_0_1 <= 4'b0;
      chn_idata_data_sva_2_431_415_1 <= 17'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_9_3_0_1 <= 4'b0;
      chn_idata_data_sva_2_463_447_1 <= 17'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_9_3_0_1 <= 4'b0;
      chn_idata_data_sva_2_495_479_1 <= 17'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_9_3_0_1 <= 4'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_9_3_0_1 <= 4'b0;
      cfg_out_precision_1_sva_st_113 <= 2'b0;
      IntShiftRightSat_49U_6U_17U_o_16_1_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_1_sva_2 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_2_sva_2 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_16_3_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_3_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_4_sva_2 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_16_5_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_5_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_6_sva_2 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_7_sva_2 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_8_sva_2 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_16_9_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_9_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_10_sva_2 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_11_sva_2 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_12_sva_2 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_13_sva_2 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_14_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_15_sva_2 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_sva_2 <= 1'b0;
      cfg_proc_precision_1_sva_st_65 <= 2'b0;
      IsNaN_5U_10U_land_3_lpi_1_dfm_4 <= 1'b0;
      IsNaN_5U_10U_land_4_lpi_1_dfm_4 <= 1'b0;
      IsNaN_5U_10U_land_5_lpi_1_dfm_4 <= 1'b0;
      IsNaN_5U_10U_land_6_lpi_1_dfm_4 <= 1'b0;
      IsNaN_5U_10U_land_7_lpi_1_dfm_5 <= 1'b0;
      IsNaN_5U_10U_land_8_lpi_1_dfm_4 <= 1'b0;
      IsNaN_5U_10U_land_9_lpi_1_dfm_4 <= 1'b0;
      IsNaN_5U_10U_land_10_lpi_1_dfm_4 <= 1'b0;
      IsNaN_5U_10U_land_11_lpi_1_dfm_4 <= 1'b0;
      IsNaN_5U_10U_land_12_lpi_1_dfm_4 <= 1'b0;
      IsNaN_5U_10U_land_13_lpi_1_dfm_4 <= 1'b0;
      IsNaN_5U_10U_land_14_lpi_1_dfm_5 <= 1'b0;
      IsNaN_5U_10U_land_lpi_1_dfm_4 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_9_4_1 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_9_4_1 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_9_4_1 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_9_4_1 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_9_4_1 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_9_4_1 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_9_4_1 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_9_4_1 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_9_4_1 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_9_4_1 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_9_4_1 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_9_4_1 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_9_4_1 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_9_4_1 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_9_4_1 <= 1'b0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_9_4_1 <= 1'b0;
      cfg_mode_eql_1_sva_5 <= 1'b0;
      cvt_unequal_tmp_20 <= 1'b0;
    end
    else if ( chn_idata_data_and_16_cse ) begin
      chn_idata_data_sva_2_47_31_1 <= chn_idata_data_sva_1_59_31_1[16:0];
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_9_3_0_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_7_3_0_mx0w0;
      chn_idata_data_sva_2_79_63_1 <= chn_idata_data_sva_1_91_63_1[16:0];
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_9_3_0_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_7_3_0_mx0w0;
      chn_idata_data_sva_2_111_95_1 <= chn_idata_data_sva_1_123_95_1[16:0];
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_9_3_0_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_7_3_0_mx0w0;
      chn_idata_data_sva_2_143_127_1 <= chn_idata_data_sva_1_155_127_1[16:0];
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_9_3_0_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_7_3_0_mx0w0;
      chn_idata_data_sva_2_175_159_1 <= chn_idata_data_sva_1_187_159_1[16:0];
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_9_3_0_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_7_3_0_mx0w0;
      chn_idata_data_sva_2_207_191_1 <= chn_idata_data_sva_1_219_191_1[16:0];
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_9_3_0_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_7_3_0_mx0w0;
      chn_idata_data_sva_2_239_223_1 <= chn_idata_data_sva_1_251_223_1[16:0];
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_9_3_0_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_7_3_0_mx0w0;
      chn_idata_data_sva_2_271_255_1 <= chn_idata_data_sva_1_283_255_1[16:0];
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_9_3_0_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_7_3_0_mx0w0;
      chn_idata_data_sva_2_303_287_1 <= chn_idata_data_sva_1_315_287_1[16:0];
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_9_3_0_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_7_3_0_mx0w0;
      chn_idata_data_sva_2_335_319_1 <= chn_idata_data_sva_1_347_319_1[16:0];
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_9_3_0_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_7_3_0_mx0w0;
      chn_idata_data_sva_2_367_351_1 <= chn_idata_data_sva_1_379_351_1[16:0];
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_9_3_0_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_7_3_0_mx0w0;
      chn_idata_data_sva_2_399_383_1 <= chn_idata_data_sva_1_411_383_1[16:0];
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_9_3_0_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_7_3_0_mx0w0;
      chn_idata_data_sva_2_431_415_1 <= chn_idata_data_sva_1_443_415_1[16:0];
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_9_3_0_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_7_3_0_mx0w0;
      chn_idata_data_sva_2_463_447_1 <= chn_idata_data_sva_1_475_447_1[16:0];
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_9_3_0_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_7_3_0_mx0w0;
      chn_idata_data_sva_2_495_479_1 <= chn_idata_data_sva_1_507_479_1[16:0];
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_9_3_0_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_7_3_0_mx0w0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_9_3_0_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_7_3_0_mx0w0;
      cfg_out_precision_1_sva_st_113 <= cfg_out_precision_1_sva_st_154;
      IntShiftRightSat_49U_6U_17U_o_16_1_sva_3 <= IntShiftRightSat_49U_6U_17U_o_16_1_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_0_1_sva_2 <= IntShiftRightSat_49U_6U_17U_o_0_1_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_0_2_sva_2 <= IntShiftRightSat_49U_6U_17U_o_0_2_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_16_3_sva_3 <= IntShiftRightSat_49U_6U_17U_o_16_3_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_0_3_sva_3 <= IntShiftRightSat_49U_6U_17U_o_0_3_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_0_4_sva_2 <= IntShiftRightSat_49U_6U_17U_o_0_4_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_16_5_sva_3 <= IntShiftRightSat_49U_6U_17U_o_16_5_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_0_5_sva_3 <= IntShiftRightSat_49U_6U_17U_o_0_5_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_0_6_sva_2 <= IntShiftRightSat_49U_6U_17U_o_0_6_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_0_7_sva_2 <= IntShiftRightSat_49U_6U_17U_o_0_7_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_0_8_sva_2 <= IntShiftRightSat_49U_6U_17U_o_0_8_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_16_9_sva_3 <= IntShiftRightSat_49U_6U_17U_o_16_9_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_0_9_sva_3 <= IntShiftRightSat_49U_6U_17U_o_0_9_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_0_10_sva_2 <= IntShiftRightSat_49U_6U_17U_o_0_10_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_0_11_sva_2 <= IntShiftRightSat_49U_6U_17U_o_0_11_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_0_12_sva_2 <= IntShiftRightSat_49U_6U_17U_o_0_12_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_0_13_sva_2 <= IntShiftRightSat_49U_6U_17U_o_0_13_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_0_14_sva_3 <= IntShiftRightSat_49U_6U_17U_o_0_14_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_0_15_sva_2 <= IntShiftRightSat_49U_6U_17U_o_0_15_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_0_sva_2 <= IntShiftRightSat_49U_6U_17U_o_0_sva_mx0w0;
      cfg_proc_precision_1_sva_st_65 <= cfg_proc_precision_1_sva_st_64;
      IsNaN_5U_10U_land_3_lpi_1_dfm_4 <= ~((~((FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_3_lpi_1_dfm_5_mx0!=10'b0000000000)))
          | (~(FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_7_4_mx0w0 & (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_7_3_0_mx0w0==4'b1111))));
      IsNaN_5U_10U_land_4_lpi_1_dfm_4 <= ~((~((FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_4_lpi_1_dfm_5_mx0!=10'b0000000000)))
          | (~(FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_7_4_mx0w0 & (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_7_3_0_mx0w0==4'b1111))));
      IsNaN_5U_10U_land_5_lpi_1_dfm_4 <= ~((~((FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_5_lpi_1_dfm_5_mx0!=10'b0000000000)))
          | (~(FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_7_4_mx0w0 & (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_7_3_0_mx0w0==4'b1111))));
      IsNaN_5U_10U_land_6_lpi_1_dfm_4 <= ~((~((FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_6_lpi_1_dfm_5_mx0!=10'b0000000000)))
          | (~(FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_7_4_mx0w0 & (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_7_3_0_mx0w0==4'b1111))));
      IsNaN_5U_10U_land_7_lpi_1_dfm_5 <= ~((~((FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_7_lpi_1_dfm_5_mx0!=10'b0000000000)))
          | (~(FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_7_4_mx0w0 & (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_7_3_0_mx0w0==4'b1111))));
      IsNaN_5U_10U_land_8_lpi_1_dfm_4 <= ~((~((FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_8_lpi_1_dfm_5_mx0!=10'b0000000000)))
          | (~(FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_7_4_mx0w0 & (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_7_3_0_mx0w0==4'b1111))));
      IsNaN_5U_10U_land_9_lpi_1_dfm_4 <= ~((~((FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_9_lpi_1_dfm_5_mx0!=10'b0000000000)))
          | (~(FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_7_4_mx0w0 & (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_7_3_0_mx0w0==4'b1111))));
      IsNaN_5U_10U_land_10_lpi_1_dfm_4 <= ~((~((FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_10_lpi_1_dfm_5_mx0!=10'b0000000000)))
          | (~(FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_7_4_mx0w0 & (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_7_3_0_mx0w0==4'b1111))));
      IsNaN_5U_10U_land_11_lpi_1_dfm_4 <= ~((~((FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_11_lpi_1_dfm_5_mx0!=10'b0000000000)))
          | (~(FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_7_4_mx0w0 & (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_7_3_0_mx0w0==4'b1111))));
      IsNaN_5U_10U_land_12_lpi_1_dfm_4 <= ~((~((FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_12_lpi_1_dfm_5_mx0!=10'b0000000000)))
          | (~(FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_7_4_mx0w0 & (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_7_3_0_mx0w0==4'b1111))));
      IsNaN_5U_10U_land_13_lpi_1_dfm_4 <= ~((~((FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_13_lpi_1_dfm_5_mx0!=10'b0000000000)))
          | (~(FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_7_4_mx0w0 & (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_7_3_0_mx0w0==4'b1111))));
      IsNaN_5U_10U_land_14_lpi_1_dfm_5 <= ~((~((FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_14_lpi_1_dfm_5_mx0!=10'b0000000000)))
          | (~(FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_7_4_mx0w0 & (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_7_3_0_mx0w0==4'b1111))));
      IsNaN_5U_10U_land_lpi_1_dfm_4 <= ~((~((FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_lpi_1_dfm_5_mx0!=10'b0000000000)))
          | (~(FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_7_4_mx0w0 & (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_7_3_0_mx0w0==4'b1111))));
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_9_4_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_7_4_mx0w0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_9_4_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_7_4_mx0w0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_9_4_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_7_4_mx0w0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_9_4_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_7_4_mx0w0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_9_4_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_7_4_mx0w0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_9_4_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_7_4_mx0w0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_9_4_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_7_4_mx0w0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_9_4_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_7_4_mx0w0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_9_4_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_7_4_mx0w0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_9_4_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_7_4_mx0w0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_9_4_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_7_4_mx0w0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_9_4_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_7_4_mx0w0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_9_4_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_7_4_mx0w0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_9_4_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_7_4_mx0w0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_9_4_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_7_4_mx0w0;
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_9_4_1 <= FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_7_4_mx0w0;
      cfg_mode_eql_1_sva_5 <= cfg_mode_eql_1_sva_4;
      cvt_unequal_tmp_20 <= cvt_unequal_tmp_19;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_1_lpi_1_dfm_8 <= 10'b0;
    end
    else if ( core_wen & ((or_5189_cse & IsNaN_8U_23U_land_1_lpi_1_dfm_3) | and_637_rgt)
        & mux_tmp_161 ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_1_lpi_1_dfm_8 <= MUX_v_10_2_2((chn_idata_data_sva_1_27_0_1[9:0]),
          FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_mx0w1,
          and_637_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_1_FpFloatToInt_16U_5U_10U_shift_acc_itm_2 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_162_nl) ) begin
      cvt_1_FpFloatToInt_16U_5U_10U_shift_acc_itm_2 <= nl_cvt_1_FpFloatToInt_16U_5U_10U_shift_acc_itm_2[4:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_2_lpi_1_dfm_8 <= 10'b0;
    end
    else if ( core_wen & ((or_5189_cse & IsNaN_8U_23U_land_2_lpi_1_dfm_3) | and_639_rgt)
        & mux_tmp_161 ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_2_lpi_1_dfm_8 <= MUX_v_10_2_2((chn_idata_data_sva_1_59_31_1[10:1]),
          FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_1_mx0w1,
          and_639_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_2_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2 <= 5'b0;
      cvt_3_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2 <= 5'b0;
      cvt_4_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 <= 5'b0;
    end
    else if ( FpFloatToInt_16U_5U_10U_shift_and_1_cse ) begin
      cvt_2_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2 <= nl_cvt_2_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2[4:0];
      cvt_3_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2 <= nl_cvt_3_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2[4:0];
      cvt_4_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 <= nl_cvt_4_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2[4:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_3_lpi_1_dfm_8 <= 10'b0;
    end
    else if ( core_wen & ((or_5189_cse & IsNaN_8U_23U_land_3_lpi_1_dfm_3) | and_641_rgt)
        & mux_tmp_161 ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_3_lpi_1_dfm_8 <= MUX_v_10_2_2((chn_idata_data_sva_1_91_63_1[10:1]),
          FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_2_mx0w1,
          and_641_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_4_lpi_1_dfm_8 <= 10'b0;
    end
    else if ( core_wen & ((or_5189_cse & IsNaN_8U_23U_land_4_lpi_1_dfm_3) | and_643_rgt)
        & mux_tmp_161 ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_4_lpi_1_dfm_8 <= MUX_v_10_2_2((chn_idata_data_sva_1_123_95_1[10:1]),
          FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_3_mx0w1,
          and_643_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_5_lpi_1_dfm_8 <= 10'b0;
    end
    else if ( core_wen & ((nor_1099_cse & or_5189_cse) | and_646_rgt) & mux_tmp_161
        ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_5_lpi_1_dfm_8 <= MUX_v_10_2_2((chn_idata_data_sva_1_155_127_1[10:1]),
          FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_4_mx0w1,
          and_646_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_5_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_167_nl)) ) begin
      cvt_5_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2 <= nl_cvt_5_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2[4:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_6_lpi_1_dfm_8 <= 10'b0;
    end
    else if ( core_wen & ((or_5189_cse & IsNaN_8U_23U_land_6_lpi_1_dfm_3) | and_648_rgt)
        & mux_tmp_161 ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_6_lpi_1_dfm_8 <= MUX_v_10_2_2((chn_idata_data_sva_1_187_159_1[10:1]),
          FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_5_mx0w1,
          and_648_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_6_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 <= 5'b0;
      cvt_7_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 <= 5'b0;
      cvt_8_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2 <= 5'b0;
      cvt_10_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 <= 5'b0;
      cvt_11_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 <= 5'b0;
      cvt_13_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 <= 5'b0;
      cvt_15_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2 <= 5'b0;
    end
    else if ( FpFloatToInt_16U_5U_10U_shift_and_5_cse ) begin
      cvt_6_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 <= nl_cvt_6_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2[4:0];
      cvt_7_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 <= nl_cvt_7_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2[4:0];
      cvt_8_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2 <= nl_cvt_8_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2[4:0];
      cvt_10_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 <= nl_cvt_10_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2[4:0];
      cvt_11_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 <= nl_cvt_11_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2[4:0];
      cvt_13_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 <= nl_cvt_13_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2[4:0];
      cvt_15_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2 <= nl_cvt_15_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2[4:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_7_lpi_1_dfm_8 <= 10'b0;
    end
    else if ( core_wen & ((or_5189_cse & IsNaN_8U_23U_land_7_lpi_1_dfm_3) | and_650_rgt)
        & mux_tmp_161 ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_7_lpi_1_dfm_8 <= MUX_v_10_2_2((chn_idata_data_sva_1_219_191_1[10:1]),
          FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_6_mx0w1,
          and_650_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_8_lpi_1_dfm_8 <= 10'b0;
    end
    else if ( core_wen & ((or_5189_cse & IsNaN_8U_23U_land_8_lpi_1_dfm_3) | and_652_rgt)
        & mux_tmp_161 ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_8_lpi_1_dfm_8 <= MUX_v_10_2_2((chn_idata_data_sva_1_251_223_1[10:1]),
          FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_7_mx0w1,
          and_652_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_9_lpi_1_dfm_8 <= 10'b0;
    end
    else if ( core_wen & ((or_5189_cse & IsNaN_8U_23U_land_9_lpi_1_dfm_3) | and_654_rgt)
        & mux_tmp_161 ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_9_lpi_1_dfm_8 <= MUX_v_10_2_2((chn_idata_data_sva_1_283_255_1[10:1]),
          FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_8_mx0w1,
          and_654_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_9_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2 <= 5'b0;
      cvt_12_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2 <= 5'b0;
      cvt_14_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2 <= 5'b0;
    end
    else if ( FpFloatToInt_16U_5U_10U_shift_and_8_cse ) begin
      cvt_9_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2 <= nl_cvt_9_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2[4:0];
      cvt_12_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2 <= nl_cvt_12_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2[4:0];
      cvt_14_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2 <= nl_cvt_14_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2[4:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_10_lpi_1_dfm_8 <= 10'b0;
    end
    else if ( core_wen & ((or_5189_cse & IsNaN_8U_23U_land_10_lpi_1_dfm_3) | and_656_rgt)
        & mux_tmp_161 ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_10_lpi_1_dfm_8 <= MUX_v_10_2_2((chn_idata_data_sva_1_315_287_1[10:1]),
          FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_9_mx0w1,
          and_656_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_11_lpi_1_dfm_8 <= 10'b0;
    end
    else if ( core_wen & ((or_5189_cse & IsNaN_8U_23U_land_11_lpi_1_dfm_3) | and_658_rgt)
        & mux_tmp_161 ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_11_lpi_1_dfm_8 <= MUX_v_10_2_2((chn_idata_data_sva_1_347_319_1[10:1]),
          FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_10_mx0w1,
          and_658_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_12_lpi_1_dfm_8 <= 10'b0;
    end
    else if ( core_wen & ((or_5189_cse & IsNaN_8U_23U_land_12_lpi_1_dfm_3) | and_660_rgt)
        & mux_tmp_161 ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_12_lpi_1_dfm_8 <= MUX_v_10_2_2((chn_idata_data_sva_1_379_351_1[10:1]),
          FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_11_mx0w1,
          and_660_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_13_lpi_1_dfm_8 <= 10'b0;
    end
    else if ( core_wen & ((or_5189_cse & IsNaN_8U_23U_land_13_lpi_1_dfm_3) | and_662_rgt)
        & mux_tmp_161 ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_13_lpi_1_dfm_8 <= MUX_v_10_2_2((chn_idata_data_sva_1_411_383_1[10:1]),
          FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_12_mx0w1,
          and_662_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_14_lpi_1_dfm_8 <= 10'b0;
    end
    else if ( core_wen & ((or_5189_cse & IsNaN_8U_23U_land_14_lpi_1_dfm_3) | and_664_rgt)
        & mux_tmp_161 ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_14_lpi_1_dfm_8 <= MUX_v_10_2_2((chn_idata_data_sva_1_443_415_1[10:1]),
          FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_13_mx0w1,
          and_664_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_15_lpi_1_dfm_8 <= 10'b0;
    end
    else if ( core_wen & ((or_5189_cse & IsNaN_8U_23U_land_15_lpi_1_dfm_3) | and_666_rgt)
        & mux_tmp_161 ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_15_lpi_1_dfm_8 <= MUX_v_10_2_2((chn_idata_data_sva_1_475_447_1[10:1]),
          FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_14_mx0w1,
          and_666_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_idata_data_sva_2_511_1 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_191_nl)) ) begin
      chn_idata_data_sva_2_511_1 <= chn_idata_data_sva_1_511_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_lpi_1_dfm_9 <= 10'b0;
    end
    else if ( core_wen & ((or_5189_cse & IsNaN_8U_23U_land_lpi_1_dfm_3) | and_668_rgt)
        & mux_tmp_161 ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_lpi_1_dfm_9 <= MUX_v_10_2_2((chn_idata_data_sva_1_507_479_1[10:1]),
          FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_2_nor_15_mx0w1,
          and_668_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_16_FpFloatToInt_16U_5U_10U_shift_acc_4_itm_2 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_192_nl)) ) begin
      cvt_16_FpFloatToInt_16U_5U_10U_shift_acc_4_itm_2 <= nl_cvt_16_FpFloatToInt_16U_5U_10U_shift_acc_4_itm_2[4:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_i_1_sva_2 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_235_nl) ) begin
      IntShiftRightSat_49U_6U_17U_i_1_sva_2 <= IntShiftRightSat_49U_6U_17U_i_1_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_2 <= 15'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_27_cse
        & (mux_243_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_2 <= MUX_v_15_2_2(IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_15_1_1_sva, and_dcpl_4);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_15_1_1_lpi_1_dfm_5 <= 15'b0;
      FpIntToFloat_17U_5U_10U_else_i_abs_0_1_lpi_1_dfm_5 <= 1'b0;
    end
    else if ( FpIntToFloat_17U_5U_10U_else_i_abs_and_cse ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_15_1_1_lpi_1_dfm_5 <= MUX_v_15_2_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_1_sva[15:1]),
          IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_mx0w0, and_dcpl_209);
      FpIntToFloat_17U_5U_10U_else_i_abs_0_1_lpi_1_dfm_5 <= MUX_s_1_2_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_1_sva[0]),
          IntShiftRightSat_49U_6U_17U_o_0_1_sva_mx0w0, and_dcpl_209);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_1_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ mux_tmp_245) ) begin
      cvt_1_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_itm_2
          <= FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_1_sva[16];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_svs_st_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_247_nl) ) begin
      cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_svs_st_2 <= cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_i_2_sva_2 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_248_nl) ) begin
      IntShiftRightSat_49U_6U_17U_i_2_sva_2 <= IntShiftRightSat_49U_6U_17U_i_2_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_16_2_sva_2 <= 1'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
        & (mux_257_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_16_2_sva_2 <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_16_2_sva, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_2 <= 15'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
        & (mux_267_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_2 <= MUX_v_15_2_2(IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_15_1_2_sva, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_15_1_2_lpi_1_dfm_6 <= 15'b0;
      FpIntToFloat_17U_5U_10U_else_i_abs_0_2_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( FpIntToFloat_17U_5U_10U_else_i_abs_and_13_cse ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_15_1_2_lpi_1_dfm_6 <= MUX_v_15_2_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_2_sva[15:1]),
          IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_mx0w0, and_dcpl_217);
      FpIntToFloat_17U_5U_10U_else_i_abs_0_2_lpi_1_dfm_6 <= MUX_s_1_2_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_2_sva[0]),
          IntShiftRightSat_49U_6U_17U_o_0_2_sva_mx0w0, and_dcpl_217);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_2_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & not_tmp_249 ) begin
      cvt_2_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2
          <= FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_2_sva[16];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 <=
          1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_271_nl) ) begin
      cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 <=
          cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2
          <= 1'b0;
      cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2
          <= 1'b0;
    end
    else if ( IntShiftRightSat_49U_6U_17U_if_and_cse ) begin
      cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2
          <= cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp;
      cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2
          <= cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_i_3_sva_2 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_275_nl) ) begin
      IntShiftRightSat_49U_6U_17U_i_3_sva_2 <= IntShiftRightSat_49U_6U_17U_i_3_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_2 <= 15'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
        & (mux_285_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_2 <= MUX_v_15_2_2(IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_15_1_3_sva, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_15_1_3_lpi_1_dfm_6 <= 15'b0;
      FpIntToFloat_17U_5U_10U_else_i_abs_0_3_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( FpIntToFloat_17U_5U_10U_else_i_abs_and_15_cse ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_15_1_3_lpi_1_dfm_6 <= MUX_v_15_2_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_3_sva[15:1]),
          IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_mx0w0, and_dcpl_224);
      FpIntToFloat_17U_5U_10U_else_i_abs_0_3_lpi_1_dfm_6 <= MUX_s_1_2_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_3_sva[0]),
          IntShiftRightSat_49U_6U_17U_o_0_3_sva_mx0w0, and_dcpl_224);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_3_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & not_tmp_269 ) begin
      cvt_3_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2
          <= FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_3_sva[16];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 <=
          1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_289_nl) ) begin
      cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 <=
          cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_i_4_sva_2 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_291_nl) ) begin
      IntShiftRightSat_49U_6U_17U_i_4_sva_2 <= IntShiftRightSat_49U_6U_17U_i_4_sva_mx0w1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_16_4_sva_2 <= 1'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
        & (mux_302_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_16_4_sva_2 <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_16_4_sva, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_2 <= 15'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
        & (mux_316_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_2 <= MUX_v_15_2_2(IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_15_1_4_sva, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_4_lpi_1_dfm_6_reg <= 5'b0;
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_5_lpi_1_dfm_5_reg <= 5'b0;
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_6_lpi_1_dfm_6_reg <= 5'b0;
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_7_lpi_1_dfm_6_reg <= 5'b0;
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_8_lpi_1_dfm_7_reg <= 5'b0;
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_10_lpi_1_dfm_6_reg <= 5'b0;
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_11_lpi_1_dfm_6_reg <= 5'b0;
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_12_lpi_1_dfm_7_reg <= 5'b0;
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_13_lpi_1_dfm_6_reg <= 5'b0;
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_15_lpi_1_dfm_7_reg <= 5'b0;
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_lpi_1_dfm_8_reg <= 5'b0;
    end
    else if ( and_2257_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_4_lpi_1_dfm_6_reg <= FpIntToFloat_17U_5U_10U_else_if_mux1h_9_rgt[14:10];
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_5_lpi_1_dfm_5_reg <= FpIntToFloat_17U_5U_10U_else_if_mux1h_12_rgt[14:10];
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_6_lpi_1_dfm_6_reg <= FpIntToFloat_17U_5U_10U_else_if_mux1h_15_rgt[14:10];
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_7_lpi_1_dfm_6_reg <= FpIntToFloat_17U_5U_10U_else_if_mux1h_18_rgt[14:10];
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_8_lpi_1_dfm_7_reg <= FpIntToFloat_17U_5U_10U_else_if_mux1h_21_rgt[14:10];
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_10_lpi_1_dfm_6_reg <= FpIntToFloat_17U_5U_10U_else_if_mux1h_27_rgt[14:10];
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_11_lpi_1_dfm_6_reg <= FpIntToFloat_17U_5U_10U_else_if_mux1h_30_rgt[14:10];
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_12_lpi_1_dfm_7_reg <= FpIntToFloat_17U_5U_10U_else_if_mux1h_33_rgt[14:10];
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_13_lpi_1_dfm_6_reg <= FpIntToFloat_17U_5U_10U_else_if_mux1h_36_rgt[14:10];
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_15_lpi_1_dfm_7_reg <= FpIntToFloat_17U_5U_10U_else_if_mux1h_41_rgt[14:10];
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_lpi_1_dfm_8_reg <= FpIntToFloat_17U_5U_10U_else_if_mux1h_44_rgt[14:10];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_4_lpi_1_dfm_6_1_reg <= 10'b0;
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_10_lpi_1_dfm_6_1_reg <= 10'b0;
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_11_lpi_1_dfm_6_1_reg <= 10'b0;
    end
    else if ( and_2259_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_4_lpi_1_dfm_6_1_reg <= FpIntToFloat_17U_5U_10U_else_if_mux1h_9_rgt[9:0];
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_10_lpi_1_dfm_6_1_reg <= FpIntToFloat_17U_5U_10U_else_if_mux1h_27_rgt[9:0];
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_11_lpi_1_dfm_6_1_reg <= FpIntToFloat_17U_5U_10U_else_if_mux1h_30_rgt[9:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_0_4_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & (~ cvt_4_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp)
        & or_dcpl_108) | and_704_rgt) & not_tmp_312 ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_0_4_lpi_1_dfm_7 <= MUX_s_1_2_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_4_sva[0]),
          IntShiftRightSat_49U_6U_17U_o_0_4_sva_mx0w0, and_704_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_4_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & not_tmp_312 ) begin
      cvt_4_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2
          <= FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_4_sva[16];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_322_nl) ) begin
      cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2
          <= cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_i_5_sva_2 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_329_nl) ) begin
      IntShiftRightSat_49U_6U_17U_i_5_sva_2 <= IntShiftRightSat_49U_6U_17U_i_5_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_2 <= 15'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
        & (mux_338_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_2 <= MUX_v_15_2_2(IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_15_1_5_sva, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_5_lpi_1_dfm_5_1_reg <= 10'b0;
    end
    else if ( (~((mux_2176_nl) | nor_2040_cse)) & core_wen ) begin
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_5_lpi_1_dfm_5_1_reg <= FpIntToFloat_17U_5U_10U_else_if_mux1h_12_rgt[9:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_0_5_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & (~ cvt_5_IntShiftRight_49U_6U_17U_obits_fixed_nor_5_tmp)
        & or_dcpl_110) | and_719_rgt) & not_tmp_336 ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_0_5_lpi_1_dfm_6 <= MUX_s_1_2_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_5_sva[0]),
          IntShiftRightSat_49U_6U_17U_o_0_5_sva_mx0w0, and_719_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_5_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & not_tmp_336 ) begin
      cvt_5_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2
          <= FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_5_sva[16];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 <=
          1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_342_nl) ) begin
      cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 <=
          cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_i_6_sva_2 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_348_nl) ) begin
      IntShiftRightSat_49U_6U_17U_i_6_sva_2 <= IntShiftRightSat_49U_6U_17U_i_6_sva_mx0w1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_16_6_sva_2 <= 1'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
        & (mux_359_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_16_6_sva_2 <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_16_6_sva, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_2 <= 15'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
        & (mux_373_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_2 <= MUX_v_15_2_2(IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_15_1_6_sva, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_6_lpi_1_dfm_6_1_reg <= 10'b0;
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_7_lpi_1_dfm_6_1_reg <= 10'b0;
    end
    else if ( and_2275_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_6_lpi_1_dfm_6_1_reg <= FpIntToFloat_17U_5U_10U_else_if_mux1h_15_rgt[9:0];
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_7_lpi_1_dfm_6_1_reg <= FpIntToFloat_17U_5U_10U_else_if_mux1h_18_rgt[9:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_0_6_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & (~ cvt_6_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp)
        & or_dcpl_113) | and_734_rgt) & not_tmp_388 ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_0_6_lpi_1_dfm_7 <= MUX_s_1_2_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_6_sva[0]),
          IntShiftRightSat_49U_6U_17U_o_0_6_sva_mx0w0, and_734_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_6_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & not_tmp_388 ) begin
      cvt_6_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2
          <= FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_6_sva[16];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2
          <= 1'b0;
      cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2
          <= 1'b0;
    end
    else if ( IntShiftRightSat_49U_6U_17U_if_and_3_cse ) begin
      cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2
          <= cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp;
      cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2
          <= cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_i_7_sva_2 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_383_nl) ) begin
      IntShiftRightSat_49U_6U_17U_i_7_sva_2 <= IntShiftRightSat_49U_6U_17U_i_7_sva_mx0w1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_16_7_sva_2 <= 1'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
        & (mux_394_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_16_7_sva_2 <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_16_7_sva, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_2 <= 15'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
        & (mux_408_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_2 <= MUX_v_15_2_2(IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_15_1_7_sva, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_0_7_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & (~ cvt_7_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp)
        & or_dcpl_115) | and_749_rgt) & not_tmp_436 ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_0_7_lpi_1_dfm_7 <= MUX_s_1_2_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_7_sva[0]),
          IntShiftRightSat_49U_6U_17U_o_0_7_sva_mx0w0, and_749_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_7_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & not_tmp_436 ) begin
      cvt_7_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2
          <= FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_7_sva[16];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_i_8_sva_2 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_418_nl) ) begin
      IntShiftRightSat_49U_6U_17U_i_8_sva_2 <= IntShiftRightSat_49U_6U_17U_i_8_sva_mx0w1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_16_8_sva_2 <= 1'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
        & (mux_431_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_16_8_sva_2 <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_16_8_sva, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_2 <= 15'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
        & (mux_444_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_2 <= MUX_v_15_2_2(IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_15_1_8_sva, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_8_lpi_1_dfm_7_1_reg <= 10'b0;
    end
    else if ( (~((mux_2186_nl) | nor_2040_cse)) & core_wen ) begin
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_8_lpi_1_dfm_7_1_reg <= FpIntToFloat_17U_5U_10U_else_if_mux1h_21_rgt[9:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_0_8_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & (~ cvt_8_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp)
        & or_dcpl_119) | and_766_rgt) & not_tmp_497 ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_0_8_lpi_1_dfm_8 <= MUX_s_1_2_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_8_sva[0]),
          IntShiftRightSat_49U_6U_17U_o_0_8_sva_mx0w0, and_766_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_8_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & not_tmp_497 ) begin
      cvt_8_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2
          <= FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_8_sva[16];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_450_nl) ) begin
      cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_svs_st_2
          <= cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_453_nl) ) begin
      cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2
          <= cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_i_9_sva_2 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_458_nl) ) begin
      IntShiftRightSat_49U_6U_17U_i_9_sva_2 <= IntShiftRightSat_49U_6U_17U_i_9_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_2 <= 15'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
        & (mux_467_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_2 <= MUX_v_15_2_2(IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_15_1_9_sva, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_15_1_9_lpi_1_dfm_6 <= 15'b0;
      FpIntToFloat_17U_5U_10U_else_i_abs_0_9_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( FpIntToFloat_17U_5U_10U_else_i_abs_and_22_cse ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_15_1_9_lpi_1_dfm_6 <= MUX_v_15_2_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_9_sva[15:1]),
          IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_mx0w0, and_dcpl_301);
      FpIntToFloat_17U_5U_10U_else_i_abs_0_9_lpi_1_dfm_6 <= MUX_s_1_2_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_9_sva[0]),
          IntShiftRightSat_49U_6U_17U_o_0_9_sva_mx0w0, and_dcpl_301);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_9_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & not_tmp_520 ) begin
      cvt_9_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_1_itm_2
          <= FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_9_sva[16];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 <=
          1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_472_nl) ) begin
      cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 <=
          cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_i_10_sva_2 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_478_nl) ) begin
      IntShiftRightSat_49U_6U_17U_i_10_sva_2 <= IntShiftRightSat_49U_6U_17U_i_10_sva_mx0w1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_16_10_sva_2 <= 1'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
        & (mux_490_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_16_10_sva_2 <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_16_10_sva, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_2 <= 15'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
        & (mux_505_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_2 <= MUX_v_15_2_2(IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_15_1_10_sva, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_0_10_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & (~ cvt_10_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp)
        & or_dcpl_124) | and_787_rgt) & not_tmp_580 ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_0_10_lpi_1_dfm_7 <= MUX_s_1_2_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_10_sva[0]),
          IntShiftRightSat_49U_6U_17U_o_0_10_sva_mx0w0, and_787_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_10_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & not_tmp_580 ) begin
      cvt_10_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2
          <= FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_10_sva[16];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_i_11_sva_2 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_516_nl) ) begin
      IntShiftRightSat_49U_6U_17U_i_11_sva_2 <= IntShiftRightSat_49U_6U_17U_i_11_sva_mx0w1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_16_11_sva_2 <= 1'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
        & (mux_528_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_16_11_sva_2 <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_16_11_sva, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_2 <= 15'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
        & (mux_544_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_2 <= MUX_v_15_2_2(IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_15_1_11_sva, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_0_11_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & (~ cvt_11_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp)
        & or_dcpl_126) | and_801_rgt) & not_tmp_638 ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_0_11_lpi_1_dfm_7 <= MUX_s_1_2_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_11_sva[0]),
          IntShiftRightSat_49U_6U_17U_o_0_11_sva_mx0w0, and_801_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_11_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & not_tmp_638 ) begin
      cvt_11_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2
          <= FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_11_sva[16];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_i_12_sva_2 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_556_nl) ) begin
      IntShiftRightSat_49U_6U_17U_i_12_sva_2 <= IntShiftRightSat_49U_6U_17U_i_12_sva_mx0w1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_16_12_sva_2 <= 1'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
        & (mux_569_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_16_12_sva_2 <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_16_12_sva, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_2 <= 15'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
        & (mux_583_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_2 <= MUX_v_15_2_2(IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_15_1_12_sva, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_12_lpi_1_dfm_7_1_reg <= 10'b0;
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_13_lpi_1_dfm_6_1_reg <= 10'b0;
    end
    else if ( and_2317_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_12_lpi_1_dfm_7_1_reg <= FpIntToFloat_17U_5U_10U_else_if_mux1h_33_rgt[9:0];
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_13_lpi_1_dfm_6_1_reg <= FpIntToFloat_17U_5U_10U_else_if_mux1h_36_rgt[9:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_0_12_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & (~ cvt_12_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp)
        & or_dcpl_130) | and_816_rgt) & (~ mux_tmp_585) ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_0_12_lpi_1_dfm_8 <= MUX_s_1_2_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_12_sva[0]),
          IntShiftRightSat_49U_6U_17U_o_0_12_sva_mx0w0, and_816_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_12_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ mux_tmp_585) ) begin
      cvt_12_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2
          <= FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_12_sva[16];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_i_13_sva_2 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_594_nl) ) begin
      IntShiftRightSat_49U_6U_17U_i_13_sva_2 <= IntShiftRightSat_49U_6U_17U_i_13_sva_mx0w1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_16_13_sva_2 <= 1'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
        & (mux_605_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_16_13_sva_2 <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_16_13_sva, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_2 <= 15'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
        & (mux_617_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_2 <= MUX_v_15_2_2(IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_15_1_13_sva, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_0_13_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & (~ cvt_13_IntShiftRight_49U_6U_17U_obits_fixed_nor_10_tmp)
        & or_dcpl_132) | and_830_rgt) & not_tmp_757 ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_0_13_lpi_1_dfm_7 <= MUX_s_1_2_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_13_sva[0]),
          IntShiftRightSat_49U_6U_17U_o_0_13_sva_mx0w0, and_830_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_13_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & not_tmp_757 ) begin
      cvt_13_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_2_itm_2
          <= FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_13_sva[16];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_i_14_sva_2 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_630_nl) ) begin
      IntShiftRightSat_49U_6U_17U_i_14_sva_2 <= IntShiftRightSat_49U_6U_17U_i_14_sva_mx0w1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_16_14_sva_2 <= 1'b0;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm_3 <= 1'b0;
    end
    else if ( IntShiftRightSat_49U_6U_17U_o_and_90_cse ) begin
      IntShiftRightSat_49U_6U_17U_o_16_14_sva_2 <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_16_14_sva, and_685_rgt);
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm_3 <= MUX_s_1_2_2(IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm_mx0w0,
          IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_2 <= 15'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
        & (mux_644_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_2 <= MUX_v_15_2_2(IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_15_1_14_sva, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_14_lpi_1_dfm_7_reg <= 5'b0;
    end
    else if ( or_4550_cse & or_183_cse_1 & or_5189_cse & main_stage_v_1 & (cfg_out_precision_1_sva_st_154==2'b10)
        & core_wen ) begin
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_14_lpi_1_dfm_7_reg <= FpIntToFloat_17U_5U_10U_else_i_abs_mux1h_17_rgt[14:10];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_14_lpi_1_dfm_7_1_reg <= 10'b0;
    end
    else if ( ((mux_2214_nl) | (fsm_output[0])) & core_wen ) begin
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_14_lpi_1_dfm_7_1_reg <= FpIntToFloat_17U_5U_10U_else_i_abs_mux1h_17_rgt[9:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_0_14_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & (~ cvt_14_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp)
        & or_dcpl_136) | and_849_rgt) & not_tmp_811 ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_0_14_lpi_1_dfm_8 <= MUX_s_1_2_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_14_sva[0]),
          IntShiftRightSat_49U_6U_17U_o_0_14_sva_mx0w0, and_849_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_14_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & not_tmp_811 ) begin
      cvt_14_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2
          <= FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_14_sva[16];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_i_15_sva_2 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_671_nl) ) begin
      IntShiftRightSat_49U_6U_17U_i_15_sva_2 <= IntShiftRightSat_49U_6U_17U_i_15_sva_mx0w1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_16_15_sva_2 <= 1'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
        & (mux_684_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_16_15_sva_2 <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_16_15_sva, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_2 <= 15'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
        & (mux_698_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_2 <= MUX_v_15_2_2(IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_15_1_15_sva, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_15_lpi_1_dfm_7_1_reg <= 10'b0;
    end
    else if ( (~((mux_2218_nl) | nor_2040_cse)) & core_wen ) begin
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_15_lpi_1_dfm_7_1_reg <= FpIntToFloat_17U_5U_10U_else_if_mux1h_41_rgt[9:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_0_15_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & (~ cvt_15_IntShiftRight_49U_6U_17U_obits_fixed_nor_15_tmp)
        & or_dcpl_139) | and_866_rgt) & not_tmp_899 ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_0_15_lpi_1_dfm_8 <= MUX_s_1_2_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_15_sva[0]),
          IntShiftRightSat_49U_6U_17U_o_0_15_sva_mx0w0, and_866_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_15_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & not_tmp_899 ) begin
      cvt_15_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_3_itm_2
          <= FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_15_sva[16];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_i_sva_2 <= 49'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_715_nl) ) begin
      IntShiftRightSat_49U_6U_17U_i_sva_2 <= IntShiftRightSat_49U_6U_17U_i_sva_mx0w1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_16_sva_2 <= 1'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
        & (mux_730_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_16_sva_2 <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_16_sva, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_sva_2 <= 15'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_26_cse
        & (mux_746_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_sva_2 <= MUX_v_15_2_2(IntShiftRightSat_49U_6U_17U_o_15_1_sva_mx0w0,
          IntShiftRightSat_49U_6U_17U_o_15_1_sva, and_685_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_lpi_1_dfm_8_1_reg <= 10'b0;
    end
    else if ( (~((mux_2223_nl) | nor_2040_cse)) & core_wen ) begin
      reg_FpIntToFloat_17U_5U_10U_else_i_abs_15_1_lpi_1_dfm_8_1_reg <= FpIntToFloat_17U_5U_10U_else_if_mux1h_44_rgt[9:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_0_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & (~ cvt_16_IntShiftRight_49U_6U_17U_obits_fixed_nor_20_tmp)
        & or_dcpl_143) | and_881_rgt) & not_tmp_989 ) begin
      FpIntToFloat_17U_5U_10U_else_i_abs_0_lpi_1_dfm_9 <= MUX_s_1_2_2((FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_sva[0]),
          IntShiftRightSat_49U_6U_17U_o_0_sva_mx0w0, and_881_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_16_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_4_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & not_tmp_989 ) begin
      cvt_16_FpIntToFloat_17U_5U_10U_else_if_slc_FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_16_4_itm_2
          <= FpIntToFloat_17U_5U_10U_else_if_ac_int_cctor_sva[16];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_out_precision_1_sva_st_149 <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_794_nl) ) begin
      cfg_out_precision_1_sva_st_149 <= cfg_out_precision_1_sva_st_154;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_proc_precision_1_sva_st_101 <= 2'b0;
      cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_2
          <= 1'b0;
    end
    else if ( cfg_proc_precision_and_24_cse ) begin
      cfg_proc_precision_1_sva_st_101 <= reg_cfg_proc_precision_1_sva_st_40_cse;
      cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_2
          <= cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_proc_precision_1_sva_st_89 <= 2'b0;
      cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_svs_2
          <= 1'b0;
    end
    else if ( cfg_proc_precision_and_27_cse ) begin
      cfg_proc_precision_1_sva_st_89 <= reg_cfg_proc_precision_1_sva_st_40_cse;
      cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_svs_2
          <= cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_3 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_401 | main_stage_v_3_mx0c1) ) begin
      main_stage_v_3 <= ~ main_stage_v_3_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_2 <= 1'b0;
      FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_2 <= 1'b0;
      FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_2 <= 1'b0;
      FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_2 <= 1'b0;
      FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_2 <= 1'b0;
      FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_2 <= 1'b0;
      FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_2 <= 1'b0;
      FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_2 <= 1'b0;
      FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_2 <= 1'b0;
      FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_2 <= 1'b0;
      FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_2 <= 1'b0;
      FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_2 <= 1'b0;
      FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_2 <= 1'b0;
      FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_2 <= 1'b0;
      FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_2 <= 1'b0;
    end
    else if ( FpFloatToInt_16U_5U_10U_internal_int_and_cse ) begin
      FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_2 <= MUX1HOT_s_1_3_2(FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_mx0w0,
          FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_9_4_1, (readslicef_11_1_10((cvt_10_IntSaturation_17U_8U_if_acc_2_nl))),
          {and_dcpl_407 , and_dcpl_409 , and_dcpl_411});
      FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_2 <= MUX1HOT_s_1_3_2(FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_mx0w0,
          FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_9_4_1, (readslicef_11_1_10((cvt_2_IntSaturation_17U_8U_if_acc_1_nl))),
          {and_dcpl_407 , and_dcpl_409 , and_dcpl_411});
      FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_2 <= MUX1HOT_s_1_3_2(FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_mx0w0,
          FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_9_4_1, cvt_3_IntSaturation_17U_8U_if_acc_1_itm_10_1,
          {and_dcpl_407 , and_dcpl_409 , and_dcpl_411});
      FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_2 <= MUX1HOT_s_1_3_2(FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_mx0w0,
          FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_9_4_1, (readslicef_11_1_10((cvt_4_IntSaturation_17U_8U_if_acc_2_nl))),
          {and_dcpl_407 , and_dcpl_409 , and_dcpl_411});
      FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_2 <= MUX1HOT_s_1_3_2(FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_mx0w0,
          FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_9_4_1, cvt_5_IntSaturation_17U_8U_if_acc_1_itm_10_1,
          {and_dcpl_407 , and_dcpl_409 , and_dcpl_411});
      FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_2 <= MUX1HOT_s_1_3_2(FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_mx0w0,
          FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_9_4_1, (readslicef_11_1_10((cvt_6_IntSaturation_17U_8U_if_acc_2_nl))),
          {and_dcpl_407 , and_dcpl_409 , and_dcpl_411});
      FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_2 <= MUX1HOT_s_1_3_2(FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_mx0w0,
          FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_9_4_1, cvt_1_IntSaturation_17U_8U_if_acc_itm_10_1,
          {and_dcpl_407 , and_dcpl_409 , and_dcpl_411});
      FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_2 <= MUX1HOT_s_1_3_2(FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_mx0w0,
          FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_9_4_1, (readslicef_11_1_10((cvt_7_IntSaturation_17U_8U_if_acc_2_nl))),
          {and_dcpl_407 , and_dcpl_409 , and_dcpl_411});
      FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_2 <= MUX1HOT_s_1_3_2(FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_mx0w0,
          FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_9_4_1, (readslicef_11_1_10((cvt_16_IntSaturation_17U_8U_if_acc_4_nl))),
          {and_dcpl_407 , and_dcpl_409 , and_dcpl_411});
      FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_2 <= MUX1HOT_s_1_3_2(FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_mx0w0,
          FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_9_4_1, (readslicef_11_1_10((cvt_8_IntSaturation_17U_8U_if_acc_3_nl))),
          {and_dcpl_407 , and_dcpl_409 , and_dcpl_411});
      FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_2 <= MUX1HOT_s_1_3_2(FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_mx0w0,
          FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_9_4_1, (readslicef_11_1_10((cvt_15_IntSaturation_17U_8U_if_acc_3_nl))),
          {and_dcpl_407 , and_dcpl_409 , and_dcpl_411});
      FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_2 <= MUX1HOT_s_1_3_2(FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_mx0w0,
          FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_9_4_1, cvt_9_IntSaturation_17U_8U_if_acc_1_itm_10_1,
          {and_dcpl_407 , and_dcpl_409 , and_dcpl_411});
      FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_2 <= MUX1HOT_s_1_3_2(FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_mx0w0,
          FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_9_4_1, (readslicef_11_1_10((cvt_13_IntSaturation_17U_8U_if_acc_2_nl))),
          {and_dcpl_407 , and_dcpl_409 , and_dcpl_411});
      FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_2 <= MUX1HOT_s_1_3_2(FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_mx0w0,
          FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_9_4_1, (readslicef_11_1_10((cvt_11_IntSaturation_17U_8U_if_acc_2_nl))),
          {and_dcpl_407 , and_dcpl_409 , and_dcpl_411});
      FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_2 <= MUX1HOT_s_1_3_2(FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_mx0w0,
          FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_9_4_1, (readslicef_11_1_10((cvt_12_IntSaturation_17U_8U_if_acc_3_nl))),
          {and_dcpl_407 , and_dcpl_409 , and_dcpl_411});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_1_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (and_896_rgt | and_900_rgt | and_dcpl_420) & (mux_811_nl)
        ) begin
      cvt_1_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_itm_2
          <= MUX1HOT_s_1_3_2((FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_1_sva[0]),
          (FpFloatToInt_16U_5U_10U_if_qr_1_lpi_1_dfm_mx0[0]), IntSaturation_17U_16U_IntSaturation_17U_16U_or_4_itm_2,
          {and_896_rgt , and_900_rgt , and_dcpl_420});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_idata_data_sva_3_47_31_1 <= 17'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_815_nl) ) begin
      chn_idata_data_sva_3_47_31_1 <= chn_idata_data_sva_2_47_31_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_1_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_svs_2
          <= 1'b0;
      cvt_2_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2
          <= 1'b0;
      cvt_3_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2
          <= 1'b0;
      cvt_4_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2
          <= 1'b0;
      cvt_5_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2
          <= 1'b0;
      cvt_16_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_4_svs_2
          <= 1'b0;
      cvt_6_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2
          <= 1'b0;
      cvt_15_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2
          <= 1'b0;
      cvt_7_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2
          <= 1'b0;
      cvt_14_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2
          <= 1'b0;
      cvt_8_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2
          <= 1'b0;
      cvt_13_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2
          <= 1'b0;
      cvt_9_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2
          <= 1'b0;
      cvt_12_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2
          <= 1'b0;
      cvt_10_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2
          <= 1'b0;
      cvt_11_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2
          <= 1'b0;
    end
    else if ( FpFloatToInt_16U_5U_10U_if_and_cse ) begin
      cvt_1_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_svs_2
          <= cvt_1_FpFloatToInt_16U_5U_10U_if_acc_itm_11_1;
      cvt_2_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2
          <= cvt_2_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1;
      cvt_3_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2
          <= cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1;
      cvt_4_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2
          <= cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1;
      cvt_5_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2
          <= cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1;
      cvt_16_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_4_svs_2
          <= cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_itm_11_1;
      cvt_6_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2
          <= cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1;
      cvt_15_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2
          <= cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1;
      cvt_7_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2
          <= cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1;
      cvt_14_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2
          <= cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1;
      cvt_8_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2
          <= cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1;
      cvt_13_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2
          <= cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1;
      cvt_9_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2
          <= cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1;
      cvt_12_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2
          <= cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1;
      cvt_10_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2
          <= cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1;
      cvt_11_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2
          <= cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_5U_10U_land_1_lpi_1_dfm_3 <= 1'b0;
      IsNaN_5U_10U_land_15_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( IsNaN_5U_10U_aelse_and_cse ) begin
      IsNaN_5U_10U_land_1_lpi_1_dfm_3 <= MUX_s_1_2_2(IsNaN_5U_10U_land_1_lpi_1_dfm_mx0w0,
          cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2,
          and_dcpl_424);
      IsNaN_5U_10U_land_15_lpi_1_dfm_3 <= MUX_s_1_2_2(IsNaN_5U_10U_land_15_lpi_1_dfm_mx0w0,
          cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_svs_2,
          and_dcpl_424);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1
          <= 1'b0;
    end
    else if ( core_wen & (cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c0
        | cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c1
        | and_dcpl_420) ) begin
      cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1
          <= MUX1HOT_s_1_3_2((FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_2_sva[0]),
          (FpFloatToInt_16U_5U_10U_if_qr_2_lpi_1_dfm_mx0[0]), IntSaturation_17U_16U_IntSaturation_17U_16U_or_5_itm_2,
          {cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c0
          , cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c1
          , and_dcpl_420});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_idata_data_sva_3_79_63_1 <= 17'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_822_nl) ) begin
      chn_idata_data_sva_3_79_63_1 <= chn_idata_data_sva_2_79_63_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_5U_10U_land_2_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( core_wen & IsNaN_5U_10U_aelse_or_cse & (mux_829_nl) ) begin
      IsNaN_5U_10U_land_2_lpi_1_dfm_4 <= MUX_s_1_2_2(IsNaN_5U_10U_land_2_lpi_1_dfm_mx0w0,
          IsNaN_5U_10U_IsNaN_5U_10U_nand_1_itm_2, and_dcpl_424);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_reg <= 5'b0;
    end
    else if ( (mux_2224_nl) & or_5189_cse & core_wen ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_1_rgt[14:10];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_1_reg <= 10'b0;
    end
    else if ( (((cfg_out_precision_1_sva_st_113==2'b10) & or_4714_cse) | and_2360_cse
        | cvt_unequal_tmp_20) & or_5189_cse & core_wen ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_1_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_1_rgt[9:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1
          <= 1'b0;
    end
    else if ( core_wen & (cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c0
        | cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c1
        | and_dcpl_420) ) begin
      cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1
          <= MUX1HOT_s_1_3_2((FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_3_sva[0]),
          (FpFloatToInt_16U_5U_10U_if_qr_3_lpi_1_dfm_mx0[0]), IntSaturation_17U_16U_IntSaturation_17U_16U_or_6_itm_2,
          {cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c0
          , cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c1
          , and_dcpl_420});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_idata_data_sva_3_111_95_1 <= 17'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_833_nl) ) begin
      chn_idata_data_sva_3_111_95_1 <= chn_idata_data_sva_2_111_95_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_5U_10U_land_3_lpi_1_dfm_5 <= 1'b0;
      IsNaN_5U_10U_land_4_lpi_1_dfm_5 <= 1'b0;
      IsNaN_5U_10U_land_5_lpi_1_dfm_5 <= 1'b0;
      IsNaN_5U_10U_land_lpi_1_dfm_5 <= 1'b0;
      IsNaN_5U_10U_land_6_lpi_1_dfm_5 <= 1'b0;
      IsNaN_5U_10U_land_8_lpi_1_dfm_5 <= 1'b0;
      IsNaN_5U_10U_land_13_lpi_1_dfm_5 <= 1'b0;
      IsNaN_5U_10U_land_9_lpi_1_dfm_5 <= 1'b0;
      IsNaN_5U_10U_land_12_lpi_1_dfm_5 <= 1'b0;
      IsNaN_5U_10U_land_10_lpi_1_dfm_5 <= 1'b0;
      IsNaN_5U_10U_land_11_lpi_1_dfm_5 <= 1'b0;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_1_itm_3 <= 1'b0;
      FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_7_itm_1 <= 10'b0;
    end
    else if ( IsNaN_5U_10U_aelse_and_1_cse ) begin
      IsNaN_5U_10U_land_3_lpi_1_dfm_5 <= MUX_s_1_2_2(IsNaN_5U_10U_land_3_lpi_1_dfm_4,
          cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2, and_dcpl_420);
      IsNaN_5U_10U_land_4_lpi_1_dfm_5 <= MUX_s_1_2_2(IsNaN_5U_10U_land_4_lpi_1_dfm_4,
          cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2, and_dcpl_420);
      IsNaN_5U_10U_land_5_lpi_1_dfm_5 <= MUX_s_1_2_2(IsNaN_5U_10U_land_5_lpi_1_dfm_4,
          cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2, and_dcpl_420);
      IsNaN_5U_10U_land_lpi_1_dfm_5 <= MUX_s_1_2_2(IsNaN_5U_10U_land_lpi_1_dfm_4,
          cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2, and_dcpl_420);
      IsNaN_5U_10U_land_6_lpi_1_dfm_5 <= MUX_s_1_2_2(IsNaN_5U_10U_land_6_lpi_1_dfm_4,
          cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2, and_dcpl_420);
      IsNaN_5U_10U_land_8_lpi_1_dfm_5 <= MUX_s_1_2_2(IsNaN_5U_10U_land_8_lpi_1_dfm_4,
          cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2, and_dcpl_420);
      IsNaN_5U_10U_land_13_lpi_1_dfm_5 <= MUX_s_1_2_2(IsNaN_5U_10U_land_13_lpi_1_dfm_4,
          cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2,
          and_dcpl_420);
      IsNaN_5U_10U_land_9_lpi_1_dfm_5 <= MUX_s_1_2_2(IsNaN_5U_10U_land_9_lpi_1_dfm_4,
          cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2, and_dcpl_420);
      IsNaN_5U_10U_land_12_lpi_1_dfm_5 <= MUX_s_1_2_2(IsNaN_5U_10U_land_12_lpi_1_dfm_4,
          cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2,
          and_dcpl_420);
      IsNaN_5U_10U_land_10_lpi_1_dfm_5 <= MUX_s_1_2_2(IsNaN_5U_10U_land_10_lpi_1_dfm_4,
          cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2,
          and_dcpl_420);
      IsNaN_5U_10U_land_11_lpi_1_dfm_5 <= MUX_s_1_2_2(IsNaN_5U_10U_land_11_lpi_1_dfm_4,
          cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2,
          and_dcpl_420);
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_1_itm_3 <= MUX_s_1_2_2(IntSaturation_17U_16U_IntSaturation_17U_16U_or_1_itm_2,
          chn_idata_data_sva_2_511_1, and_dcpl_408);
      FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_7_itm_1 <= MUX_v_10_2_2((FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_7_nl),
          FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_9_lpi_1_dfm_8, and_dcpl_408);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_reg <= 5'b0;
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_reg <= 5'b0;
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_reg <= 5'b0;
    end
    else if ( and_2365_cse ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_2_rgt[14:10];
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_5_rgt[14:10];
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_13_rgt[14:10];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_1_reg <= 10'b0;
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_1_reg <= 10'b0;
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_1_reg <= 10'b0;
    end
    else if ( and_2369_cse ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_1_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_2_rgt[9:0];
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_1_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_5_rgt[9:0];
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_1_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_13_rgt[9:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1
          <= 1'b0;
    end
    else if ( core_wen & (cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0
        | cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1
        | and_dcpl_420) ) begin
      cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1
          <= MUX1HOT_s_1_3_2((FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_4_sva[0]),
          (FpFloatToInt_16U_5U_10U_if_qr_4_lpi_1_dfm_mx0[0]), IntSaturation_17U_16U_IntSaturation_17U_16U_or_7_itm_2,
          {cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0
          , cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1
          , and_dcpl_420});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_idata_data_sva_3_143_127_1 <= 17'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_837_nl) ) begin
      chn_idata_data_sva_3_143_127_1 <= chn_idata_data_sva_2_143_127_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5 <= 15'b0;
    end
    else if ( core_wen & (and_dcpl_408 | FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c1
        | FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c2) ) begin
      FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5 <= MUX1HOT_v_15_6_2((FpFloatToInt_16U_5U_10U_internal_int_24_1_4_sva[14:0]),
          (FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_4_sva[15:1]), (FpFloatToInt_16U_5U_10U_if_qr_4_lpi_1_dfm_mx0[15:1]),
          15'b100000000000000, IntSaturation_17U_16U_o_15_1_4_lpi_1_dfm_7, IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_2,
          {(FpFloatToInt_16U_5U_10U_and_37_nl) , (FpFloatToInt_16U_5U_10U_and_38_nl)
          , (FpFloatToInt_16U_5U_10U_and_7_nl) , (FpFloatToInt_16U_5U_10U_o_int_and_28_nl)
          , FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c1 , FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5_mx0c2});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_reg <= 5'b0;
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_reg <= 5'b0;
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_reg <= 5'b0;
    end
    else if ( and_2372_cse ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_4_rgt[14:10];
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_14_rgt[14:10];
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_15_rgt[14:10];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_1_reg <= 10'b0;
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_1_reg <= 10'b0;
    end
    else if ( and_2380_cse ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_1_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_4_rgt[9:0];
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_1_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_11_rgt[9:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_idata_data_sva_3_495_479_1 <= 17'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_841_nl) ) begin
      chn_idata_data_sva_3_495_479_1 <= chn_idata_data_sva_2_495_479_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_5_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (and_954_rgt | and_956_rgt | and_dcpl_420) & (mux_849_nl)
        ) begin
      cvt_5_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_2
          <= MUX1HOT_s_1_3_2((FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_5_sva[0]),
          (FpFloatToInt_16U_5U_10U_if_qr_5_lpi_1_dfm_mx0[0]), IntSaturation_17U_16U_IntSaturation_17U_16U_or_8_itm_2,
          {and_954_rgt , and_956_rgt , and_dcpl_420});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_idata_data_sva_3_175_159_1 <= 17'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_853_nl) ) begin
      chn_idata_data_sva_3_175_159_1 <= chn_idata_data_sva_2_175_159_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpFloatToInt_16U_5U_10U_internal_int_0_sva_3 <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_407 | and_957_rgt) & (mux_859_nl) ) begin
      FpFloatToInt_16U_5U_10U_internal_int_0_sva_3 <= MUX_s_1_2_2(FpFloatToInt_16U_5U_10U_internal_int_0_sva_mx0w0,
          FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_9_4_1, and_957_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1
          <= 1'b0;
    end
    else if ( core_wen & (cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1_mx0c0
        | cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1_mx0c1
        | and_dcpl_420) ) begin
      cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1
          <= MUX1HOT_s_1_3_2((FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_sva[0]),
          (FpFloatToInt_16U_5U_10U_if_qr_lpi_1_dfm_mx0[0]), IntSaturation_17U_16U_IntSaturation_17U_16U_or_3_itm_2,
          {cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1_mx0c0
          , cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1_mx0c1
          , and_dcpl_420});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_reg <= 5'b0;
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_reg <= 5'b0;
    end
    else if ( and_2389_cse ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_6_rgt[14:10];
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_12_rgt[14:10];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_1_reg <= 10'b0;
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_1_reg <= 10'b0;
    end
    else if ( and_2393_cse ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_1_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_6_rgt[9:0];
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_1_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_12_rgt[9:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_idata_data_sva_3_463_447_1 <= 17'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_863_nl) ) begin
      chn_idata_data_sva_3_463_447_1 <= chn_idata_data_sva_2_463_447_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1
          <= 1'b0;
    end
    else if ( core_wen & (cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0
        | cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1
        | and_dcpl_420) ) begin
      cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1
          <= MUX1HOT_s_1_3_2((FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_6_sva[0]),
          (FpFloatToInt_16U_5U_10U_if_qr_6_lpi_1_dfm_mx0[0]), IntSaturation_17U_16U_IntSaturation_17U_16U_or_9_itm_2,
          {cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0
          , cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1
          , and_dcpl_420});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_idata_data_sva_3_207_191_1 <= 17'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_867_nl) ) begin
      chn_idata_data_sva_3_207_191_1 <= chn_idata_data_sva_2_207_191_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_reg <= 5'b0;
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_reg <= 5'b0;
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_reg <= 5'b0;
    end
    else if ( and_2396_cse ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_7_rgt[14:10];
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_9_rgt[14:10];
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_11_rgt[14:10];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_1_reg <= 10'b0;
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_1_reg <= 10'b0;
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_1_reg <= 10'b0;
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_1_reg <= 10'b0;
    end
    else if ( and_2402_cse ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_1_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_7_rgt[9:0];
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_1_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_9_rgt[9:0];
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_1_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_14_rgt[9:0];
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_1_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_15_rgt[9:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_15_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (and_984_rgt | and_986_rgt | and_dcpl_420) & (mux_875_nl)
        ) begin
      cvt_15_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_2
          <= MUX1HOT_s_1_3_2((FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_15_sva[0]),
          (FpFloatToInt_16U_5U_10U_if_qr_15_lpi_1_dfm_mx0[0]), IntSaturation_17U_16U_IntSaturation_17U_16U_or_2_itm_2,
          {and_984_rgt , and_986_rgt , and_dcpl_420});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_reg <= 5'b0;
    end
    else if ( (((cfg_out_precision_1_sva_st_113==2'b01) & (cfg_proc_precision_1_sva_st_65==2'b10))
        | cvt_unequal_tmp_20) & or_5189_cse & core_wen ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_8_rgt[14:10];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_1_reg <= 10'b0;
    end
    else if ( (((cfg_out_precision_1_sva_st_113==2'b01)) | cvt_unequal_tmp_20 | and_2360_cse)
        & or_5189_cse & core_wen ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_1_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_8_rgt[9:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_idata_data_sva_3_431_415_1 <= 17'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_879_nl) ) begin
      chn_idata_data_sva_3_431_415_1 <= chn_idata_data_sva_2_431_415_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_7_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (and_987_rgt | and_989_rgt | and_dcpl_420) & (mux_887_nl)
        ) begin
      cvt_7_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_2
          <= MUX1HOT_s_1_3_2((FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_7_sva[0]),
          (FpFloatToInt_16U_5U_10U_if_qr_7_lpi_1_dfm_mx0[0]), IntSaturation_17U_16U_IntSaturation_17U_16U_or_itm_2,
          {and_987_rgt , and_989_rgt , and_dcpl_420});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_idata_data_sva_3_239_223_1 <= 17'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_891_nl) ) begin
      chn_idata_data_sva_3_239_223_1 <= chn_idata_data_sva_2_239_223_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_5U_10U_land_7_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & IsNaN_5U_10U_aelse_or_1_cse & (~ (mux_899_nl)) ) begin
      IsNaN_5U_10U_land_7_lpi_1_dfm_6 <= MUX_s_1_2_2(IsNaN_5U_10U_land_7_lpi_1_dfm_5,
          cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2, and_dcpl_420);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1
          <= 1'b0;
    end
    else if ( core_wen & (cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c0
        | cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c1
        | and_dcpl_420) ) begin
      cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1
          <= MUX1HOT_s_1_3_2((FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_14_sva[0]),
          (FpFloatToInt_16U_5U_10U_if_qr_14_lpi_1_dfm_mx0[0]), IntSaturation_17U_16U_IntSaturation_17U_16U_or_15_itm_2,
          {cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c0
          , cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c1
          , and_dcpl_420});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_5U_10U_land_14_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & IsNaN_5U_10U_aelse_or_1_cse & (mux_909_nl) ) begin
      IsNaN_5U_10U_land_14_lpi_1_dfm_6 <= MUX_s_1_2_2(IsNaN_5U_10U_land_14_lpi_1_dfm_5,
          cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2,
          and_dcpl_420);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_reg <= 5'b0;
    end
    else if ( (mux_2237_nl) & or_5189_cse & core_wen ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_10_rgt[14:10];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_1_reg <= 10'b0;
    end
    else if ( ((mux_2239_nl) | and_2360_cse) & or_5189_cse & core_wen ) begin
      reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_1_reg <= FpFloatToInt_16U_5U_10U_o_int_mux1h_10_rgt[9:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_idata_data_sva_3_399_383_1 <= 17'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_913_nl) ) begin
      chn_idata_data_sva_3_399_383_1 <= chn_idata_data_sva_2_399_383_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_8_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_2
          <= 1'b0;
    end
    else if ( core_wen & (and_1009_rgt | and_1011_rgt | and_dcpl_420) & (mux_921_nl)
        ) begin
      cvt_8_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_2
          <= MUX1HOT_s_1_3_2((FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_8_sva[0]),
          (FpFloatToInt_16U_5U_10U_if_qr_8_lpi_1_dfm_mx0[0]), IntShiftRightSat_49U_6U_17U_o_0_1_sva_2,
          {and_1009_rgt , and_1011_rgt , and_dcpl_420});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_idata_data_sva_3_271_255_1 <= 17'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_925_nl) ) begin
      chn_idata_data_sva_3_271_255_1 <= chn_idata_data_sva_2_271_255_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1
          <= 1'b0;
    end
    else if ( core_wen & (cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0
        | cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1
        | and_dcpl_420) ) begin
      cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1
          <= MUX1HOT_s_1_3_2((FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_13_sva[0]),
          (FpFloatToInt_16U_5U_10U_if_qr_13_lpi_1_dfm_mx0[0]), IntSaturation_17U_16U_IntSaturation_17U_16U_or_14_itm_2,
          {cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0
          , cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1
          , and_dcpl_420});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_idata_data_sva_3_367_351_1 <= 17'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_929_nl) ) begin
      chn_idata_data_sva_3_367_351_1 <= chn_idata_data_sva_2_367_351_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1
          <= 1'b0;
    end
    else if ( core_wen & (cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c0
        | cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c1
        | and_dcpl_420) ) begin
      cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1
          <= MUX1HOT_s_1_3_2((FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_9_sva[0]),
          (FpFloatToInt_16U_5U_10U_if_qr_9_lpi_1_dfm_mx0[0]), IntShiftRightSat_49U_6U_17U_o_0_10_sva_2,
          {cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c0
          , cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1_mx0c1
          , and_dcpl_420});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_idata_data_sva_3_303_287_1 <= 17'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_933_nl) ) begin
      chn_idata_data_sva_3_303_287_1 <= chn_idata_data_sva_2_303_287_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1
          <= 1'b0;
    end
    else if ( core_wen & (cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c0
        | cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c1
        | and_dcpl_420) ) begin
      cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1
          <= MUX1HOT_s_1_3_2((FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_12_sva[0]),
          (FpFloatToInt_16U_5U_10U_if_qr_12_lpi_1_dfm_mx0[0]), IntSaturation_17U_16U_IntSaturation_17U_16U_or_12_itm_2,
          {cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c0
          , cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1_mx0c1
          , and_dcpl_420});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_idata_data_sva_3_335_319_1 <= 17'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_937_nl) ) begin
      chn_idata_data_sva_3_335_319_1 <= chn_idata_data_sva_2_335_319_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1
          <= 1'b0;
    end
    else if ( core_wen & (cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0
        | cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1
        | and_dcpl_420) ) begin
      cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1
          <= MUX1HOT_s_1_3_2((FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_10_sva[0]),
          (FpFloatToInt_16U_5U_10U_if_qr_10_lpi_1_dfm_mx0[0]), IntSaturation_17U_16U_IntSaturation_17U_16U_or_10_itm_2,
          {cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0
          , cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1
          , and_dcpl_420});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1
          <= 1'b0;
    end
    else if ( core_wen & (cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0
        | cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1
        | and_dcpl_420) ) begin
      cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1
          <= MUX1HOT_s_1_3_2((FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_11_sva[0]),
          (FpFloatToInt_16U_5U_10U_if_qr_11_lpi_1_dfm_mx0[0]), IntSaturation_17U_16U_IntSaturation_17U_16U_or_11_itm_2,
          {cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c0
          , cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1_mx0c1
          , and_dcpl_420});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_out_precision_1_sva_6 <= 2'b0;
      cvt_16_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= 1'b0;
      cvt_unequal_tmp_21 <= 1'b0;
      cfg_mode_eql_1_sva_6 <= 1'b0;
      cvt_15_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= 1'b0;
      cvt_14_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= 1'b0;
      cvt_13_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= 1'b0;
      cvt_12_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= 1'b0;
      cvt_11_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= 1'b0;
      cvt_10_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= 1'b0;
      cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= 1'b0;
      cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= 1'b0;
      cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= 1'b0;
      cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= 1'b0;
      cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= 1'b0;
      cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= 1'b0;
      cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= 1'b0;
      cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= 1'b0;
      cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= 1'b0;
      cfg_proc_precision_1_sva_st_66 <= 2'b0;
    end
    else if ( cfg_out_precision_and_32_cse ) begin
      cfg_out_precision_1_sva_6 <= cfg_out_precision_1_sva_st_113;
      cvt_16_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= ~((IntShiftRightSat_49U_6U_17U_i_sva_2 == conv_s2s_18_49(cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl))
          | (IntShiftRightSat_49U_6U_17U_oelse_mux_24_nl));
      cvt_unequal_tmp_21 <= cvt_unequal_tmp_20;
      cfg_mode_eql_1_sva_6 <= cfg_mode_eql_1_sva_5;
      cvt_15_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= ~((IntShiftRightSat_49U_6U_17U_i_15_sva_2 == conv_s2s_18_49(cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl))
          | (IntShiftRightSat_49U_6U_17U_oelse_mux_26_nl));
      cvt_14_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= ~((IntShiftRightSat_49U_6U_17U_i_14_sva_2 == conv_s2s_18_49(cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl))
          | (IntShiftRightSat_49U_6U_17U_oelse_mux_22_nl));
      cvt_13_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= ~((IntShiftRightSat_49U_6U_17U_i_13_sva_2 == conv_s2s_18_49(cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl))
          | (IntShiftRightSat_49U_6U_17U_oelse_mux_28_nl));
      cvt_12_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= ~((IntShiftRightSat_49U_6U_17U_i_12_sva_2 == conv_s2s_18_49(cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl))
          | (IntShiftRightSat_49U_6U_17U_oelse_mux_18_nl));
      cvt_11_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= ~((IntShiftRightSat_49U_6U_17U_i_11_sva_2 == conv_s2s_18_49(cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl))
          | (IntShiftRightSat_49U_6U_17U_oelse_mux_20_nl));
      cvt_10_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= ~((IntShiftRightSat_49U_6U_17U_i_10_sva_2 == conv_s2s_18_49(cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl))
          | (IntShiftRightSat_49U_6U_17U_oelse_mux_16_nl));
      cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= ~((IntShiftRightSat_49U_6U_17U_i_9_sva_2 == conv_s2s_18_49(cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl))
          | (IntShiftRightSat_49U_6U_17U_oelse_mux_30_nl));
      cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= ~((IntShiftRightSat_49U_6U_17U_i_8_sva_2 == conv_s2s_18_49(cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl))
          | (IntShiftRightSat_49U_6U_17U_oelse_mux_10_nl));
      cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= ~((IntShiftRightSat_49U_6U_17U_i_7_sva_2 == conv_s2s_18_49(cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl))
          | (IntShiftRightSat_49U_6U_17U_oelse_mux_12_nl));
      cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= ~((IntShiftRightSat_49U_6U_17U_i_6_sva_2 == conv_s2s_18_49(cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl))
          | (IntShiftRightSat_49U_6U_17U_oelse_mux_8_nl));
      cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= ~((IntShiftRightSat_49U_6U_17U_i_5_sva_2 == conv_s2s_18_49(cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl))
          | (IntShiftRightSat_49U_6U_17U_oelse_mux_14_nl));
      cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= ~((IntShiftRightSat_49U_6U_17U_i_4_sva_2 == conv_s2s_18_49(cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl))
          | (IntShiftRightSat_49U_6U_17U_oelse_mux_4_nl));
      cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= ~((IntShiftRightSat_49U_6U_17U_i_3_sva_2 == conv_s2s_18_49(cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl))
          | (IntShiftRightSat_49U_6U_17U_oelse_mux_6_nl));
      cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= ~((IntShiftRightSat_49U_6U_17U_i_2_sva_2 == conv_s2s_18_49(cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl))
          | (IntShiftRightSat_49U_6U_17U_oelse_mux_2_nl));
      cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_if_nor_itm_2
          <= ~((IntShiftRightSat_49U_6U_17U_i_1_sva_2 == conv_s2s_18_49(cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl))
          | (IntShiftRightSat_49U_6U_17U_oelse_mux_32_nl));
      cfg_proc_precision_1_sva_st_66 <= cfg_proc_precision_1_sva_st_65;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_16_1_sva_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_943_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_16_1_sva_4 <= IntShiftRightSat_49U_6U_17U_o_16_1_sva_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_16_2_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_2_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_16_4_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_4_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_16_6_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_6_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_16_7_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_16_8_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_8_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_7_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_16_10_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_16_11_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_16_12_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_12_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_11_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_16_13_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_16_14_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_16_15_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_16_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_15_sva_3 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_13_sva_3 <= 1'b0;
      cvt_14_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_3_svs_1 <=
          1'b0;
    end
    else if ( IntShiftRightSat_49U_6U_17U_o_and_cse ) begin
      IntShiftRightSat_49U_6U_17U_o_16_2_sva_3 <= IntShiftRightSat_49U_6U_17U_o_16_2_sva_2;
      IntShiftRightSat_49U_6U_17U_o_0_2_sva_3 <= IntShiftRightSat_49U_6U_17U_o_0_2_sva_2;
      IntShiftRightSat_49U_6U_17U_o_16_4_sva_3 <= IntShiftRightSat_49U_6U_17U_o_16_4_sva_2;
      IntShiftRightSat_49U_6U_17U_o_0_4_sva_3 <= IntShiftRightSat_49U_6U_17U_o_0_4_sva_2;
      IntShiftRightSat_49U_6U_17U_o_16_6_sva_3 <= IntShiftRightSat_49U_6U_17U_o_16_6_sva_2;
      IntShiftRightSat_49U_6U_17U_o_0_6_sva_3 <= IntShiftRightSat_49U_6U_17U_o_0_6_sva_2;
      IntShiftRightSat_49U_6U_17U_o_16_7_sva_3 <= IntShiftRightSat_49U_6U_17U_o_16_7_sva_2;
      IntShiftRightSat_49U_6U_17U_o_16_8_sva_3 <= IntShiftRightSat_49U_6U_17U_o_16_8_sva_2;
      IntShiftRightSat_49U_6U_17U_o_0_8_sva_3 <= IntShiftRightSat_49U_6U_17U_o_0_8_sva_2;
      IntShiftRightSat_49U_6U_17U_o_0_7_sva_3 <= IntShiftRightSat_49U_6U_17U_o_0_7_sva_2;
      IntShiftRightSat_49U_6U_17U_o_16_10_sva_3 <= IntShiftRightSat_49U_6U_17U_o_16_10_sva_2;
      IntShiftRightSat_49U_6U_17U_o_16_11_sva_3 <= IntShiftRightSat_49U_6U_17U_o_16_11_sva_2;
      IntShiftRightSat_49U_6U_17U_o_16_12_sva_3 <= IntShiftRightSat_49U_6U_17U_o_16_12_sva_2;
      IntShiftRightSat_49U_6U_17U_o_0_12_sva_3 <= IntShiftRightSat_49U_6U_17U_o_0_12_sva_2;
      IntShiftRightSat_49U_6U_17U_o_0_11_sva_3 <= IntShiftRightSat_49U_6U_17U_o_0_11_sva_2;
      IntShiftRightSat_49U_6U_17U_o_16_13_sva_3 <= IntShiftRightSat_49U_6U_17U_o_16_13_sva_2;
      IntShiftRightSat_49U_6U_17U_o_16_14_sva_3 <= IntShiftRightSat_49U_6U_17U_o_16_14_sva_2;
      IntShiftRightSat_49U_6U_17U_o_16_15_sva_3 <= IntShiftRightSat_49U_6U_17U_o_16_15_sva_2;
      IntShiftRightSat_49U_6U_17U_o_16_sva_3 <= IntShiftRightSat_49U_6U_17U_o_16_sva_2;
      IntShiftRightSat_49U_6U_17U_o_0_sva_3 <= IntShiftRightSat_49U_6U_17U_o_0_sva_2;
      IntShiftRightSat_49U_6U_17U_o_0_15_sva_3 <= IntShiftRightSat_49U_6U_17U_o_0_15_sva_2;
      IntShiftRightSat_49U_6U_17U_o_0_13_sva_3 <= IntShiftRightSat_49U_6U_17U_o_0_13_sva_2;
      cvt_14_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_3_svs_1 <=
          readslicef_11_1_10((cvt_14_IntSaturation_17U_8U_if_acc_3_nl));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_else_nor_dfs_2 <= 1'b0;
      cvt_else_equal_tmp_5 <= 1'b0;
    end
    else if ( cvt_else_and_24_cse ) begin
      cvt_else_nor_dfs_2 <= cvt_else_nor_dfs;
      cvt_else_equal_tmp_5 <= cvt_else_equal_tmp_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_else_equal_tmp_9 <= 1'b0;
    end
    else if ( cvt_else_and_cse & (~(or_dcpl_178 | and_dcpl_535 | (~ main_stage_v_3)))
        & (~ (mux_954_nl)) ) begin
      cvt_else_equal_tmp_9 <= cvt_else_equal_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_16_3_sva_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_959_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_16_3_sva_4 <= IntShiftRightSat_49U_6U_17U_o_16_3_sva_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_else_equal_tmp_16 <= 1'b0;
    end
    else if ( cvt_else_and_cse & (~((~ and_tmp_165) | and_dcpl_535 | (~ main_stage_v_3)))
        & (~ (mux_964_nl)) ) begin
      cvt_else_equal_tmp_16 <= cvt_else_equal_tmp_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_16_5_sva_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_982_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_16_5_sva_4 <= IntShiftRightSat_49U_6U_17U_o_16_5_sva_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_cvt_else_nor_dfs_9_cse <= 1'b0;
      cvt_else_equal_tmp_28 <= 1'b0;
    end
    else if ( cvt_else_and_10_cse ) begin
      reg_cvt_else_nor_dfs_9_cse <= cvt_else_nor_dfs;
      cvt_else_equal_tmp_28 <= cvt_else_equal_tmp_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_else_nor_dfs_11 <= 1'b0;
      cvt_else_equal_tmp_34 <= 1'b0;
      cvt_else_equal_tmp_33 <= 1'b0;
    end
    else if ( cvt_else_and_34_cse ) begin
      cvt_else_nor_dfs_11 <= cvt_else_nor_dfs;
      cvt_else_equal_tmp_34 <= cvt_else_equal_tmp_1;
      cvt_else_equal_tmp_33 <= cvt_else_equal_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_else_nor_dfs_10 <= 1'b0;
    end
    else if ( cvt_else_and_cse & reg_cvt_else_cvt_else_nor_4_cse & (~ (mux_995_nl))
        ) begin
      cvt_else_nor_dfs_10 <= cvt_else_nor_dfs;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_else_nor_dfs_15 <= 1'b0;
      cvt_else_equal_tmp_46 <= 1'b0;
      cvt_else_equal_tmp_45 <= 1'b0;
    end
    else if ( cvt_else_and_19_cse ) begin
      cvt_else_nor_dfs_15 <= cvt_else_nor_dfs;
      cvt_else_equal_tmp_46 <= cvt_else_equal_tmp_1;
      cvt_else_equal_tmp_45 <= cvt_else_equal_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_odata_data_13_0_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_195 | or_dcpl_4)) ) begin
      chn_odata_data_13_0_lpi_1_dfm_1 <= chn_odata_data_13_0_lpi_1_dfm_1_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_16_9_sva_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1000_nl) ) begin
      IntShiftRightSat_49U_6U_17U_o_16_9_sva_4 <= IntShiftRightSat_49U_6U_17U_o_16_9_sva_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_0_3_sva_4 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_5_sva_4 <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_0_9_sva_4 <= 1'b0;
    end
    else if ( IntShiftRightSat_49U_6U_17U_o_and_103_cse ) begin
      IntShiftRightSat_49U_6U_17U_o_0_3_sva_4 <= IntShiftRightSat_49U_6U_17U_o_0_3_sva_3;
      IntShiftRightSat_49U_6U_17U_o_0_5_sva_4 <= IntShiftRightSat_49U_6U_17U_o_0_5_sva_3;
      IntShiftRightSat_49U_6U_17U_o_0_9_sva_4 <= IntShiftRightSat_49U_6U_17U_o_0_9_sva_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_is_inf_1_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1004_nl) ) begin
      FpIntToFloat_17U_5U_10U_is_inf_1_lpi_1_dfm_6 <= ~(((~((~ cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_1_itm_4)
          & (FpMantRNE_17U_11U_else_mux_1_nl))) & (FpIntToFloat_17U_5U_10U_else_mux_1_nl))
          | IsNaN_5U_10U_IsNaN_5U_10U_nand_1_itm_2);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_1_lpi_1_dfm_7_itm <= 1'b0;
    end
    else if ( (mux_2250_nl) & or_4862_cse & core_wen & (~ cfg_mode_eql_1_sva_5) &
        main_stage_v_2 & (cfg_out_precision_1_sva_st_113==2'b10) & (~ IsNaN_5U_10U_IsNaN_5U_10U_nand_1_itm_2)
        & (~ cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_svs_st_2)
        & or_5189_cse & cvt_unequal_tmp_20 ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_1_lpi_1_dfm_7_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_1_itm[4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_1_lpi_1_dfm_7_1_itm <= 4'b0;
    end
    else if ( (mux_2251_nl) & core_wen & (~ cfg_mode_eql_1_sva_5) & main_stage_v_2
        & or_5189_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_1_lpi_1_dfm_7_1_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_1_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_1_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_svs_st_2 <=
          1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1011_nl) ) begin
      cvt_1_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_svs_st_2 <=
          cvt_1_IntSaturation_17U_8U_if_acc_itm_10_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_is_inf_2_lpi_1_dfm_6 <= 1'b0;
    end
    else if ( cvt_else_and_cse & ((and_tmp_50 & and_dcpl_401) | and_1077_rgt) & (~
        (mux_1018_nl)) ) begin
      FpIntToFloat_17U_5U_10U_is_inf_2_lpi_1_dfm_6 <= MUX_s_1_2_2((FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_nor_1_nl),
          cvt_else_equal_tmp, and_1077_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_2_lpi_1_dfm_8_itm <= 1'b0;
    end
    else if ( (mux_2252_nl) & or_4714_cse & or_4862_cse & core_wen & (~ cfg_mode_eql_1_sva_5)
        & main_stage_v_2 & (cfg_out_precision_1_sva_st_113==2'b10) & (~ cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2)
        & (~ cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2)
        & (cfg_out_precision_1_sva_st_149==2'b10) & or_5189_cse & cvt_unequal_tmp_20
        ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_2_lpi_1_dfm_8_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_3_itm[4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_2_lpi_1_dfm_8_1_itm <= 4'b0;
    end
    else if ( (mux_2253_nl) & (~ cfg_mode_eql_1_sva_5) & main_stage_v_2 & core_wen
        & or_5189_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_2_lpi_1_dfm_8_1_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_3_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_is_inf_3_lpi_1_dfm_7 <= 1'b0;
      FpIntToFloat_17U_5U_10U_is_inf_5_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( FpIntToFloat_17U_5U_10U_is_inf_and_14_cse ) begin
      FpIntToFloat_17U_5U_10U_is_inf_3_lpi_1_dfm_7 <= ~(((~((~ cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4)
          & (FpMantRNE_17U_11U_else_mux_5_nl))) & (FpIntToFloat_17U_5U_10U_else_mux_7_nl))
          | cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2);
      FpIntToFloat_17U_5U_10U_is_inf_5_lpi_1_dfm_7 <= ~(((~((~ cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4)
          & (FpMantRNE_17U_11U_else_mux_9_nl))) & (FpIntToFloat_17U_5U_10U_else_mux_13_nl))
          | cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_3_lpi_1_dfm_8_itm <= 1'b0;
    end
    else if ( (mux_2254_nl) & or_4714_cse & or_4862_cse & core_wen & (~ cfg_mode_eql_1_sva_5)
        & main_stage_v_2 & (cfg_out_precision_1_sva_st_113==2'b10) & (~ cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2)
        & (~ cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2)
        & (cfg_out_precision_1_sva_st_149==2'b10) & or_5189_cse & cvt_unequal_tmp_20
        ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_3_lpi_1_dfm_8_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_5_itm[4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_3_lpi_1_dfm_8_1_itm <= 4'b0;
    end
    else if ( (mux_2255_nl) & (~ cfg_mode_eql_1_sva_5) & main_stage_v_2 & core_wen
        & or_5189_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_3_lpi_1_dfm_8_1_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_5_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_3_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1035_nl) ) begin
      cvt_3_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2
          <= cvt_3_IntSaturation_17U_8U_if_acc_1_itm_10_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( cvt_else_and_cse & ((mux_tmp_321 & and_dcpl_401) | and_1091_rgt) &
        (~ (mux_1054_nl)) ) begin
      FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_7 <= MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_2_mx1w0,
          cvt_else_equal_tmp_1, and_1091_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_4_lpi_1_dfm_9_itm <= 1'b0;
    end
    else if ( cvt_unequal_tmp_20 & (mux_2256_nl) & or_400_cse_1 & or_4714_cse & or_4862_cse
        & core_wen & (~ cfg_mode_eql_1_sva_5) & main_stage_v_2 & (cfg_out_precision_1_sva_st_113==2'b10)
        & (~ cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2)
        & (~ FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_3) & (cfg_out_precision_1_sva_st_149==2'b10)
        & or_5189_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_4_lpi_1_dfm_9_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_7_itm[4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_4_lpi_1_dfm_9_1_itm <= 4'b0;
    end
    else if ( (mux_2257_nl) & and_dcpl_1319 & (~ cfg_mode_eql_1_sva_5) & or_5189_cse
        ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_4_lpi_1_dfm_9_1_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_7_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_5_lpi_1_dfm_8_itm <= 1'b0;
    end
    else if ( (mux_2258_nl) & or_4714_cse & or_4862_cse & core_wen & (~ cfg_mode_eql_1_sva_5)
        & main_stage_v_2 & (cfg_out_precision_1_sva_st_113==2'b10) & (~ cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2)
        & (~ cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2)
        & (cfg_out_precision_1_sva_st_149==2'b10) & or_5189_cse & cvt_unequal_tmp_20
        ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_5_lpi_1_dfm_8_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_9_itm[4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_5_lpi_1_dfm_8_1_itm <= 4'b0;
    end
    else if ( (mux_2259_nl) & (~ cfg_mode_eql_1_sva_5) & main_stage_v_2 & core_wen
        & or_5189_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_5_lpi_1_dfm_8_1_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_9_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_5_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1070_nl) ) begin
      cvt_5_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2
          <= cvt_5_IntSaturation_17U_8U_if_acc_1_itm_10_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( cvt_else_and_cse & FpIntToFloat_17U_5U_10U_is_inf_FpIntToFloat_17U_5U_10U_is_inf_or_15_cse
        & (~ (mux_1077_nl)) ) begin
      FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_7 <= MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_2_mx1w0,
          cvt_else_equal_tmp, and_1104_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_6_lpi_1_dfm_9_itm <= 1'b0;
    end
    else if ( cvt_unequal_tmp_20 & (mux_2260_nl) & or_400_cse_1 & or_4714_cse & or_4862_cse
        & core_wen & (~ cfg_mode_eql_1_sva_5) & main_stage_v_2 & (cfg_out_precision_1_sva_st_113==2'b10)
        & (~ cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2)
        & (~ FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_3) & (cfg_out_precision_1_sva_st_149==2'b10)
        & or_5189_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_6_lpi_1_dfm_9_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_11_itm[4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_6_lpi_1_dfm_9_1_itm <= 4'b0;
    end
    else if ( (mux_2261_nl) & main_stage_v_2 & (~ cfg_mode_eql_1_sva_5) & core_wen
        & or_5189_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_6_lpi_1_dfm_9_1_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_11_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( cvt_else_and_cse & FpIntToFloat_17U_5U_10U_is_inf_FpIntToFloat_17U_5U_10U_is_inf_or_15_cse
        & (~ (mux_1091_nl)) ) begin
      FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_7 <= MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_2_mx1w0,
          cvt_else_equal_tmp, and_1104_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_7_lpi_1_dfm_9_itm <= 1'b0;
    end
    else if ( cvt_unequal_tmp_20 & (mux_2262_nl) & or_400_cse_1 & or_4714_cse & or_4862_cse
        & core_wen & (~ cfg_mode_eql_1_sva_5) & main_stage_v_2 & (cfg_out_precision_1_sva_st_113==2'b10)
        & (~ cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2)
        & (~ FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_3) & (cfg_out_precision_1_sva_st_149==2'b10)
        & or_5189_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_7_lpi_1_dfm_9_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_13_itm[4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_7_lpi_1_dfm_9_1_itm <= 4'b0;
    end
    else if ( (mux_2263_nl) & main_stage_v_2 & (~ cfg_mode_eql_1_sva_5) & core_wen
        & or_5189_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_7_lpi_1_dfm_9_1_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_13_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( cvt_else_and_cse & FpIntToFloat_17U_5U_10U_is_inf_FpIntToFloat_17U_5U_10U_is_inf_or_15_cse
        & (~ (mux_1116_nl)) ) begin
      FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_8 <= MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_2_mx1w0,
          cvt_else_equal_tmp_1, and_1104_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_8_lpi_1_dfm_10_itm <= 1'b0;
    end
    else if ( cvt_unequal_tmp_20 & (mux_2264_nl) & or_400_cse_1 & or_4714_cse & or_4862_cse
        & core_wen & (~ cfg_mode_eql_1_sva_5) & main_stage_v_2 & (cfg_out_precision_1_sva_st_113==2'b10)
        & (~ cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2)
        & (~ FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_3) & (cfg_out_precision_1_sva_st_149==2'b10)
        & or_5189_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_8_lpi_1_dfm_10_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_15_itm[4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_8_lpi_1_dfm_10_1_itm <= 4'b0;
    end
    else if ( (mux_2265_nl) & (~ cfg_mode_eql_1_sva_5) & core_wen & main_stage_v_2
        & or_5189_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_8_lpi_1_dfm_10_1_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_15_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_is_inf_9_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1127_nl) ) begin
      FpIntToFloat_17U_5U_10U_is_inf_9_lpi_1_dfm_7 <= ~(((~((~ cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4)
          & (FpMantRNE_17U_11U_else_mux_17_nl))) & (FpIntToFloat_17U_5U_10U_else_mux_25_nl))
          | cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_9_lpi_1_dfm_8_itm <= 1'b0;
    end
    else if ( (mux_2266_nl) & or_4714_cse & or_4862_cse & core_wen & (~ cfg_mode_eql_1_sva_5)
        & main_stage_v_2 & (cfg_out_precision_1_sva_st_113==2'b10) & (~ cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2)
        & (~ cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2)
        & (cfg_out_precision_1_sva_st_149==2'b10) & or_5189_cse & cvt_unequal_tmp_20
        ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_9_lpi_1_dfm_8_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_17_itm[4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_9_lpi_1_dfm_8_1_itm <= 4'b0;
    end
    else if ( (mux_2267_nl) & (~ cfg_mode_eql_1_sva_5) & main_stage_v_2 & core_wen
        & or_5189_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_9_lpi_1_dfm_8_1_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_17_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_9_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2
          <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1134_nl) ) begin
      cvt_9_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2
          <= cvt_9_IntSaturation_17U_8U_if_acc_1_itm_10_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( core_wen & FpIntToFloat_17U_5U_10U_is_inf_or_cse ) begin
      FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_7 <= MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_2_mx0w0,
          cvt_else_equal_tmp, and_dcpl_617);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_10_lpi_1_dfm_9_itm <= 1'b0;
    end
    else if ( cvt_unequal_tmp_20 & (mux_2268_nl) & or_400_cse_1 & or_4714_cse & or_4862_cse
        & core_wen & (~ cfg_mode_eql_1_sva_5) & main_stage_v_2 & (cfg_out_precision_1_sva_st_113==2'b10)
        & (~ cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2)
        & (~ FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_3) & (cfg_out_precision_1_sva_st_149==2'b10)
        & or_5189_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_10_lpi_1_dfm_9_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_19_itm[4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_10_lpi_1_dfm_9_1_itm <= 4'b0;
    end
    else if ( (mux_2269_nl) & main_stage_v_2 & (~ cfg_mode_eql_1_sva_5) & core_wen
        & or_5189_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_10_lpi_1_dfm_9_1_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_19_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_7 <= 1'b0;
    end
    else if ( cvt_else_and_cse & FpIntToFloat_17U_5U_10U_is_inf_or_cse & (~ (mux_1163_nl))
        ) begin
      FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_7 <= MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_2_mx1w0,
          cvt_else_equal_tmp, and_dcpl_617);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_11_lpi_1_dfm_9_itm <= 1'b0;
    end
    else if ( cvt_unequal_tmp_20 & (mux_2270_nl) & or_4714_cse & or_400_cse_1 & or_4862_cse
        & core_wen & (~ cfg_mode_eql_1_sva_5) & main_stage_v_2 & (cfg_out_precision_1_sva_st_113==2'b10)
        & (~ cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2)
        & (~ FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_3) & (cfg_out_precision_1_sva_st_149==2'b10)
        & or_5189_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_11_lpi_1_dfm_9_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_21_itm[4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_11_lpi_1_dfm_9_1_itm <= 4'b0;
    end
    else if ( (mux_2271_nl) & main_stage_v_2 & (~ cfg_mode_eql_1_sva_5) & core_wen
        & or_5189_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_11_lpi_1_dfm_9_1_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_21_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( cvt_else_and_cse & FpIntToFloat_17U_5U_10U_is_inf_or_cse & (~ (mux_1179_nl))
        ) begin
      FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_8 <= MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_2_mx1w0,
          cvt_else_equal_tmp_1, and_dcpl_617);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_12_lpi_1_dfm_10_itm <= 1'b0;
    end
    else if ( cvt_unequal_tmp_20 & (mux_2272_nl) & or_4714_cse & or_400_cse_1 & or_4862_cse
        & core_wen & (~ cfg_mode_eql_1_sva_5) & main_stage_v_2 & (cfg_out_precision_1_sva_st_113==2'b10)
        & (~ cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2)
        & (~ FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_3) & (cfg_out_precision_1_sva_st_149==2'b10)
        & or_5189_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_12_lpi_1_dfm_10_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_23_itm[4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_12_lpi_1_dfm_10_1_itm <= 4'b0;
    end
    else if ( (mux_2273_nl) & main_stage_v_2 & (~ cfg_mode_eql_1_sva_5) & core_wen
        & or_5189_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_12_lpi_1_dfm_10_1_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_23_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_7 <= 1'b0;
      FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_8 <= 1'b0;
    end
    else if ( FpIntToFloat_17U_5U_10U_is_inf_and_8_cse ) begin
      FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_7 <= MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_2_mx0w0,
          cvt_else_equal_tmp, and_dcpl_631);
      FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_8 <= MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2_mx0w0,
          cvt_else_equal_tmp_1, and_dcpl_631);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_13_lpi_1_dfm_9_itm <= 1'b0;
    end
    else if ( cvt_unequal_tmp_20 & (mux_2274_nl) & or_4714_cse & or_400_cse_1 & or_4862_cse
        & core_wen & (~ cfg_mode_eql_1_sva_5) & main_stage_v_2 & (cfg_out_precision_1_sva_st_113==2'b10)
        & (~ cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2)
        & (~ FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_3) & (cfg_out_precision_1_sva_st_149==2'b10)
        & or_5189_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_13_lpi_1_dfm_9_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_25_itm[4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_13_lpi_1_dfm_9_1_itm <= 4'b0;
    end
    else if ( (mux_2275_nl) & main_stage_v_2 & (~ cfg_mode_eql_1_sva_5) & core_wen
        & or_5189_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_13_lpi_1_dfm_9_1_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_25_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_0_14_sva_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_1204_nl)) ) begin
      IntShiftRightSat_49U_6U_17U_o_0_14_sva_4 <= IntShiftRightSat_49U_6U_17U_o_0_14_sva_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm_4 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_1213_nl)) ) begin
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm_4 <= IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_14_lpi_1_dfm_10_itm <= 1'b0;
    end
    else if ( cvt_unequal_tmp_20 & (mux_2276_nl) & or_4714_cse & or_400_cse_1 & or_4862_cse
        & core_wen & (~ cfg_mode_eql_1_sva_5) & main_stage_v_2 & (cfg_out_precision_1_sva_st_113==2'b10)
        & (~ cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2)
        & (~ FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2) & (cfg_out_precision_1_sva_st_149==2'b10)
        & or_5189_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_14_lpi_1_dfm_10_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_27_itm[4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_14_lpi_1_dfm_10_1_itm <= 4'b0;
    end
    else if ( (mux_2277_nl) & and_dcpl_1319 & (~ cfg_mode_eql_1_sva_5) & or_5189_cse
        ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_14_lpi_1_dfm_10_1_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_27_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRightSat_49U_6U_17U_o_15_1_14_1_reg <= 5'b0;
    end
    else if ( or_5189_cse & core_wen & (~ (cfg_out_precision_1_sva_st_149[1])) )
        begin
      reg_IntShiftRightSat_49U_6U_17U_o_15_1_14_1_reg <= IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_mux_rgt[14:10];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_IntShiftRightSat_49U_6U_17U_o_15_1_14_3_reg <= 10'b0;
    end
    else if ( or_5189_cse & core_wen ) begin
      reg_IntShiftRightSat_49U_6U_17U_o_15_1_14_3_reg <= IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_mux_rgt[9:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_8 <= 1'b0;
      FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_9 <= 1'b0;
    end
    else if ( FpIntToFloat_17U_5U_10U_is_inf_and_10_cse ) begin
      FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_8 <= MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_2_mx0w0,
          cvt_else_equal_tmp, and_dcpl_648);
      FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_9 <= MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_2_mx0w0,
          cvt_else_equal_tmp_1, and_dcpl_648);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_15_lpi_1_dfm_10_itm <= 1'b0;
    end
    else if ( cvt_unequal_tmp_20 & (mux_2278_nl) & or_4714_cse & or_400_cse_1 & or_4862_cse
        & core_wen & (~ cfg_mode_eql_1_sva_5) & main_stage_v_2 & (cfg_out_precision_1_sva_st_113==2'b10)
        & (~ cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2)
        & (~ FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_3) & (cfg_out_precision_1_sva_st_149==2'b10)
        & or_5189_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_15_lpi_1_dfm_10_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_29_itm[4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_15_lpi_1_dfm_10_1_itm <= 4'b0;
    end
    else if ( (mux_2279_nl) & and_dcpl_1319 & (~ cfg_mode_eql_1_sva_5) & or_5189_cse
        ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_15_lpi_1_dfm_10_1_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_29_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_lpi_1_dfm_11_itm <= 1'b0;
    end
    else if ( cvt_unequal_tmp_20 & (mux_2280_nl) & or_4714_cse & or_400_cse_1 & or_4862_cse
        & core_wen & (~ cfg_mode_eql_1_sva_5) & main_stage_v_2 & (cfg_out_precision_1_sva_st_113==2'b10)
        & (~ cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_svs_2)
        & (~ FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_3) & (cfg_out_precision_1_sva_st_149==2'b10)
        & or_5189_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_lpi_1_dfm_11_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_31_itm[4];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_lpi_1_dfm_11_1_itm <= 4'b0;
    end
    else if ( (mux_2281_nl) & (~ cfg_mode_eql_1_sva_5) & core_wen & main_stage_v_2
        & or_5189_cse ) begin
      reg_FpIntToFloat_17U_5U_10U_o_expo_lpi_1_dfm_11_1_itm <= FpIntToFloat_17U_5U_10U_o_expo_mux1h_31_itm[3:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_out_precision_1_sva_st_156 <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1262_nl) ) begin
      cfg_out_precision_1_sva_st_156 <= cfg_out_precision_1_sva_st_149;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_proc_precision_1_sva_st_108 <= 2'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1266_nl) ) begin
      cfg_proc_precision_1_sva_st_108 <= cfg_proc_precision_1_sva_st_101;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_proc_precision_1_sva_st_102 <= 2'b0;
      cfg_out_precision_1_sva_st_144 <= 2'b0;
    end
    else if ( cfg_proc_precision_and_40_cse ) begin
      cfg_proc_precision_1_sva_st_102 <= cfg_proc_precision_1_sva_st_101;
      cfg_out_precision_1_sva_st_144 <= cfg_out_precision_1_sva_st_149;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cfg_proc_precision_1_sva_st_90 <= 2'b0;
      cfg_out_precision_1_sva_st_136 <= 2'b0;
    end
    else if ( cfg_proc_precision_and_43_cse ) begin
      cfg_proc_precision_1_sva_st_90 <= cfg_proc_precision_1_sva_st_89;
      cfg_out_precision_1_sva_st_136 <= cfg_out_precision_1_sva_st_113;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_idata_data_sva_3_15_0_reg <= 1'b0;
    end
    else if ( or_5189_cse & cfg_mode_eql_1_sva_5 & core_wen ) begin
      reg_chn_idata_data_sva_3_15_0_reg <= chn_idata_data_mux1h_65_rgt[15];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_idata_data_sva_3_15_0_1_reg <= 5'b0;
    end
    else if ( ((~((~((cfg_proc_precision_1_sva_st_65!=2'b10) | (cfg_out_precision_1_sva_st_113[0])))
        | (cfg_out_precision_1_sva_st_113[1]))) | cfg_mode_eql_1_sva_5) & or_5189_cse
        & core_wen ) begin
      reg_chn_idata_data_sva_3_15_0_1_reg <= chn_idata_data_mux1h_65_rgt[14:10];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_idata_data_sva_3_15_0_2_reg <= 10'b0;
    end
    else if ( ((~ (mux_2249_nl)) | cfg_mode_eql_1_sva_5) & or_5189_cse & core_wen
        ) begin
      reg_chn_idata_data_sva_3_15_0_2_reg <= chn_idata_data_mux1h_65_rgt[9:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_3 <= 1'b0;
      FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( FpIntToFloat_17U_5U_10U_is_inf_and_23_cse ) begin
      FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_3 <= MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_2_mx1w0,
          cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp, and_1249_cse);
      FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_3 <= MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_2_mx1w0,
          cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp, and_1249_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2 <= 1'b0;
    end
    else if ( cvt_else_and_cse & ((or_tmp_3032 & or_4862_cse & or_4714_cse & or_5189_cse
        & (cfg_out_precision_1_sva_st_149==2'b10) & main_stage_v_2 & or_400_cse_1)
        | and_1213_rgt) & (mux_1429_nl) ) begin
      FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2 <= MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2_mx0w0,
          cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp, and_1213_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_3 <= 1'b0;
      FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( FpIntToFloat_17U_5U_10U_is_inf_and_26_cse ) begin
      FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_3 <= MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_2_mx0w0,
          cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp, and_1249_cse);
      FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_3 <= MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_2_mx0w0,
          cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_tmp, and_1249_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 <= 1'b0;
      cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 <= 1'b0;
      cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 <= 1'b0;
    end
    else if ( FpIntToFloat_17U_5U_10U_if_and_16_cse ) begin
      cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 <= cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp;
      cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 <= cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp;
      cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 <= cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 <= 1'b0;
      cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 <= 1'b0;
      cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 <= 1'b0;
      cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 <= 1'b0;
      cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 <= 1'b0;
    end
    else if ( FpIntToFloat_17U_5U_10U_if_and_18_cse ) begin
      cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 <= MUX_s_1_2_2(cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp,
          cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs, and_1247_rgt);
      cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 <= MUX_s_1_2_2(cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp,
          cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs, and_1247_rgt);
      cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 <= MUX_s_1_2_2(cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp,
          cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs, and_1247_rgt);
      cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 <= MUX_s_1_2_2(cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp,
          cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs, and_1247_rgt);
      cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 <= MUX_s_1_2_2(cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp,
          cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs, and_1247_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 <= 1'b0;
    end
    else if ( core_wen & (and_1249_cse | and_1250_rgt) & (mux_1472_nl) ) begin
      cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 <= MUX_s_1_2_2(cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp,
          cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs, and_1250_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2 <= 1'b0;
      cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2 <= 1'b0;
    end
    else if ( FpIntToFloat_17U_5U_10U_if_and_22_cse ) begin
      cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2 <= MUX_s_1_2_2(cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp,
          cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs, and_1247_rgt);
      cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2 <= MUX_s_1_2_2(cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp,
          cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs, and_1247_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 <= 1'b0;
      cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2 <= 1'b0;
      cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_svs_2 <= 1'b0;
    end
    else if ( FpIntToFloat_17U_5U_10U_if_and_27_cse ) begin
      cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 <= MUX_s_1_2_2(cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp,
          cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs, and_1247_rgt);
      cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2 <= MUX_s_1_2_2(cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp,
          cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs, and_1247_rgt);
      cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_svs_2 <= MUX_s_1_2_2(cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_tmp,
          cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_svs, and_1247_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2 <= 1'b0;
    end
    else if ( core_wen & ((and_tmp_12 & (cfg_out_precision_1_sva_st_154==2'b10) &
        or_5189_cse) | and_1247_rgt) & mux_1521_cse ) begin
      cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2 <= MUX_s_1_2_2(cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp,
          cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs, and_1247_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_16_7_sva <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_15_1_6_sva <= 15'b0;
      IntShiftRightSat_49U_6U_17U_o_16_6_sva <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_15_1_7_sva <= 15'b0;
    end
    else if ( IntShiftRightSat_49U_6U_17U_o_and_107_cse ) begin
      IntShiftRightSat_49U_6U_17U_o_16_7_sva <= IntShiftRightSat_49U_6U_17U_o_16_7_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_15_1_6_sva <= IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_16_6_sva <= IntShiftRightSat_49U_6U_17U_o_16_6_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_15_1_7_sva <= IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_16_8_sva <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_15_1_8_sva <= 15'b0;
    end
    else if ( IntShiftRightSat_49U_6U_17U_o_and_108_cse ) begin
      IntShiftRightSat_49U_6U_17U_o_16_8_sva <= IntShiftRightSat_49U_6U_17U_o_16_8_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_15_1_8_sva <= IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_16_10_sva <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_16_11_sva <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_15_1_2_sva <= 15'b0;
      IntShiftRightSat_49U_6U_17U_o_16_2_sva <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_15_1_3_sva <= 15'b0;
      IntShiftRightSat_49U_6U_17U_o_15_1_9_sva <= 15'b0;
      IntShiftRightSat_49U_6U_17U_o_15_1_10_sva <= 15'b0;
      IntShiftRightSat_49U_6U_17U_o_15_1_11_sva <= 15'b0;
    end
    else if ( IntShiftRightSat_49U_6U_17U_o_and_109_cse ) begin
      IntShiftRightSat_49U_6U_17U_o_16_10_sva <= IntShiftRightSat_49U_6U_17U_o_16_10_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_16_11_sva <= IntShiftRightSat_49U_6U_17U_o_16_11_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_15_1_2_sva <= IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_16_2_sva <= IntShiftRightSat_49U_6U_17U_o_16_2_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_15_1_3_sva <= IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_15_1_9_sva <= IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_15_1_10_sva <= IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_15_1_11_sva <= IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_16_12_sva <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_15_1_12_sva <= 15'b0;
    end
    else if ( IntShiftRightSat_49U_6U_17U_o_and_111_cse ) begin
      IntShiftRightSat_49U_6U_17U_o_16_12_sva <= IntShiftRightSat_49U_6U_17U_o_16_12_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_15_1_12_sva <= IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_16_13_sva <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_16_14_sva <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_15_1_4_sva <= 15'b0;
      IntShiftRightSat_49U_6U_17U_o_16_4_sva <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_15_1_13_sva <= 15'b0;
      IntShiftRightSat_49U_6U_17U_o_15_1_14_sva <= 15'b0;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm <= 1'b0;
    end
    else if ( IntShiftRightSat_49U_6U_17U_o_and_112_cse ) begin
      IntShiftRightSat_49U_6U_17U_o_16_13_sva <= IntShiftRightSat_49U_6U_17U_o_16_13_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_16_14_sva <= IntShiftRightSat_49U_6U_17U_o_16_14_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_15_1_4_sva <= IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_16_4_sva <= IntShiftRightSat_49U_6U_17U_o_16_4_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_15_1_13_sva <= IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_15_1_14_sva <= IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_mx0w0;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm <= IntSaturation_17U_16U_IntSaturation_17U_16U_or_13_itm_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_16_15_sva <= 1'b0;
      IntShiftRightSat_49U_6U_17U_o_15_1_15_sva <= 15'b0;
    end
    else if ( IntShiftRightSat_49U_6U_17U_o_and_114_cse ) begin
      IntShiftRightSat_49U_6U_17U_o_16_15_sva <= IntShiftRightSat_49U_6U_17U_o_16_15_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_15_1_15_sva <= IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_sva <= 15'b0;
      IntShiftRightSat_49U_6U_17U_o_16_sva <= 1'b0;
    end
    else if ( IntShiftRightSat_49U_6U_17U_o_and_115_cse ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_sva <= IntShiftRightSat_49U_6U_17U_o_15_1_sva_mx0w0;
      IntShiftRightSat_49U_6U_17U_o_16_sva <= IntShiftRightSat_49U_6U_17U_o_16_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_idata_data_sva_1_511_1 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_1533_nl)) ) begin
      chn_idata_data_sva_1_511_1 <= chn_in_rsci_d_mxwt[511];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_1_sva_2 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1534_nl) ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_1_sva_2 <= nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_1_sva_2[4:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_24U_11U_else_carry_1_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1535_nl) ) begin
      FpMantRNE_24U_11U_else_carry_1_sva_2 <= FpMantRNE_24U_11U_else_carry_1_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_2_sva_2 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1536_nl) ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_2_sva_2 <= nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_2_sva_2[4:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_24U_11U_else_carry_2_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1537_nl) ) begin
      FpMantRNE_24U_11U_else_carry_2_sva_2 <= FpMantRNE_24U_11U_else_carry_2_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_3_sva_2 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1538_nl) ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_3_sva_2 <= nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_3_sva_2[4:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_24U_11U_else_carry_3_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1539_nl) ) begin
      FpMantRNE_24U_11U_else_carry_3_sva_2 <= FpMantRNE_24U_11U_else_carry_3_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_4_sva_2 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1540_nl) ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_4_sva_2 <= nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_4_sva_2[4:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_24U_11U_else_carry_4_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1541_nl) ) begin
      FpMantRNE_24U_11U_else_carry_4_sva_2 <= FpMantRNE_24U_11U_else_carry_4_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_5_sva_2 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1542_nl) ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_5_sva_2 <= nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_5_sva_2[4:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_24U_11U_else_carry_5_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1543_nl) ) begin
      FpMantRNE_24U_11U_else_carry_5_sva_2 <= FpMantRNE_24U_11U_else_carry_5_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_6_sva_2 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1544_nl) ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_6_sva_2 <= nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_6_sva_2[4:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_24U_11U_else_carry_6_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1545_nl) ) begin
      FpMantRNE_24U_11U_else_carry_6_sva_2 <= FpMantRNE_24U_11U_else_carry_6_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_7_sva_2 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1546_nl) ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_7_sva_2 <= nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_7_sva_2[4:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_24U_11U_else_carry_7_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1547_nl) ) begin
      FpMantRNE_24U_11U_else_carry_7_sva_2 <= FpMantRNE_24U_11U_else_carry_7_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_8_sva_2 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1548_nl) ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_8_sva_2 <= nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_8_sva_2[4:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_24U_11U_else_carry_8_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1549_nl) ) begin
      FpMantRNE_24U_11U_else_carry_8_sva_2 <= FpMantRNE_24U_11U_else_carry_8_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_9_sva_2 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1550_nl) ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_9_sva_2 <= nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_9_sva_2[4:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_24U_11U_else_carry_9_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1551_nl) ) begin
      FpMantRNE_24U_11U_else_carry_9_sva_2 <= FpMantRNE_24U_11U_else_carry_9_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_10_sva_2 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1552_nl) ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_10_sva_2 <= nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_10_sva_2[4:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_24U_11U_else_carry_10_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1553_nl) ) begin
      FpMantRNE_24U_11U_else_carry_10_sva_2 <= FpMantRNE_24U_11U_else_carry_10_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_11_sva_2 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1554_nl) ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_11_sva_2 <= nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_11_sva_2[4:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_24U_11U_else_carry_11_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1555_nl) ) begin
      FpMantRNE_24U_11U_else_carry_11_sva_2 <= FpMantRNE_24U_11U_else_carry_11_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_12_sva_2 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1556_nl) ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_12_sva_2 <= nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_12_sva_2[4:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_24U_11U_else_carry_12_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1557_nl) ) begin
      FpMantRNE_24U_11U_else_carry_12_sva_2 <= FpMantRNE_24U_11U_else_carry_12_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_13_sva_2 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1558_nl) ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_13_sva_2 <= nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_13_sva_2[4:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_24U_11U_else_carry_13_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1559_nl) ) begin
      FpMantRNE_24U_11U_else_carry_13_sva_2 <= FpMantRNE_24U_11U_else_carry_13_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_14_sva_2 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1560_nl) ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_14_sva_2 <= nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_14_sva_2[4:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_24U_11U_else_carry_14_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1561_nl) ) begin
      FpMantRNE_24U_11U_else_carry_14_sva_2 <= FpMantRNE_24U_11U_else_carry_14_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_15_sva_2 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1562_nl) ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_15_sva_2 <= nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_15_sva_2[4:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_24U_11U_else_carry_15_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1563_nl) ) begin
      FpMantRNE_24U_11U_else_carry_15_sva_2 <= FpMantRNE_24U_11U_else_carry_15_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva_2 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1564_nl) ) begin
      FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva_2 <= nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva_2[4:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_24U_11U_else_carry_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1565_nl) ) begin
      FpMantRNE_24U_11U_else_carry_sva_2 <= FpMantRNE_24U_11U_else_carry_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_sva_9 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_1569_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_sva_9 <= cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_4_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_16_FpMantRNE_24U_11U_else_and_4_svs_2 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_itm_8_1
        & (~ cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_itm_7_1) & cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_itm_8_1)
        | and_1321_rgt) & (~ mux_tmp_6) ) begin
      cvt_16_FpMantRNE_24U_11U_else_and_4_svs_2 <= MUX_s_1_2_2(cvt_16_FpMantRNE_24U_11U_else_and_4_tmp,
          cvt_16_FpMantRNE_24U_11U_else_and_4_svs, and_1321_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_sva_9 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_1573_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_sva_9 <= cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_15_FpMantRNE_24U_11U_else_and_3_svs_2 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1
        & (~ cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1) & cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1)
        | and_1325_rgt) & (~ mux_tmp_6) ) begin
      cvt_15_FpMantRNE_24U_11U_else_and_3_svs_2 <= MUX_s_1_2_2(cvt_15_FpMantRNE_24U_11U_else_and_3_tmp,
          cvt_15_FpMantRNE_24U_11U_else_and_3_svs, and_1325_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_sva_9 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_1577_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_sva_9 <= cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_14_FpMantRNE_24U_11U_else_and_3_svs_2 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1
        & (~ cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1) & cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1)
        | and_1329_rgt) & (~ mux_tmp_6) ) begin
      cvt_14_FpMantRNE_24U_11U_else_and_3_svs_2 <= MUX_s_1_2_2(cvt_14_FpMantRNE_24U_11U_else_and_3_tmp,
          cvt_14_FpMantRNE_24U_11U_else_and_3_svs, and_1329_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_sva_9 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_1581_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_sva_9 <= cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_13_FpMantRNE_24U_11U_else_and_2_svs_2 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1
        & (~ cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1) & cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1)
        | and_1333_rgt) & (~ mux_tmp_6) ) begin
      cvt_13_FpMantRNE_24U_11U_else_and_2_svs_2 <= MUX_s_1_2_2(cvt_13_FpMantRNE_24U_11U_else_and_2_tmp,
          cvt_13_FpMantRNE_24U_11U_else_and_2_svs, and_1333_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_sva_9 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_1585_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_sva_9 <= cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_12_FpMantRNE_24U_11U_else_and_3_svs_2 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1
        & (~ cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1) & cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1)
        | and_1337_rgt) & (~ mux_tmp_6) ) begin
      cvt_12_FpMantRNE_24U_11U_else_and_3_svs_2 <= MUX_s_1_2_2(cvt_12_FpMantRNE_24U_11U_else_and_3_tmp,
          cvt_12_FpMantRNE_24U_11U_else_and_3_svs, and_1337_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_sva_9 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_1589_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_sva_9 <= cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_11_FpMantRNE_24U_11U_else_and_2_svs_2 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1
        & (~ cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1) & cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1)
        | and_1341_rgt) & (~ mux_tmp_6) ) begin
      cvt_11_FpMantRNE_24U_11U_else_and_2_svs_2 <= MUX_s_1_2_2(cvt_11_FpMantRNE_24U_11U_else_and_2_tmp,
          cvt_11_FpMantRNE_24U_11U_else_and_2_svs, and_1341_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_sva_9 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1591_nl) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_sva_9 <= cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_10_FpMantRNE_24U_11U_else_and_2_svs_2 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1
        & (~ cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1) & cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1)
        | and_1345_rgt) & (~ mux_tmp_6) ) begin
      cvt_10_FpMantRNE_24U_11U_else_and_2_svs_2 <= MUX_s_1_2_2(cvt_10_FpMantRNE_24U_11U_else_and_2_tmp,
          cvt_10_FpMantRNE_24U_11U_else_and_2_svs, and_1345_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_sva_9 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_1595_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_sva_9 <= cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_9_FpMantRNE_24U_11U_else_and_1_svs_2 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1
        & (~ cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1) & cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1)
        | and_1349_rgt) & (~ mux_tmp_6) ) begin
      cvt_9_FpMantRNE_24U_11U_else_and_1_svs_2 <= MUX_s_1_2_2(cvt_9_FpMantRNE_24U_11U_else_and_1_tmp,
          cvt_9_FpMantRNE_24U_11U_else_and_1_svs, and_1349_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_sva_9 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_1599_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_sva_9 <= cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_8_FpMantRNE_24U_11U_else_and_3_svs_2 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1
        & (~ cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1) & cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1)
        | and_1353_rgt) & (~ mux_tmp_6) ) begin
      cvt_8_FpMantRNE_24U_11U_else_and_3_svs_2 <= MUX_s_1_2_2(cvt_8_FpMantRNE_24U_11U_else_and_3_tmp,
          cvt_8_FpMantRNE_24U_11U_else_and_3_svs, and_1353_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_sva_9 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_1603_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_sva_9 <= cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_7_FpMantRNE_24U_11U_else_and_2_svs_2 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1
        & (~ cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1) & cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1)
        | and_1357_rgt) & (~ mux_tmp_6) ) begin
      cvt_7_FpMantRNE_24U_11U_else_and_2_svs_2 <= MUX_s_1_2_2(cvt_7_FpMantRNE_24U_11U_else_and_2_tmp,
          cvt_7_FpMantRNE_24U_11U_else_and_2_svs, and_1357_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_sva_9 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1605_nl) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_sva_9 <= cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_6_FpMantRNE_24U_11U_else_and_2_svs_2 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1
        & (~ cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1) & cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1)
        | and_1361_rgt) & (~ mux_tmp_6) ) begin
      cvt_6_FpMantRNE_24U_11U_else_and_2_svs_2 <= MUX_s_1_2_2(cvt_6_FpMantRNE_24U_11U_else_and_2_tmp,
          cvt_6_FpMantRNE_24U_11U_else_and_2_svs, and_1361_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_sva_9 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_1609_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_sva_9 <= cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_5_FpMantRNE_24U_11U_else_and_1_svs_2 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1
        & (~ cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1) & cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1)
        | and_1365_rgt) & (~ mux_tmp_6) ) begin
      cvt_5_FpMantRNE_24U_11U_else_and_1_svs_2 <= MUX_s_1_2_2(cvt_5_FpMantRNE_24U_11U_else_and_1_tmp,
          cvt_5_FpMantRNE_24U_11U_else_and_1_svs, and_1365_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_sva_9 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_1613_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_sva_9 <= cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_4_FpMantRNE_24U_11U_else_and_2_svs_2 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1
        & (~ cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1) & cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1)
        | and_1369_rgt) & (~ mux_tmp_6) ) begin
      cvt_4_FpMantRNE_24U_11U_else_and_2_svs_2 <= MUX_s_1_2_2(cvt_4_FpMantRNE_24U_11U_else_and_2_tmp,
          cvt_4_FpMantRNE_24U_11U_else_and_2_svs, and_1369_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_sva_9 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_1617_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_sva_9 <= cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_3_FpMantRNE_24U_11U_else_and_1_svs_2 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1
        & (~ cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1) & cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1)
        | and_1373_rgt) & (~ mux_tmp_6) ) begin
      cvt_3_FpMantRNE_24U_11U_else_and_1_svs_2 <= MUX_s_1_2_2(cvt_3_FpMantRNE_24U_11U_else_and_1_tmp,
          cvt_3_FpMantRNE_24U_11U_else_and_1_svs, and_1373_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_sva_9 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_1621_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_sva_9 <= cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_2_FpMantRNE_24U_11U_else_and_1_svs_2 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1
        & (~ cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1) & cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1)
        | and_1377_rgt) & (~ mux_tmp_6) ) begin
      cvt_2_FpMantRNE_24U_11U_else_and_1_svs_2 <= MUX_s_1_2_2(cvt_2_FpMantRNE_24U_11U_else_and_1_tmp,
          cvt_2_FpMantRNE_24U_11U_else_and_1_svs, and_1377_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_sva_9 <= 5'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (~ (mux_1625_nl)) ) begin
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_sva_9 <= cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_1_FpMantRNE_24U_11U_else_and_svs_2 <= 1'b0;
    end
    else if ( core_wen & ((or_5189_cse & cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_itm_8_1
        & (~ cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1) & cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_itm_8_1)
        | and_1381_rgt) & (~ mux_tmp_6) ) begin
      cvt_1_FpMantRNE_24U_11U_else_and_svs_2 <= MUX_s_1_2_2(cvt_1_FpMantRNE_24U_11U_else_and_tmp,
          cvt_1_FpMantRNE_24U_11U_else_and_svs, and_1381_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_17U_16U_o_15_1_lpi_1_dfm_9 <= 15'b0;
    end
    else if ( core_wen & (IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_rgt
        | IntSaturation_17U_16U_and_31_rgt | IntSaturation_17U_16U_o_and_31_rgt)
        & mux_tmp_161 ) begin
      IntSaturation_17U_16U_o_15_1_lpi_1_dfm_9 <= MUX1HOT_v_15_3_2(IntShiftRightSat_49U_6U_17U_o_15_1_sva_mx0w0,
          15'b100000000000000, 15'b11111111111111, {IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_rgt
          , IntSaturation_17U_16U_and_31_rgt , IntSaturation_17U_16U_o_and_31_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_17U_16U_o_15_1_15_lpi_1_dfm_8 <= 15'b0;
    end
    else if ( core_wen & (IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_1_rgt
        | IntSaturation_17U_16U_and_29_rgt | IntSaturation_17U_16U_o_and_29_rgt)
        & mux_tmp_161 ) begin
      IntSaturation_17U_16U_o_15_1_15_lpi_1_dfm_8 <= MUX1HOT_v_15_3_2(IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_mx0w0,
          15'b100000000000000, 15'b11111111111111, {IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_1_rgt
          , IntSaturation_17U_16U_and_29_rgt , IntSaturation_17U_16U_o_and_29_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_17U_16U_o_15_1_14_lpi_1_dfm_8 <= 15'b0;
    end
    else if ( core_wen & (IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_2_rgt
        | IntSaturation_17U_16U_and_27_rgt | IntSaturation_17U_16U_o_and_27_rgt)
        & mux_tmp_161 ) begin
      IntSaturation_17U_16U_o_15_1_14_lpi_1_dfm_8 <= MUX1HOT_v_15_3_2(IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_mx0w0,
          15'b100000000000000, 15'b11111111111111, {IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_2_rgt
          , IntSaturation_17U_16U_and_27_rgt , IntSaturation_17U_16U_o_and_27_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_17U_16U_o_15_1_13_lpi_1_dfm_7 <= 15'b0;
    end
    else if ( core_wen & (IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_3_rgt
        | IntSaturation_17U_16U_and_25_rgt | IntSaturation_17U_16U_o_and_25_rgt)
        & mux_tmp_161 ) begin
      IntSaturation_17U_16U_o_15_1_13_lpi_1_dfm_7 <= MUX1HOT_v_15_3_2(IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_mx0w0,
          15'b100000000000000, 15'b11111111111111, {IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_3_rgt
          , IntSaturation_17U_16U_and_25_rgt , IntSaturation_17U_16U_o_and_25_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_17U_16U_o_15_1_12_lpi_1_dfm_8 <= 15'b0;
    end
    else if ( core_wen & (IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_4_rgt
        | IntSaturation_17U_16U_and_23_rgt | IntSaturation_17U_16U_o_and_23_rgt)
        & mux_tmp_161 ) begin
      IntSaturation_17U_16U_o_15_1_12_lpi_1_dfm_8 <= MUX1HOT_v_15_3_2(IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_mx0w0,
          15'b100000000000000, 15'b11111111111111, {IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_4_rgt
          , IntSaturation_17U_16U_and_23_rgt , IntSaturation_17U_16U_o_and_23_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_17U_16U_o_15_1_11_lpi_1_dfm_7 <= 15'b0;
    end
    else if ( core_wen & (IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_5_rgt
        | IntSaturation_17U_16U_and_21_rgt | IntSaturation_17U_16U_o_and_21_rgt)
        & mux_tmp_161 ) begin
      IntSaturation_17U_16U_o_15_1_11_lpi_1_dfm_7 <= MUX1HOT_v_15_3_2(IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_mx0w0,
          15'b100000000000000, 15'b11111111111111, {IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_5_rgt
          , IntSaturation_17U_16U_and_21_rgt , IntSaturation_17U_16U_o_and_21_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_17U_16U_o_15_1_10_lpi_1_dfm_7 <= 15'b0;
    end
    else if ( core_wen & (IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_6_rgt
        | IntSaturation_17U_16U_and_19_rgt | IntSaturation_17U_16U_o_and_19_rgt)
        & mux_tmp_161 ) begin
      IntSaturation_17U_16U_o_15_1_10_lpi_1_dfm_7 <= MUX1HOT_v_15_3_2(IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_mx0w0,
          15'b100000000000000, 15'b11111111111111, {IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_6_rgt
          , IntSaturation_17U_16U_and_19_rgt , IntSaturation_17U_16U_o_and_19_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_17U_16U_o_15_1_9_lpi_1_dfm_6 <= 15'b0;
    end
    else if ( core_wen & (IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_7_rgt
        | IntSaturation_17U_16U_and_17_rgt | IntSaturation_17U_16U_o_and_17_rgt)
        & mux_tmp_161 ) begin
      IntSaturation_17U_16U_o_15_1_9_lpi_1_dfm_6 <= MUX1HOT_v_15_3_2(IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_mx0w0,
          15'b100000000000000, 15'b11111111111111, {IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_7_rgt
          , IntSaturation_17U_16U_and_17_rgt , IntSaturation_17U_16U_o_and_17_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_17U_16U_o_15_1_8_lpi_1_dfm_8 <= 15'b0;
    end
    else if ( core_wen & (IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_8_rgt
        | IntSaturation_17U_16U_and_15_rgt | IntSaturation_17U_16U_o_and_15_rgt)
        & mux_tmp_161 ) begin
      IntSaturation_17U_16U_o_15_1_8_lpi_1_dfm_8 <= MUX1HOT_v_15_3_2(IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_mx0w0,
          15'b100000000000000, 15'b11111111111111, {IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_8_rgt
          , IntSaturation_17U_16U_and_15_rgt , IntSaturation_17U_16U_o_and_15_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_17U_16U_o_15_1_7_lpi_1_dfm_7 <= 15'b0;
    end
    else if ( core_wen & (IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_9_rgt
        | IntSaturation_17U_16U_and_13_rgt | IntSaturation_17U_16U_o_and_13_rgt)
        & mux_tmp_161 ) begin
      IntSaturation_17U_16U_o_15_1_7_lpi_1_dfm_7 <= MUX1HOT_v_15_3_2(IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_mx0w0,
          15'b100000000000000, 15'b11111111111111, {IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_9_rgt
          , IntSaturation_17U_16U_and_13_rgt , IntSaturation_17U_16U_o_and_13_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_17U_16U_o_15_1_6_lpi_1_dfm_7 <= 15'b0;
    end
    else if ( core_wen & (IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_10_rgt
        | IntSaturation_17U_16U_and_11_rgt | IntSaturation_17U_16U_o_and_11_rgt)
        & mux_tmp_161 ) begin
      IntSaturation_17U_16U_o_15_1_6_lpi_1_dfm_7 <= MUX1HOT_v_15_3_2(IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_mx0w0,
          15'b100000000000000, 15'b11111111111111, {IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_10_rgt
          , IntSaturation_17U_16U_and_11_rgt , IntSaturation_17U_16U_o_and_11_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_17U_16U_o_15_1_5_lpi_1_dfm_6 <= 15'b0;
    end
    else if ( core_wen & (IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_11_rgt
        | IntSaturation_17U_16U_and_9_rgt | IntSaturation_17U_16U_o_and_9_rgt) &
        mux_tmp_161 ) begin
      IntSaturation_17U_16U_o_15_1_5_lpi_1_dfm_6 <= MUX1HOT_v_15_3_2(IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_mx0w0,
          15'b100000000000000, 15'b11111111111111, {IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_11_rgt
          , IntSaturation_17U_16U_and_9_rgt , IntSaturation_17U_16U_o_and_9_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_17U_16U_o_15_1_4_lpi_1_dfm_7 <= 15'b0;
    end
    else if ( core_wen & (IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_12_rgt
        | IntSaturation_17U_16U_and_7_rgt | IntSaturation_17U_16U_o_and_7_rgt) &
        mux_tmp_161 ) begin
      IntSaturation_17U_16U_o_15_1_4_lpi_1_dfm_7 <= MUX1HOT_v_15_3_2(IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_mx0w0,
          15'b100000000000000, 15'b11111111111111, {IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_12_rgt
          , IntSaturation_17U_16U_and_7_rgt , IntSaturation_17U_16U_o_and_7_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_17U_16U_o_15_1_3_lpi_1_dfm_6 <= 15'b0;
    end
    else if ( core_wen & (IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_13_rgt
        | IntSaturation_17U_16U_and_5_rgt | IntSaturation_17U_16U_o_and_5_rgt) &
        mux_tmp_161 ) begin
      IntSaturation_17U_16U_o_15_1_3_lpi_1_dfm_6 <= MUX1HOT_v_15_3_2(IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_mx0w0,
          15'b100000000000000, 15'b11111111111111, {IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_13_rgt
          , IntSaturation_17U_16U_and_5_rgt , IntSaturation_17U_16U_o_and_5_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_17U_16U_o_15_1_2_lpi_1_dfm_6 <= 15'b0;
    end
    else if ( core_wen & (IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_14_rgt
        | IntSaturation_17U_16U_and_3_rgt | IntSaturation_17U_16U_o_and_3_rgt) &
        mux_tmp_161 ) begin
      IntSaturation_17U_16U_o_15_1_2_lpi_1_dfm_6 <= MUX1HOT_v_15_3_2(IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_mx0w0,
          15'b100000000000000, 15'b11111111111111, {IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_14_rgt
          , IntSaturation_17U_16U_and_3_rgt , IntSaturation_17U_16U_o_and_3_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_17U_16U_o_15_1_1_lpi_1_dfm_5 <= 15'b0;
    end
    else if ( core_wen & (IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_15_rgt
        | IntSaturation_17U_16U_and_1_rgt | IntSaturation_17U_16U_o_and_1_rgt) &
        mux_tmp_161 ) begin
      IntSaturation_17U_16U_o_15_1_1_lpi_1_dfm_5 <= MUX1HOT_v_15_3_2(IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_mx0w0,
          15'b100000000000000, 15'b11111111111111, {IntSaturation_17U_16U_o_IntSaturation_17U_16U_o_nor_15_rgt
          , IntSaturation_17U_16U_and_1_rgt , IntSaturation_17U_16U_o_and_1_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_8_itm_2 <= 1'b0;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_4_itm_2 <= 1'b0;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_2_itm_2 <= 1'b0;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_itm_2 <= 1'b0;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_15_itm_2 <= 1'b0;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_14_itm_2 <= 1'b0;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_12_itm_2 <= 1'b0;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_11_itm_2 <= 1'b0;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_10_itm_2 <= 1'b0;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_9_itm_2 <= 1'b0;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_7_itm_2 <= 1'b0;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_6_itm_2 <= 1'b0;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_5_itm_2 <= 1'b0;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_3_itm_2 <= 1'b0;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_1_itm_2 <= 1'b0;
    end
    else if ( IntSaturation_17U_16U_and_33_cse ) begin
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_8_itm_2 <= (IntShiftRightSat_49U_6U_17U_o_0_9_sva_mx0w0
          & (~ cvt_9_IntSaturation_17U_16U_else_if_acc_1_itm_2_1)) | cvt_9_IntSaturation_17U_16U_if_acc_1_itm_2_1;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_4_itm_2 <= (IntShiftRightSat_49U_6U_17U_o_0_5_sva_mx0w0
          & (~ cvt_5_IntSaturation_17U_16U_else_if_acc_1_itm_2_1)) | cvt_5_IntSaturation_17U_16U_if_acc_1_itm_2_1;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_2_itm_2 <= (IntShiftRightSat_49U_6U_17U_o_0_3_sva_mx0w0
          & (~ cvt_3_IntSaturation_17U_16U_else_if_acc_1_itm_2_1)) | cvt_3_IntSaturation_17U_16U_if_acc_1_itm_2_1;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_itm_2 <= (IntShiftRightSat_49U_6U_17U_o_0_1_sva_mx0w0
          & (~ cvt_1_IntSaturation_17U_16U_else_if_acc_itm_2_1)) | cvt_1_IntSaturation_17U_16U_if_acc_itm_2_1;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_15_itm_2 <= (IntShiftRightSat_49U_6U_17U_o_0_sva_mx0w0
          & (~ cvt_16_IntSaturation_17U_16U_else_if_acc_4_itm_2_1)) | cvt_16_IntSaturation_17U_16U_if_acc_4_itm_2_1;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_14_itm_2 <= (IntShiftRightSat_49U_6U_17U_o_0_15_sva_mx0w0
          & (~ cvt_15_IntSaturation_17U_16U_else_if_acc_3_itm_2_1)) | cvt_15_IntSaturation_17U_16U_if_acc_3_itm_2_1;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_12_itm_2 <= (IntShiftRightSat_49U_6U_17U_o_0_13_sva_mx0w0
          & (~ cvt_13_IntSaturation_17U_16U_else_if_acc_2_itm_2_1)) | cvt_13_IntSaturation_17U_16U_if_acc_2_itm_2_1;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_11_itm_2 <= (IntShiftRightSat_49U_6U_17U_o_0_12_sva_mx0w0
          & (~ cvt_12_IntSaturation_17U_16U_else_if_acc_3_itm_2_1)) | cvt_12_IntSaturation_17U_16U_if_acc_3_itm_2_1;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_10_itm_2 <= (IntShiftRightSat_49U_6U_17U_o_0_11_sva_mx0w0
          & (~ cvt_11_IntSaturation_17U_16U_else_if_acc_2_itm_2_1)) | cvt_11_IntSaturation_17U_16U_if_acc_2_itm_2_1;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_9_itm_2 <= (IntShiftRightSat_49U_6U_17U_o_0_10_sva_mx0w0
          & (~ cvt_10_IntSaturation_17U_16U_else_if_acc_2_itm_2_1)) | cvt_10_IntSaturation_17U_16U_if_acc_2_itm_2_1;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_7_itm_2 <= (IntShiftRightSat_49U_6U_17U_o_0_8_sva_mx0w0
          & (~ cvt_8_IntSaturation_17U_16U_else_if_acc_3_itm_2_1)) | cvt_8_IntSaturation_17U_16U_if_acc_3_itm_2_1;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_6_itm_2 <= (IntShiftRightSat_49U_6U_17U_o_0_7_sva_mx0w0
          & (~ cvt_7_IntSaturation_17U_16U_else_if_acc_2_itm_2_1)) | cvt_7_IntSaturation_17U_16U_if_acc_2_itm_2_1;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_5_itm_2 <= (IntShiftRightSat_49U_6U_17U_o_0_6_sva_mx0w0
          & (~ cvt_6_IntSaturation_17U_16U_else_if_acc_2_itm_2_1)) | cvt_6_IntSaturation_17U_16U_if_acc_2_itm_2_1;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_3_itm_2 <= (IntShiftRightSat_49U_6U_17U_o_0_4_sva_mx0w0
          & (~ cvt_4_IntSaturation_17U_16U_else_if_acc_2_itm_2_1)) | cvt_4_IntSaturation_17U_16U_if_acc_2_itm_2_1;
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_1_itm_2 <= (IntShiftRightSat_49U_6U_17U_o_0_2_sva_mx0w0
          & (~ cvt_2_IntSaturation_17U_16U_else_if_acc_1_itm_2_1)) | cvt_2_IntSaturation_17U_16U_if_acc_1_itm_2_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_idata_data_sva_2_15_0_1 <= 16'b0;
    end
    else if ( core_wen & (~ and_dcpl_93) & (mux_1627_nl) ) begin
      chn_idata_data_sva_2_15_0_1 <= chn_idata_data_sva_1_27_0_1[15:0];
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_5U_10U_nor_itm_2 <= 1'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_27_cse
        & (mux_1640_nl) ) begin
      IsNaN_5U_10U_nor_itm_2 <= MUX_s_1_2_2((IsNaN_5U_10U_nor_nl), cvt_16_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_4_tmp,
          and_dcpl_204);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_5U_10U_IsNaN_5U_10U_nand_itm_2 <= 1'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_27_cse
        & (mux_1649_nl) ) begin
      IsNaN_5U_10U_IsNaN_5U_10U_nand_itm_2 <= MUX_s_1_2_2((IsNaN_5U_10U_IsNaN_5U_10U_nand_nl),
          cvt_13_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp,
          and_dcpl_204);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_5U_10U_nor_1_itm_2 <= 1'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_27_cse
        & (mux_1660_nl) ) begin
      IsNaN_5U_10U_nor_1_itm_2 <= MUX_s_1_2_2((IsNaN_5U_10U_nor_1_nl), cvt_14_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp,
          and_dcpl_204);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_5U_10U_IsNaN_5U_10U_nand_1_itm_2 <= 1'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_27_cse
        & (mux_1663_nl) ) begin
      IsNaN_5U_10U_IsNaN_5U_10U_nand_1_itm_2 <= MUX_s_1_2_2((IsNaN_5U_10U_IsNaN_5U_10U_nand_1_nl),
          cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_tmp, and_dcpl_204);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_5U_10U_nor_14_itm_2 <= 1'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_27_cse
        & (mux_1674_nl) ) begin
      IsNaN_5U_10U_nor_14_itm_2 <= MUX_s_1_2_2((IsNaN_5U_10U_nor_14_nl), cvt_15_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp,
          and_dcpl_204);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_5U_10U_IsNaN_5U_10U_nand_14_itm_2 <= 1'b0;
    end
    else if ( core_wen & IntShiftRightSat_49U_6U_17U_o_IntShiftRightSat_49U_6U_17U_o_or_27_cse
        & (mux_1685_nl) ) begin
      IsNaN_5U_10U_IsNaN_5U_10U_nand_14_itm_2 <= MUX_s_1_2_2((IsNaN_5U_10U_IsNaN_5U_10U_nand_14_nl),
          cvt_12_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp,
          and_dcpl_204);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_lor_3_lpi_1_dfm <= 1'b0;
      IntShiftRightSat_49U_6U_17U_lor_4_lpi_1_dfm <= 1'b0;
    end
    else if ( IntShiftRightSat_49U_6U_17U_oelse_and_cse ) begin
      IntShiftRightSat_49U_6U_17U_lor_3_lpi_1_dfm <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_3_lpi_1_dfm_mx1w0,
          cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp,
          and_1385_rgt);
      IntShiftRightSat_49U_6U_17U_lor_4_lpi_1_dfm <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_4_lpi_1_dfm_mx1w0,
          cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp,
          and_1385_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_lor_5_lpi_1_dfm <= 1'b0;
    end
    else if ( cvt_else_and_cse & IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_18_cse
        & mux_320_cse ) begin
      IntShiftRightSat_49U_6U_17U_lor_5_lpi_1_dfm <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_5_lpi_1_dfm_mx1w0,
          cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp,
          and_1385_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_lor_7_lpi_1_dfm <= 1'b0;
      IntShiftRightSat_49U_6U_17U_lor_8_lpi_1_dfm <= 1'b0;
    end
    else if ( IntShiftRightSat_49U_6U_17U_oelse_and_18_cse ) begin
      IntShiftRightSat_49U_6U_17U_lor_7_lpi_1_dfm <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_7_lpi_1_dfm_mx1w0,
          cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp,
          and_1385_rgt);
      IntShiftRightSat_49U_6U_17U_lor_8_lpi_1_dfm <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_8_lpi_1_dfm_mx1w0,
          cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp,
          and_1385_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_lor_9_lpi_1_dfm <= 1'b0;
    end
    else if ( cvt_else_and_cse & IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_15_cse
        & (mux_449_nl) ) begin
      IntShiftRightSat_49U_6U_17U_lor_9_lpi_1_dfm <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_9_lpi_1_dfm_mx1w0,
          cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp,
          and_1385_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_lor_6_lpi_1_dfm <= 1'b0;
    end
    else if ( cvt_else_and_cse & IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_19_cse
        & (mux_454_nl) ) begin
      IntShiftRightSat_49U_6U_17U_lor_6_lpi_1_dfm <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_6_lpi_1_dfm_mx1w0,
          cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp,
          and_1385_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_lor_11_lpi_1_dfm <= 1'b0;
      IntShiftRightSat_49U_6U_17U_lor_12_lpi_1_dfm <= 1'b0;
    end
    else if ( IntShiftRightSat_49U_6U_17U_oelse_and_22_cse ) begin
      IntShiftRightSat_49U_6U_17U_lor_11_lpi_1_dfm <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_11_lpi_1_dfm_mx1w0,
          cvt_10_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp,
          and_1385_rgt);
      IntShiftRightSat_49U_6U_17U_lor_12_lpi_1_dfm <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_12_lpi_1_dfm_mx1w0,
          cvt_11_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp,
          and_1385_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_lor_13_lpi_1_dfm <= 1'b0;
    end
    else if ( cvt_else_and_cse & IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_15_cse
        & mux_272_cse ) begin
      IntShiftRightSat_49U_6U_17U_lor_13_lpi_1_dfm <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_13_lpi_1_dfm_mx1w0,
          cvt_12_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp,
          and_1385_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_lor_15_lpi_1_dfm <= 1'b0;
      IntShiftRightSat_49U_6U_17U_lor_14_lpi_1_dfm <= 1'b0;
    end
    else if ( IntShiftRightSat_49U_6U_17U_oelse_and_25_cse ) begin
      IntShiftRightSat_49U_6U_17U_lor_15_lpi_1_dfm <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_15_lpi_1_dfm_mx1w0,
          cvt_14_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp,
          and_1385_rgt);
      IntShiftRightSat_49U_6U_17U_lor_14_lpi_1_dfm <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_14_lpi_1_dfm_mx1w0,
          cvt_13_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp,
          and_1385_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_lor_lpi_1_dfm <= 1'b0;
    end
    else if ( cvt_else_and_cse & IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_8_cse
        & (mux_770_nl) ) begin
      IntShiftRightSat_49U_6U_17U_lor_lpi_1_dfm <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_lpi_1_dfm_mx1w0,
          cvt_16_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_4_tmp,
          and_1385_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_lor_16_lpi_1_dfm <= 1'b0;
    end
    else if ( cvt_else_and_cse & IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_8_cse
        & (mux_789_nl) ) begin
      IntShiftRightSat_49U_6U_17U_lor_16_lpi_1_dfm <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_16_lpi_1_dfm_mx1w0,
          cvt_15_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp,
          and_1385_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_lor_10_lpi_1_dfm <= 1'b0;
    end
    else if ( cvt_else_and_cse & IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_oelse_or_19_cse
        & (mux_799_nl) ) begin
      IntShiftRightSat_49U_6U_17U_lor_10_lpi_1_dfm <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_10_lpi_1_dfm_mx1w0,
          cvt_10_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp,
          and_1385_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_lor_2_lpi_1_dfm <= 1'b0;
    end
    else if ( cvt_else_and_cse & ((or_dcpl_386 & or_4862_cse & and_dcpl_401) | and_1467_rgt)
        & (mux_803_nl) ) begin
      IntShiftRightSat_49U_6U_17U_lor_2_lpi_1_dfm <= MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_2_lpi_1_dfm_mx1w0,
          cvt_11_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp,
          and_1467_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_1_FpMantRNE_17U_11U_else_and_svs <= 1'b0;
    end
    else if ( core_wen & (~(and_dcpl_942 | (~ or_4862_cse) | and_dcpl_93 | cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_svs_st_2
        | or_dcpl_389)) ) begin
      cvt_1_FpMantRNE_17U_11U_else_and_svs <= cvt_1_FpMantRNE_17U_11U_else_and_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp <= 1'b0;
    end
    else if ( cvt_else_and_cse & (~((~ or_4862_cse) | cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_svs_st_2
        | or_dcpl_389)) & mux_tmp_245 ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp <= or_1202_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_2_FpMantRNE_17U_11U_else_and_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(and_dcpl_946 | or_dcpl_151 | or_dcpl_399 | cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2
        | (cfg_out_precision_1_sva_st_149!=2'b10))) ) begin
      cvt_2_FpMantRNE_17U_11U_else_and_1_svs <= cvt_2_FpMantRNE_17U_11U_else_and_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_1 <= 1'b0;
    end
    else if ( cvt_else_and_cse & (~(or_dcpl_151 | (~ main_stage_v_2) | cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2
        | (cfg_out_precision_1_sva_st_149!=2'b10))) & (mux_1687_nl) ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_1 <= or_1596_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_3_FpMantRNE_17U_11U_else_and_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(and_dcpl_950 | (~ and_tmp_50) | or_dcpl_399 | cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2
        | (cfg_out_precision_1_sva_st_149!=2'b10))) ) begin
      cvt_3_FpMantRNE_17U_11U_else_and_1_svs <= cvt_3_FpMantRNE_17U_11U_else_and_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_2 <= 1'b0;
    end
    else if ( cvt_else_and_cse & (~((~ and_tmp_50) | (~ main_stage_v_2) | cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2
        | (cfg_out_precision_1_sva_st_149!=2'b10))) & (mux_1689_nl) ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_2 <= or_1625_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_4_FpMantRNE_17U_11U_else_and_2_svs <= 1'b0;
    end
    else if ( core_wen & (~(and_dcpl_954 | (~ and_tmp_50) | and_1021_cse | and_dcpl_93
        | or_dcpl_420)) ) begin
      cvt_4_FpMantRNE_17U_11U_else_and_2_svs <= cvt_4_FpMantRNE_17U_11U_else_and_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_3 <= 1'b0;
    end
    else if ( cvt_else_and_cse & (~(or_dcpl_353 | or_dcpl_420)) & (mux_1692_nl) )
        begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_3 <= or_1659_cse_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_5_FpMantRNE_17U_11U_else_and_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(and_dcpl_958 | or_dcpl_163 | or_dcpl_399 | (cfg_out_precision_1_sva_st_149!=2'b10)
        | cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2))
        ) begin
      cvt_5_FpMantRNE_17U_11U_else_and_1_svs <= cvt_5_FpMantRNE_17U_11U_else_and_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_4 <= 1'b0;
    end
    else if ( cvt_else_and_cse & (~(or_dcpl_163 | (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
        | cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2))
        & (mux_1694_nl) ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_4 <= or_1693_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_6_FpMantRNE_17U_11U_else_and_2_svs <= 1'b0;
    end
    else if ( core_wen & (~(and_dcpl_962 | or_dcpl_163 | and_1021_cse | and_dcpl_93
        | or_dcpl_439)) ) begin
      cvt_6_FpMantRNE_17U_11U_else_and_2_svs <= cvt_6_FpMantRNE_17U_11U_else_and_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_5 <= 1'b0;
    end
    else if ( cvt_else_and_cse & (~(or_3774_cse | or_dcpl_439)) & (mux_1697_nl) )
        begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_5 <= or_1720_cse_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_7_FpMantRNE_17U_11U_else_and_2_svs <= 1'b0;
    end
    else if ( core_wen & (~(and_dcpl_966 | or_dcpl_163 | and_1021_cse | and_dcpl_93
        | or_dcpl_448)) ) begin
      cvt_7_FpMantRNE_17U_11U_else_and_2_svs <= cvt_7_FpMantRNE_17U_11U_else_and_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_6 <= 1'b0;
    end
    else if ( cvt_else_and_cse & (~(or_3774_cse | or_dcpl_448)) & (mux_1700_nl) )
        begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_6 <= or_1752_cse_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_8_FpMantRNE_17U_11U_else_and_3_svs <= 1'b0;
    end
    else if ( core_wen & (~(and_dcpl_970 | (~ or_4862_cse) | and_dcpl_479 | and_1021_cse
        | and_dcpl_93 | (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
        | FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_3)) ) begin
      cvt_8_FpMantRNE_17U_11U_else_and_3_svs <= cvt_8_FpMantRNE_17U_11U_else_and_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_7 <= 1'b0;
    end
    else if ( cvt_else_and_cse & (~(or_3774_cse | (~ main_stage_v_2) | or_578_cse
        | FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_3)) & (mux_1704_nl) ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_7 <= or_1789_cse_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_9_FpMantRNE_17U_11U_else_and_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(and_dcpl_974 | (~ mux_tmp_455) | or_dcpl_399 | (cfg_out_precision_1_sva_st_149!=2'b10)
        | cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2))
        ) begin
      cvt_9_FpMantRNE_17U_11U_else_and_1_svs <= cvt_9_FpMantRNE_17U_11U_else_and_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_8 <= 1'b0;
    end
    else if ( cvt_else_and_cse & (~((~ mux_tmp_455) | (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
        | cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2))
        & (mux_1707_nl) ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_8 <= or_1829_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_10_FpMantRNE_17U_11U_else_and_2_svs <= 1'b0;
    end
    else if ( core_wen & (~(and_dcpl_978 | (~ mux_tmp_455) | and_1021_cse | or_dcpl_480
        | and_dcpl_93 | or_578_cse)) ) begin
      cvt_10_FpMantRNE_17U_11U_else_and_2_svs <= cvt_10_FpMantRNE_17U_11U_else_and_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_9 <= 1'b0;
    end
    else if ( cvt_else_and_cse & (~(or_3817_cse | or_dcpl_480 | or_578_cse)) & (mux_1711_nl)
        ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_9 <= or_1851_cse_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_11_FpMantRNE_17U_11U_else_and_2_svs <= 1'b0;
    end
    else if ( core_wen & (~(and_dcpl_982 | (~ mux_tmp_455) | and_1021_cse | and_dcpl_93
        | or_dcpl_490)) ) begin
      cvt_11_FpMantRNE_17U_11U_else_and_2_svs <= cvt_11_FpMantRNE_17U_11U_else_and_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_10 <= 1'b0;
    end
    else if ( cvt_else_and_cse & (~(or_3817_cse | or_dcpl_490)) & (mux_1715_nl) )
        begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_10 <= or_1892_cse_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_12_FpMantRNE_17U_11U_else_and_3_svs <= 1'b0;
    end
    else if ( core_wen & (~(and_dcpl_987 | (~ or_4862_cse) | and_dcpl_479 | and_1021_cse
        | (cfg_out_precision_1_sva_st_149!=2'b10) | FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_3
        | (~ main_stage_v_2) | and_dcpl_93)) ) begin
      cvt_12_FpMantRNE_17U_11U_else_and_3_svs <= cvt_12_FpMantRNE_17U_11U_else_and_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_11 <= 1'b0;
    end
    else if ( cvt_else_and_cse & (~(or_3817_cse | (cfg_out_precision_1_sva_st_149!=2'b10)
        | FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_3 | (~ main_stage_v_2))) &
        mux_tmp_585 ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_11 <= or_1925_cse_1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_13_FpMantRNE_17U_11U_else_and_2_svs <= 1'b0;
    end
    else if ( core_wen & (~(and_dcpl_991 | (~ mux_tmp_455) | (cfg_out_precision_1_sva_st_149!=2'b10)
        | FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_3 | (~ main_stage_v_2) | or_dcpl_511))
        ) begin
      cvt_13_FpMantRNE_17U_11U_else_and_2_svs <= cvt_13_FpMantRNE_17U_11U_else_and_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_12 <= 1'b0;
    end
    else if ( cvt_else_and_cse & (~(or_tmp_3025 | (~ (cfg_out_precision_1_sva_st_149[1]))
        | FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_3 | (~ main_stage_v_2) | and_1021_cse))
        & (mux_1720_nl) ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_12 <= or_5038_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_14_FpMantRNE_17U_11U_else_and_3_svs <= 1'b0;
    end
    else if ( core_wen & (~(and_dcpl_995 | (~ or_4862_cse) | and_dcpl_479 | or_578_cse
        | (~ main_stage_v_2) | FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2 | or_dcpl_511))
        ) begin
      cvt_14_FpMantRNE_17U_11U_else_and_3_svs <= cvt_14_FpMantRNE_17U_11U_else_and_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_13 <= 1'b0;
    end
    else if ( cvt_else_and_cse & (~((~ mux_1142_cse) | or_578_cse | (~ main_stage_v_2)
        | FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2)) & (mux_1727_nl) ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_13 <= or_5053_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_15_FpMantRNE_17U_11U_else_and_3_svs <= 1'b0;
    end
    else if ( core_wen & (~(and_dcpl_999 | (~ or_4862_cse) | and_dcpl_479 | or_578_cse
        | and_dcpl_93 | and_1021_cse | (~ main_stage_v_2) | FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_3))
        ) begin
      cvt_15_FpMantRNE_17U_11U_else_and_3_svs <= cvt_15_FpMantRNE_17U_11U_else_and_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_14 <= 1'b0;
    end
    else if ( cvt_else_and_cse & (~((~ and_tmp_225) | or_578_cse | (~ main_stage_v_2)
        | FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_3)) & (mux_1734_nl) ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_14 <= or_5069_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_16_FpMantRNE_17U_11U_else_and_4_svs <= 1'b0;
    end
    else if ( core_wen & (~(and_dcpl_1003 | (~ mux_tmp_455) | or_dcpl_277 | (~ (cfg_out_precision_1_sva_st_149[1]))
        | FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_3 | or_dcpl_511)) ) begin
      cvt_16_FpMantRNE_17U_11U_else_and_4_svs <= cvt_16_FpMantRNE_17U_11U_else_and_4_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_15 <= 1'b0;
    end
    else if ( cvt_else_and_cse & (~((~ mux_tmp_455) | or_dcpl_277 | (~ (cfg_out_precision_1_sva_st_149[1]))
        | and_1021_cse | FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_3)) & (mux_1743_nl)
        ) begin
      FpIntToFloat_17U_5U_10U_else_unequal_tmp_15 <= or_5086_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_3 <= 1'b0;
      FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_3 <= 1'b0;
      FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_3 <= 1'b0;
      FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_3 <= 1'b0;
      FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( FpIntToFloat_17U_5U_10U_is_inf_and_28_cse ) begin
      FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_3 <= MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_2_mx1w0,
          cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp, and_1249_cse);
      FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_3 <= MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_2_mx1w0,
          cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp, and_1249_cse);
      FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_3 <= MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_2_mx1w0,
          cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp, and_1249_cse);
      FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_3 <= MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_2_mx0w0,
          cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp, and_1249_cse);
      FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_3 <= MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_2_mx1w0,
          cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp, and_1249_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_3 <= 1'b0;
    end
    else if ( core_wen & FpIntToFloat_17U_5U_10U_is_inf_FpIntToFloat_17U_5U_10U_is_inf_or_10_cse
        & (~ (mux_1415_nl)) ) begin
      FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_3 <= MUX_s_1_2_2(FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_2_mx0w0,
          cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp, and_1249_cse);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_1_sva <= 15'b0;
    end
    else if ( cvt_else_and_cse & (~ or_dcpl_386) & (~ mux_tmp_114) ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_1_sva <= IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs <= 1'b0;
      cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs <= 1'b0;
    end
    else if ( FpIntToFloat_17U_5U_10U_if_and_31_cse ) begin
      cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs <= cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
      cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs <= cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs <= 1'b0;
    end
    else if ( cvt_else_and_cse & (~(or_dcpl_15 | nand_171_cse | (cfg_out_precision_1_sva_st_154[0])))
        & (mux_121_nl) ) begin
      cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs <= cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_5_sva <= 15'b0;
    end
    else if ( cvt_else_and_cse & (~ or_dcpl_16) & (~ mux_tmp_122) ) begin
      IntShiftRightSat_49U_6U_17U_o_15_1_5_sva <= IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs <= 1'b0;
      cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs <= 1'b0;
    end
    else if ( FpIntToFloat_17U_5U_10U_if_and_33_cse ) begin
      cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs <= cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
      cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs <= cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs <= 1'b0;
    end
    else if ( cvt_else_and_cse & FpIntToFloat_17U_5U_10U_if_nor_6_cse & (mux_131_nl)
        ) begin
      cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs <= cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs <= 1'b0;
      cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs <= 1'b0;
    end
    else if ( FpIntToFloat_17U_5U_10U_if_and_36_cse ) begin
      cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs <= cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
      cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs <= cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs <= 1'b0;
    end
    else if ( cvt_else_and_cse & FpIntToFloat_17U_5U_10U_if_nor_6_cse & mux_134_cse
        ) begin
      cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs <= cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs <= 1'b0;
    end
    else if ( cvt_else_and_cse & (~ or_tmp_3032) & (mux_143_nl) ) begin
      cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs <= cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs <= 1'b0;
    end
    else if ( cvt_else_and_cse & FpIntToFloat_17U_5U_10U_if_nor_6_cse & (mux_150_nl)
        ) begin
      cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs <= cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_svs <= 1'b0;
    end
    else if ( cvt_else_and_cse & FpIntToFloat_17U_5U_10U_if_nor_10_cse & (mux_153_nl)
        ) begin
      cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_svs <= cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_1_FpMantRNE_24U_11U_else_and_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_612 | (cfg_proc_precision_rsci_d[0]) | (~ cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_itm_8_1)
        | cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1 | (~ cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_itm_8_1)
        | (fsm_output[0]))) ) begin
      cvt_1_FpMantRNE_24U_11U_else_and_svs <= cvt_1_FpMantRNE_24U_11U_else_and_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_2_FpMantRNE_24U_11U_else_and_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_612 | (cfg_proc_precision_rsci_d[0]) | (~ cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1)
        | cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1 | (~ cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1)
        | (fsm_output[0]))) ) begin
      cvt_2_FpMantRNE_24U_11U_else_and_1_svs <= cvt_2_FpMantRNE_24U_11U_else_and_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_3_FpMantRNE_24U_11U_else_and_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_612 | (cfg_proc_precision_rsci_d[0]) | (~ cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1)
        | cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1 | (~ cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1)
        | (fsm_output[0]))) ) begin
      cvt_3_FpMantRNE_24U_11U_else_and_1_svs <= cvt_3_FpMantRNE_24U_11U_else_and_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_4_FpMantRNE_24U_11U_else_and_2_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_612 | (cfg_proc_precision_rsci_d[0]) | (~ cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1)
        | cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1)
        | (fsm_output[0]))) ) begin
      cvt_4_FpMantRNE_24U_11U_else_and_2_svs <= cvt_4_FpMantRNE_24U_11U_else_and_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_5_FpMantRNE_24U_11U_else_and_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_612 | (cfg_proc_precision_rsci_d[0]) | (~ cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1)
        | cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1 | (~ cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1)
        | (fsm_output[0]))) ) begin
      cvt_5_FpMantRNE_24U_11U_else_and_1_svs <= cvt_5_FpMantRNE_24U_11U_else_and_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_6_FpMantRNE_24U_11U_else_and_2_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_612 | (cfg_proc_precision_rsci_d[0]) | (~ cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1)
        | cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1)
        | (fsm_output[0]))) ) begin
      cvt_6_FpMantRNE_24U_11U_else_and_2_svs <= cvt_6_FpMantRNE_24U_11U_else_and_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_7_FpMantRNE_24U_11U_else_and_2_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_612 | (cfg_proc_precision_rsci_d[0]) | (~ cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1)
        | cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1)
        | (fsm_output[0]))) ) begin
      cvt_7_FpMantRNE_24U_11U_else_and_2_svs <= cvt_7_FpMantRNE_24U_11U_else_and_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_8_FpMantRNE_24U_11U_else_and_3_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_612 | (cfg_proc_precision_rsci_d[0]) | (~ cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1)
        | cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 | (~ cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1)
        | (fsm_output[0]))) ) begin
      cvt_8_FpMantRNE_24U_11U_else_and_3_svs <= cvt_8_FpMantRNE_24U_11U_else_and_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_9_FpMantRNE_24U_11U_else_and_1_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_612 | (cfg_proc_precision_rsci_d[0]) | (~ cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1)
        | cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1 | (~ cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1)
        | (fsm_output[0]))) ) begin
      cvt_9_FpMantRNE_24U_11U_else_and_1_svs <= cvt_9_FpMantRNE_24U_11U_else_and_1_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_10_FpMantRNE_24U_11U_else_and_2_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_612 | (cfg_proc_precision_rsci_d[0]) | (~ cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1)
        | cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1)
        | (fsm_output[0]))) ) begin
      cvt_10_FpMantRNE_24U_11U_else_and_2_svs <= cvt_10_FpMantRNE_24U_11U_else_and_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_11_FpMantRNE_24U_11U_else_and_2_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_612 | (cfg_proc_precision_rsci_d[0]) | (~ cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1)
        | cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1)
        | (fsm_output[0]))) ) begin
      cvt_11_FpMantRNE_24U_11U_else_and_2_svs <= cvt_11_FpMantRNE_24U_11U_else_and_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_12_FpMantRNE_24U_11U_else_and_3_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_612 | (cfg_proc_precision_rsci_d[0]) | (~ cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1)
        | cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 | (~ cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1)
        | (fsm_output[0]))) ) begin
      cvt_12_FpMantRNE_24U_11U_else_and_3_svs <= cvt_12_FpMantRNE_24U_11U_else_and_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_13_FpMantRNE_24U_11U_else_and_2_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_612 | (cfg_proc_precision_rsci_d[0]) | (~ cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1)
        | cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1)
        | (fsm_output[0]))) ) begin
      cvt_13_FpMantRNE_24U_11U_else_and_2_svs <= cvt_13_FpMantRNE_24U_11U_else_and_2_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_14_FpMantRNE_24U_11U_else_and_3_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_612 | (cfg_proc_precision_rsci_d[0]) | (~ cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1)
        | cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 | (~ cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1)
        | (fsm_output[0]))) ) begin
      cvt_14_FpMantRNE_24U_11U_else_and_3_svs <= cvt_14_FpMantRNE_24U_11U_else_and_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_15_FpMantRNE_24U_11U_else_and_3_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_612 | (cfg_proc_precision_rsci_d[0]) | (~ cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1)
        | cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 | (~ cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1)
        | (fsm_output[0]))) ) begin
      cvt_15_FpMantRNE_24U_11U_else_and_3_svs <= cvt_15_FpMantRNE_24U_11U_else_and_3_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      cvt_16_FpMantRNE_24U_11U_else_and_4_svs <= 1'b0;
    end
    else if ( core_wen & (~(or_dcpl_612 | (cfg_proc_precision_rsci_d[0]) | (~ cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_itm_8_1)
        | cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_itm_7_1 | (~ cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_itm_8_1)
        | (fsm_output[0]))) ) begin
      cvt_16_FpMantRNE_24U_11U_else_and_4_svs <= cvt_16_FpMantRNE_24U_11U_else_and_4_tmp;
    end
  end
  assign cvt_and_261_nl = (~ FpIntToFloat_17U_5U_10U_is_inf_1_lpi_1_dfm_6) & cvt_asn_323
      & (~ or_tmp_4102);
  assign cvt_and_262_nl = FpIntToFloat_17U_5U_10U_is_inf_1_lpi_1_dfm_6 & cvt_asn_323;
  assign cvt_and_257_nl = (~ FpIntToFloat_17U_5U_10U_is_inf_3_lpi_1_dfm_7) & cvt_asn_323
      & (~ or_5175_tmp);
  assign cvt_and_258_nl = FpIntToFloat_17U_5U_10U_is_inf_3_lpi_1_dfm_7 & cvt_asn_323;
  assign cvt_and_253_nl = (~ FpIntToFloat_17U_5U_10U_is_inf_5_lpi_1_dfm_7) & cvt_asn_323
      & (~ or_5177_tmp);
  assign cvt_and_254_nl = FpIntToFloat_17U_5U_10U_is_inf_5_lpi_1_dfm_7 & cvt_asn_323;
  assign cvt_and_245_nl = (~ FpIntToFloat_17U_5U_10U_is_inf_9_lpi_1_dfm_7) & cvt_asn_323
      & (~ or_5181_tmp);
  assign cvt_and_246_nl = FpIntToFloat_17U_5U_10U_is_inf_9_lpi_1_dfm_7 & cvt_asn_323;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_nl = (reg_FpIntToFloat_17U_5U_10U_o_expo_1_lpi_1_dfm_7_itm
      & (~ IsNaN_5U_10U_land_2_lpi_1_dfm_4)) | FpIntToFloat_17U_5U_10U_is_inf_1_lpi_1_dfm_6;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_1_nl = (reg_FpIntToFloat_17U_5U_10U_o_expo_2_lpi_1_dfm_8_itm
      & (~ IsNaN_5U_10U_land_3_lpi_1_dfm_5)) | FpIntToFloat_17U_5U_10U_is_inf_2_lpi_1_dfm_6;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_2_nl = (reg_FpIntToFloat_17U_5U_10U_o_expo_3_lpi_1_dfm_8_itm
      & (~ IsNaN_5U_10U_land_4_lpi_1_dfm_5)) | FpIntToFloat_17U_5U_10U_is_inf_3_lpi_1_dfm_7;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_3_nl = (reg_FpIntToFloat_17U_5U_10U_o_expo_4_lpi_1_dfm_9_itm
      & (~ IsNaN_5U_10U_land_5_lpi_1_dfm_5)) | FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_7;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_4_nl = (reg_FpIntToFloat_17U_5U_10U_o_expo_5_lpi_1_dfm_8_itm
      & (~ IsNaN_5U_10U_land_6_lpi_1_dfm_5)) | FpIntToFloat_17U_5U_10U_is_inf_5_lpi_1_dfm_7;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_5_nl = (reg_FpIntToFloat_17U_5U_10U_o_expo_6_lpi_1_dfm_9_itm
      & (~ IsNaN_5U_10U_land_7_lpi_1_dfm_6)) | FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_7;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_6_nl = (reg_FpIntToFloat_17U_5U_10U_o_expo_7_lpi_1_dfm_9_itm
      & (~ IsNaN_5U_10U_land_8_lpi_1_dfm_5)) | FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_7;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_7_nl = (reg_FpIntToFloat_17U_5U_10U_o_expo_8_lpi_1_dfm_10_itm
      & (~ IsNaN_5U_10U_land_9_lpi_1_dfm_5)) | FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_8;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_8_nl = (reg_FpIntToFloat_17U_5U_10U_o_expo_9_lpi_1_dfm_8_itm
      & (~ IsNaN_5U_10U_land_lpi_1_dfm_5)) | FpIntToFloat_17U_5U_10U_is_inf_9_lpi_1_dfm_7;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_9_nl = (reg_FpIntToFloat_17U_5U_10U_o_expo_10_lpi_1_dfm_9_itm
      & (~ IsNaN_5U_10U_land_1_lpi_1_dfm_3)) | FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_7;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_10_nl = (reg_FpIntToFloat_17U_5U_10U_o_expo_11_lpi_1_dfm_9_itm
      & (~ IsNaN_5U_10U_land_10_lpi_1_dfm_5)) | FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_7;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_11_nl = (reg_FpIntToFloat_17U_5U_10U_o_expo_12_lpi_1_dfm_10_itm
      & (~ IsNaN_5U_10U_land_11_lpi_1_dfm_5)) | FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_8;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_12_nl = (reg_FpIntToFloat_17U_5U_10U_o_expo_13_lpi_1_dfm_9_itm
      & (~ IsNaN_5U_10U_land_12_lpi_1_dfm_5)) | FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_7;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_13_nl = (reg_FpIntToFloat_17U_5U_10U_o_expo_14_lpi_1_dfm_10_itm
      & (~ IsNaN_5U_10U_land_13_lpi_1_dfm_5)) | FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_8;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_14_nl = (reg_FpIntToFloat_17U_5U_10U_o_expo_15_lpi_1_dfm_10_itm
      & (~ IsNaN_5U_10U_land_14_lpi_1_dfm_6)) | FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_8;
  assign SetToInf_5U_10U_SetToInf_5U_10U_or_15_nl = (reg_FpIntToFloat_17U_5U_10U_o_expo_lpi_1_dfm_11_itm
      & (~ IsNaN_5U_10U_land_15_lpi_1_dfm_3)) | FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_9;
  assign cvt_or_48_nl = cvt_asn_321 | cfg_mode_eql_1_sva_6;
  assign cvt_and_259_nl = (~ FpIntToFloat_17U_5U_10U_is_inf_2_lpi_1_dfm_6) & cvt_asn_329
      & (~ or_5174_tmp);
  assign cvt_and_260_nl = FpIntToFloat_17U_5U_10U_is_inf_2_lpi_1_dfm_6 & cvt_asn_329;
  assign and_3148_nl = cvt_asn_333 & (~ or_5174_tmp);
  assign mux_2301_nl = MUX_s_1_2_2(mux_tmp_2294, (~ or_tmp), cfg_proc_precision_1_sva_st_66[1]);
  assign mux_2302_nl = MUX_s_1_2_2((mux_2301_nl), mux_tmp_2294, cfg_proc_precision_1_sva_st_66[0]);
  assign and_3140_nl = cvt_or_6_cse & (~ or_5176_tmp);
  assign cvt_and_255_nl = (~ FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_7) & cvt_asn_335
      & (~ or_5176_tmp);
  assign cvt_and_256_nl = FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_7 & cvt_asn_335;
  assign mux_2307_nl = MUX_s_1_2_2(mux_tmp_2300, (~ or_tmp_4080), cfg_proc_precision_1_sva_st_66[1]);
  assign mux_2308_nl = MUX_s_1_2_2((mux_2307_nl), mux_tmp_2300, cfg_proc_precision_1_sva_st_66[0]);
  assign cvt_and_251_nl = (~ FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_7) & cvt_asn_353
      & (~ or_5178_tmp);
  assign cvt_and_252_nl = FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_7 & cvt_asn_353;
  assign and_3136_nl = cvt_asn_357 & (~ or_5178_tmp);
  assign mux_2313_nl = MUX_s_1_2_2(mux_tmp_2306, (~ or_tmp_4081), cfg_proc_precision_1_sva_st_90[1]);
  assign mux_2314_nl = MUX_s_1_2_2((mux_2313_nl), mux_tmp_2306, cfg_proc_precision_1_sva_st_90[0]);
  assign cvt_and_249_nl = (~ FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_7) & cvt_asn_365
      & (~ or_5179_tmp);
  assign cvt_and_250_nl = FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_7 & cvt_asn_365;
  assign and_3133_nl = cvt_asn_369 & (~ or_5179_tmp);
  assign mux_2319_nl = MUX_s_1_2_2(mux_tmp_2312, (~ or_tmp_4082), cfg_proc_precision_1_sva_st_102[1]);
  assign mux_2320_nl = MUX_s_1_2_2((mux_2319_nl), mux_tmp_2312, cfg_proc_precision_1_sva_st_102[0]);
  assign and_3128_nl = cvt_or_14_cse & (~ or_5180_tmp);
  assign cvt_and_247_nl = (~ FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_8) & cvt_asn_377
      & (~ or_5180_tmp);
  assign cvt_and_248_nl = FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_8 & cvt_asn_377;
  assign and_3130_nl = cvt_asn_381 & (~ or_5180_tmp);
  assign mux_2326_nl = MUX_s_1_2_2(mux_tmp_2319, (~ or_tmp_4084), cfg_proc_precision_1_sva_st_90[1]);
  assign mux_2327_nl = MUX_s_1_2_2((mux_2326_nl), mux_tmp_2319, cfg_proc_precision_1_sva_st_90[0]);
  assign cvt_and_243_nl = (~ FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_7) & cvt_asn_371
      & (~ or_5182_tmp);
  assign cvt_and_244_nl = FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_7 & cvt_asn_371;
  assign and_3124_nl = cvt_asn_399 & (~ or_5182_tmp);
  assign mux_2331_nl = MUX_s_1_2_2(mux_tmp_2324, (~ or_tmp_4086), cfg_proc_precision_1_sva_st_90[1]);
  assign mux_2332_nl = MUX_s_1_2_2((mux_2331_nl), mux_tmp_2324, cfg_proc_precision_1_sva_st_90[0]);
  assign cvt_and_241_nl = (~ FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_7) & cvt_asn_389
      & (~ or_5183_tmp);
  assign cvt_and_242_nl = FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_7 & cvt_asn_389;
  assign and_3121_nl = cvt_asn_393 & (~ or_5183_tmp);
  assign mux_2337_nl = MUX_s_1_2_2(mux_tmp_2330, (~ or_tmp_4087), cfg_proc_precision_1_sva_st_102[1]);
  assign mux_2338_nl = MUX_s_1_2_2((mux_2337_nl), mux_tmp_2330, cfg_proc_precision_1_sva_st_102[0]);
  assign and_3116_nl = cvt_or_22_cse & (~ or_5184_tmp);
  assign cvt_and_239_nl = (~ FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_8) & cvt_asn_383
      & (~ or_5184_tmp);
  assign cvt_and_240_nl = FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_8 & cvt_asn_383;
  assign and_3118_nl = cvt_asn_387 & (~ or_5184_tmp);
  assign mux_2343_nl = MUX_s_1_2_2(mux_tmp_2336, (~ or_tmp_4084), cfg_proc_precision_1_sva_st_90[1]);
  assign mux_2344_nl = MUX_s_1_2_2((mux_2343_nl), mux_tmp_2336, cfg_proc_precision_1_sva_st_90[0]);
  assign cvt_and_237_nl = (~ FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_7) & cvt_asn_371
      & (~ or_5185_tmp);
  assign cvt_and_238_nl = FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_7 & cvt_asn_371;
  assign and_3115_nl = cvt_asn_375 & (~ or_5185_tmp);
  assign mux_2348_nl = MUX_s_1_2_2(mux_tmp_2341, (~ or_tmp_4092), cfg_proc_precision_1_sva_st_90[1]);
  assign mux_2349_nl = MUX_s_1_2_2((mux_2348_nl), mux_tmp_2341, cfg_proc_precision_1_sva_st_90[0]);
  assign and_3110_nl = cvt_or_26_cse & (~ or_5186_tmp);
  assign cvt_and_235_nl = (~ FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_8) & cvt_asn_359
      & (~ or_5186_tmp);
  assign cvt_and_236_nl = FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_8 & cvt_asn_359;
  assign and_3112_nl = cvt_asn_363 & (~ or_5186_tmp);
  assign and_3104_nl = cvt_or_30_cse & (~ or_5188_tmp);
  assign cvt_and_231_nl = (~ FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_9) & cvt_asn_341
      & (~ or_5188_tmp);
  assign cvt_and_232_nl = FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_9 & cvt_asn_341;
  assign and_3105_nl = cvt_asn_345 & (~ or_5188_tmp);
  assign cvt_and_233_nl = (~ FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_8) & cvt_asn_347
      & (~ or_5187_tmp);
  assign cvt_and_234_nl = FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_8 & cvt_asn_347;
  assign and_3109_nl = cvt_asn_351 & (~ or_5187_tmp);
  assign mux_2360_nl = MUX_s_1_2_2(mux_tmp_2353, (~ or_tmp_4097), cfg_proc_precision_1_sva_st_102[1]);
  assign mux_2361_nl = MUX_s_1_2_2((mux_2360_nl), mux_tmp_2353, cfg_proc_precision_1_sva_st_102[0]);
  assign mux_2362_nl = MUX_s_1_2_2(or_tmp_4097, (~ (mux_2361_nl)), or_5254_cse);
  assign FpFloatToInt_16U_5U_10U_else_mux_2_nl = MUX_s_1_2_2(FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_2,
      cvt_1_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_itm_2,
      chn_idata_data_sva_3_47_31_1[0]);
  assign FpFloatToInt_16U_5U_10U_mux_4_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_else_mux_2_nl),
      cvt_1_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_itm_2,
      cvt_1_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_svs_2);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_nl = (FpFloatToInt_16U_5U_10U_mux_4_nl)
      & (~ IsNaN_5U_10U_land_1_lpi_1_dfm_3);
  assign cvt_if_mux_10_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_nl),
      (reg_chn_idata_data_sva_3_15_0_2_reg[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2281_nl = MUX_s_1_2_2((cvt_if_mux_10_nl), (reg_chn_idata_data_sva_3_15_0_2_reg[0]),
      cfg_mode_eql_1_sva_6);
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_nl = (cvt_8_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_2
      & (~ cvt_1_IntSaturation_17U_8U_else_if_acc_itm_10)) | FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_2;
  assign cvt_else_mux1h_10_nl = MUX1HOT_s_1_3_2((FpIntToFloat_17U_5U_10U_o_mant_1_lpi_1_dfm_1[0]),
      cvt_7_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_2,
      (IntSaturation_17U_8U_IntSaturation_17U_8U_or_nl), {cvt_else_nor_dfs , cvt_else_equal_tmp
      , cvt_else_equal_tmp_1});
  assign cvt_mux_2280_nl = MUX_s_1_2_2((cvt_else_mux1h_10_nl), (reg_chn_idata_data_sva_3_15_0_2_reg[0]),
      cfg_mode_eql_1_sva_6);
  assign cvt_else_mux1h_8_nl = MUX1HOT_s_1_3_2(IntShiftRightSat_49U_6U_17U_o_16_1_sva_4,
      (reg_chn_idata_data_sva_3_15_0_1_reg[4]), (IntSaturation_17U_8U_o_7_1_1_lpi_1_dfm_1[6]),
      {cvt_else_nor_dfs , cvt_else_equal_tmp , cvt_else_equal_tmp_1});
  assign cvt_if_mux_8_nl = MUX_s_1_2_2((reg_chn_idata_data_sva_3_15_0_1_reg[4]),
      (chn_idata_data_sva_3_47_31_1[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2373_nl = MUX_s_1_2_2((cvt_if_mux_8_nl), (cvt_else_mux1h_8_nl),
      cvt_and_tmp_1);
  assign FpFloatToInt_16U_5U_10U_else_mux_5_nl = MUX_s_1_2_2(FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_2,
      cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1,
      chn_idata_data_sva_3_79_63_1[0]);
  assign FpFloatToInt_16U_5U_10U_mux_11_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_else_mux_5_nl),
      cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1,
      cvt_2_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_1_nl = (FpFloatToInt_16U_5U_10U_mux_11_nl)
      & (~ IsNaN_5U_10U_land_2_lpi_1_dfm_4);
  assign cvt_if_mux_25_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_1_nl),
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_1_reg[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2285_nl = MUX_s_1_2_2((cvt_if_mux_25_nl), (chn_idata_data_sva_3_47_31_1[1]),
      cfg_mode_eql_1_sva_6);
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_1_nl = (IntShiftRightSat_49U_6U_17U_o_0_2_sva_3
      & (~ cvt_2_IntSaturation_17U_8U_else_if_acc_1_itm_10)) | FpFloatToInt_16U_5U_10U_internal_int_0_2_sva_2;
  assign cvt_else_mux1h_29_nl = MUX1HOT_s_1_3_2((FpIntToFloat_17U_5U_10U_o_mant_2_lpi_1_dfm_1[0]),
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_1_itm_3, (IntSaturation_17U_8U_IntSaturation_17U_8U_or_1_nl),
      {cvt_else_nor_dfs_1_mx1 , cvt_else_equal_tmp_3_mx0 , cvt_else_equal_tmp_4_mx1});
  assign cvt_mux_2284_nl = MUX_s_1_2_2((cvt_else_mux1h_29_nl), (chn_idata_data_sva_3_47_31_1[1]),
      cfg_mode_eql_1_sva_6);
  assign cvt_else_mux1h_27_nl = MUX1HOT_s_1_3_2(IntShiftRightSat_49U_6U_17U_o_16_2_sva_3,
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_reg[4]), (IntSaturation_17U_8U_o_7_1_2_lpi_1_dfm_1[6]),
      {cvt_else_nor_dfs_1_mx1 , cvt_else_equal_tmp_3_mx0 , cvt_else_equal_tmp_4_mx1});
  assign cvt_if_mux_23_nl = MUX_s_1_2_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_reg[4]),
      (chn_idata_data_sva_3_79_63_1[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2346_nl = MUX_s_1_2_2((cvt_if_mux_23_nl), (cvt_else_mux1h_27_nl),
      cvt_and_tmp_1);
  assign FpFloatToInt_16U_5U_10U_else_mux_8_nl = MUX_s_1_2_2(FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_2,
      cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1,
      chn_idata_data_sva_3_111_95_1[0]);
  assign FpFloatToInt_16U_5U_10U_mux_18_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_else_mux_8_nl),
      cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1,
      cvt_3_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_2_nl = (FpFloatToInt_16U_5U_10U_mux_18_nl)
      & (~ IsNaN_5U_10U_land_3_lpi_1_dfm_5);
  assign cvt_if_mux_40_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_2_nl),
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_1_reg[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2289_nl = MUX_s_1_2_2((cvt_if_mux_40_nl), (chn_idata_data_sva_3_79_63_1[1]),
      cfg_mode_eql_1_sva_6);
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_2_nl = (IntShiftRightSat_49U_6U_17U_o_0_3_sva_4
      & (~ cvt_3_IntSaturation_17U_8U_else_if_acc_1_itm_10)) | FpFloatToInt_16U_5U_10U_internal_int_0_3_sva_2;
  assign cvt_else_mux1h_48_nl = MUX1HOT_s_1_3_2((FpIntToFloat_17U_5U_10U_o_mant_3_lpi_1_dfm_1[0]),
      cvt_15_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_2,
      (IntSaturation_17U_8U_IntSaturation_17U_8U_or_2_nl), {cvt_else_nor_dfs , cvt_else_equal_tmp
      , cvt_else_equal_tmp_1});
  assign cvt_mux_2288_nl = MUX_s_1_2_2((cvt_else_mux1h_48_nl), (chn_idata_data_sva_3_79_63_1[1]),
      cfg_mode_eql_1_sva_6);
  assign cvt_else_mux1h_46_nl = MUX1HOT_s_1_3_2(IntShiftRightSat_49U_6U_17U_o_16_3_sva_4,
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_reg[4]), (IntSaturation_17U_8U_o_7_1_3_lpi_1_dfm_1[6]),
      {cvt_else_nor_dfs , cvt_else_equal_tmp , cvt_else_equal_tmp_1});
  assign cvt_if_mux_38_nl = MUX_s_1_2_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_reg[4]),
      (chn_idata_data_sva_3_111_95_1[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2348_nl = MUX_s_1_2_2((cvt_if_mux_38_nl), (cvt_else_mux1h_46_nl),
      cvt_and_tmp_1);
  assign FpFloatToInt_16U_5U_10U_else_mux_11_nl = MUX_s_1_2_2(FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_2,
      cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1,
      chn_idata_data_sva_3_143_127_1[0]);
  assign FpFloatToInt_16U_5U_10U_mux_25_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_else_mux_11_nl),
      cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1,
      cvt_4_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_3_nl = (FpFloatToInt_16U_5U_10U_mux_25_nl)
      & (~ IsNaN_5U_10U_land_4_lpi_1_dfm_5);
  assign cvt_if_mux_55_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_3_nl),
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_1_reg[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2293_nl = MUX_s_1_2_2((cvt_if_mux_55_nl), (chn_idata_data_sva_3_111_95_1[1]),
      cfg_mode_eql_1_sva_6);
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_3_nl = (IntShiftRightSat_49U_6U_17U_o_0_4_sva_3
      & (~ cvt_4_IntSaturation_17U_8U_else_if_acc_2_itm_10)) | FpFloatToInt_16U_5U_10U_internal_int_0_4_sva_2;
  assign cvt_else_mux1h_67_nl = MUX1HOT_s_1_3_2((FpIntToFloat_17U_5U_10U_o_mant_4_lpi_1_dfm_1[0]),
      cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1,
      (IntSaturation_17U_8U_IntSaturation_17U_8U_or_3_nl), {cvt_else_nor_dfs_3_mx1
      , cvt_else_equal_tmp_9_mx1 , cvt_else_equal_tmp_10_mx0});
  assign cvt_mux_2292_nl = MUX_s_1_2_2((cvt_else_mux1h_67_nl), (chn_idata_data_sva_3_111_95_1[1]),
      cfg_mode_eql_1_sva_6);
  assign cvt_else_mux1h_65_nl = MUX1HOT_s_1_3_2(IntShiftRightSat_49U_6U_17U_o_16_4_sva_3,
      (FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5[14]), (IntSaturation_17U_8U_o_7_1_4_lpi_1_dfm_1[6]),
      {cvt_else_nor_dfs_3_mx1 , cvt_else_equal_tmp_9_mx1 , cvt_else_equal_tmp_10_mx0});
  assign cvt_if_mux_53_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_o_int_15_1_4_lpi_1_dfm_5[14]),
      (chn_idata_data_sva_3_143_127_1[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2350_nl = MUX_s_1_2_2((cvt_if_mux_53_nl), (cvt_else_mux1h_65_nl),
      cvt_and_tmp_1);
  assign FpFloatToInt_16U_5U_10U_else_mux_14_nl = MUX_s_1_2_2(FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_2,
      cvt_5_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_2,
      chn_idata_data_sva_3_175_159_1[0]);
  assign FpFloatToInt_16U_5U_10U_mux_32_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_else_mux_14_nl),
      cvt_5_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_2,
      cvt_5_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_4_nl = (FpFloatToInt_16U_5U_10U_mux_32_nl)
      & (~ IsNaN_5U_10U_land_5_lpi_1_dfm_5);
  assign cvt_if_mux_70_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_4_nl),
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_1_reg[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2297_nl = MUX_s_1_2_2((cvt_if_mux_70_nl), (chn_idata_data_sva_3_143_127_1[1]),
      cfg_mode_eql_1_sva_6);
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_4_nl = (IntShiftRightSat_49U_6U_17U_o_0_5_sva_4
      & (~ cvt_5_IntSaturation_17U_8U_else_if_acc_1_itm_10)) | FpFloatToInt_16U_5U_10U_internal_int_0_5_sva_2;
  assign cvt_else_mux1h_86_nl = MUX1HOT_s_1_3_2((FpIntToFloat_17U_5U_10U_o_mant_5_lpi_1_dfm_1[0]),
      cvt_1_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_itm_2,
      (IntSaturation_17U_8U_IntSaturation_17U_8U_or_4_nl), {cvt_else_nor_dfs , cvt_else_equal_tmp
      , cvt_else_equal_tmp_1});
  assign cvt_mux_2296_nl = MUX_s_1_2_2((cvt_else_mux1h_86_nl), (chn_idata_data_sva_3_143_127_1[1]),
      cfg_mode_eql_1_sva_6);
  assign cvt_else_mux1h_84_nl = MUX1HOT_s_1_3_2(IntShiftRightSat_49U_6U_17U_o_16_5_sva_4,
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_reg[4]), (IntSaturation_17U_8U_o_7_1_5_lpi_1_dfm_1[6]),
      {cvt_else_nor_dfs , cvt_else_equal_tmp , cvt_else_equal_tmp_1});
  assign cvt_if_mux_68_nl = MUX_s_1_2_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_reg[4]),
      (chn_idata_data_sva_3_175_159_1[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2352_nl = MUX_s_1_2_2((cvt_if_mux_68_nl), (cvt_else_mux1h_84_nl),
      cvt_and_tmp_1);
  assign FpFloatToInt_16U_5U_10U_else_mux_17_nl = MUX_s_1_2_2(FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_2,
      cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1,
      chn_idata_data_sva_3_207_191_1[0]);
  assign FpFloatToInt_16U_5U_10U_mux_39_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_else_mux_17_nl),
      cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1,
      cvt_6_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_5_nl = (FpFloatToInt_16U_5U_10U_mux_39_nl)
      & (~ IsNaN_5U_10U_land_6_lpi_1_dfm_5);
  assign cvt_if_mux_85_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_5_nl),
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_2_lpi_1_dfm_5_1_reg[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2301_nl = MUX_s_1_2_2((cvt_if_mux_85_nl), (chn_idata_data_sva_3_175_159_1[1]),
      cfg_mode_eql_1_sva_6);
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_5_nl = (IntShiftRightSat_49U_6U_17U_o_0_6_sva_3
      & (~ cvt_6_IntSaturation_17U_8U_else_if_acc_2_itm_10)) | FpFloatToInt_16U_5U_10U_internal_int_0_6_sva_2;
  assign cvt_else_mux1h_105_nl = MUX1HOT_s_1_3_2((FpIntToFloat_17U_5U_10U_o_mant_6_lpi_1_dfm_1[0]),
      cvt_2_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1,
      (IntSaturation_17U_8U_IntSaturation_17U_8U_or_5_nl), {cvt_else_nor_dfs_5_mx1
      , cvt_else_equal_tmp_15_mx0 , cvt_else_equal_tmp_16_mx1});
  assign cvt_mux_2300_nl = MUX_s_1_2_2((cvt_else_mux1h_105_nl), (chn_idata_data_sva_3_175_159_1[1]),
      cfg_mode_eql_1_sva_6);
  assign cvt_else_mux1h_103_nl = MUX1HOT_s_1_3_2(IntShiftRightSat_49U_6U_17U_o_16_6_sva_3,
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_reg[4]), (IntSaturation_17U_8U_o_7_1_6_lpi_1_dfm_1[6]),
      {cvt_else_nor_dfs_5_mx1 , cvt_else_equal_tmp_15_mx0 , cvt_else_equal_tmp_16_mx1});
  assign cvt_if_mux_83_nl = MUX_s_1_2_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_reg[4]),
      (chn_idata_data_sva_3_207_191_1[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2354_nl = MUX_s_1_2_2((cvt_if_mux_83_nl), (cvt_else_mux1h_103_nl),
      cvt_and_tmp_1);
  assign FpFloatToInt_16U_5U_10U_else_mux_20_nl = MUX_s_1_2_2(FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_2,
      cvt_7_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_2,
      chn_idata_data_sva_3_239_223_1[0]);
  assign FpFloatToInt_16U_5U_10U_mux_46_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_else_mux_20_nl),
      cvt_7_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_2,
      cvt_7_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_6_nl = (FpFloatToInt_16U_5U_10U_mux_46_nl)
      & (~ IsNaN_5U_10U_land_7_lpi_1_dfm_6);
  assign cvt_if_mux_100_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_6_nl),
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_1_reg[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2305_nl = MUX_s_1_2_2((cvt_if_mux_100_nl), (chn_idata_data_sva_3_207_191_1[1]),
      cfg_mode_eql_1_sva_6);
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_6_nl = (IntShiftRightSat_49U_6U_17U_o_0_7_sva_3
      & (~ cvt_7_IntSaturation_17U_8U_else_if_acc_2_itm_10)) | FpFloatToInt_16U_5U_10U_internal_int_0_7_sva_2;
  assign cvt_else_mux1h_124_nl = MUX1HOT_s_1_3_2((FpIntToFloat_17U_5U_10U_o_mant_7_lpi_1_dfm_1[0]),
      cvt_3_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1,
      (IntSaturation_17U_8U_IntSaturation_17U_8U_or_6_nl), {cvt_else_nor_dfs_6_mx1
      , cvt_else_equal_tmp_18_mx0 , cvt_else_equal_tmp_19_mx0});
  assign cvt_mux_2304_nl = MUX_s_1_2_2((cvt_else_mux1h_124_nl), (chn_idata_data_sva_3_207_191_1[1]),
      cfg_mode_eql_1_sva_6);
  assign cvt_else_mux1h_122_nl = MUX1HOT_s_1_3_2(IntShiftRightSat_49U_6U_17U_o_16_7_sva_3,
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_reg[4]), (IntSaturation_17U_8U_o_7_1_7_lpi_1_dfm_1[6]),
      {cvt_else_nor_dfs_6_mx1 , cvt_else_equal_tmp_18_mx0 , cvt_else_equal_tmp_19_mx0});
  assign cvt_if_mux_98_nl = MUX_s_1_2_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_reg[4]),
      (chn_idata_data_sva_3_239_223_1[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2358_nl = MUX_s_1_2_2((cvt_if_mux_98_nl), (cvt_else_mux1h_122_nl),
      cvt_and_tmp_1);
  assign FpFloatToInt_16U_5U_10U_else_mux_23_nl = MUX_s_1_2_2(FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_2,
      cvt_8_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_2,
      chn_idata_data_sva_3_271_255_1[0]);
  assign FpFloatToInt_16U_5U_10U_mux_53_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_else_mux_23_nl),
      cvt_8_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_2,
      cvt_8_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_7_nl = (FpFloatToInt_16U_5U_10U_mux_53_nl)
      & (~ IsNaN_5U_10U_land_8_lpi_1_dfm_5);
  assign cvt_if_mux_115_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_7_nl),
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_1_reg[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2309_nl = MUX_s_1_2_2((cvt_if_mux_115_nl), (chn_idata_data_sva_3_239_223_1[1]),
      cfg_mode_eql_1_sva_6);
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_7_nl = (IntShiftRightSat_49U_6U_17U_o_0_8_sva_3
      & (~ cvt_8_IntSaturation_17U_8U_else_if_acc_3_itm_10)) | FpFloatToInt_16U_5U_10U_internal_int_0_8_sva_2;
  assign cvt_else_mux1h_143_nl = MUX1HOT_s_1_3_2((FpIntToFloat_17U_5U_10U_o_mant_8_lpi_1_dfm_1[0]),
      cvt_4_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1,
      (IntSaturation_17U_8U_IntSaturation_17U_8U_or_7_nl), {cvt_else_nor_dfs_7_mx1
      , cvt_else_equal_tmp_21_mx1 , cvt_else_equal_tmp_22_mx1});
  assign cvt_mux_2308_nl = MUX_s_1_2_2((cvt_else_mux1h_143_nl), (chn_idata_data_sva_3_239_223_1[1]),
      cfg_mode_eql_1_sva_6);
  assign cvt_else_mux1h_141_nl = MUX1HOT_s_1_3_2(IntShiftRightSat_49U_6U_17U_o_16_8_sva_3,
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_reg[4]), (IntSaturation_17U_8U_o_7_1_8_lpi_1_dfm_1[6]),
      {cvt_else_nor_dfs_7_mx1 , cvt_else_equal_tmp_21_mx1 , cvt_else_equal_tmp_22_mx1});
  assign cvt_if_mux_113_nl = MUX_s_1_2_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_reg[4]),
      (chn_idata_data_sva_3_271_255_1[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2360_nl = MUX_s_1_2_2((cvt_if_mux_113_nl), (cvt_else_mux1h_141_nl),
      cvt_and_tmp_1);
  assign FpFloatToInt_16U_5U_10U_else_mux_26_nl = MUX_s_1_2_2(FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_2,
      cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1,
      chn_idata_data_sva_3_303_287_1[0]);
  assign FpFloatToInt_16U_5U_10U_mux_60_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_else_mux_26_nl),
      cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1,
      cvt_9_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_8_nl = (FpFloatToInt_16U_5U_10U_mux_60_nl)
      & (~ IsNaN_5U_10U_land_9_lpi_1_dfm_5);
  assign cvt_if_mux_130_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_8_nl),
      (FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_7_itm_1[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2313_nl = MUX_s_1_2_2((cvt_if_mux_130_nl), (chn_idata_data_sva_3_271_255_1[1]),
      cfg_mode_eql_1_sva_6);
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_8_nl = (IntShiftRightSat_49U_6U_17U_o_0_9_sva_4
      & (~ cvt_9_IntSaturation_17U_8U_else_if_acc_1_itm_10)) | FpFloatToInt_16U_5U_10U_internal_int_0_9_sva_2;
  assign cvt_else_mux1h_162_nl = MUX1HOT_s_1_3_2((FpIntToFloat_17U_5U_10U_o_mant_9_lpi_1_dfm_1[0]),
      cvt_5_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_2,
      (IntSaturation_17U_8U_IntSaturation_17U_8U_or_8_nl), {cvt_else_nor_dfs , cvt_else_equal_tmp
      , cvt_else_equal_tmp_1});
  assign cvt_mux_2312_nl = MUX_s_1_2_2((cvt_else_mux1h_162_nl), (chn_idata_data_sva_3_271_255_1[1]),
      cfg_mode_eql_1_sva_6);
  assign cvt_else_mux1h_160_nl = MUX1HOT_s_1_3_2(IntShiftRightSat_49U_6U_17U_o_16_9_sva_4,
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_reg[4]), (IntSaturation_17U_8U_o_7_1_9_lpi_1_dfm_1[6]),
      {cvt_else_nor_dfs , cvt_else_equal_tmp , cvt_else_equal_tmp_1});
  assign cvt_if_mux_128_nl = MUX_s_1_2_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_reg[4]),
      (chn_idata_data_sva_3_303_287_1[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2362_nl = MUX_s_1_2_2((cvt_if_mux_128_nl), (cvt_else_mux1h_160_nl),
      cvt_and_tmp_1);
  assign FpFloatToInt_16U_5U_10U_else_mux_29_nl = MUX_s_1_2_2(FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_2,
      cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1,
      chn_idata_data_sva_3_335_319_1[0]);
  assign FpFloatToInt_16U_5U_10U_mux_67_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_else_mux_29_nl),
      cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1,
      cvt_10_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_9_nl = (FpFloatToInt_16U_5U_10U_mux_67_nl)
      & (~ IsNaN_5U_10U_land_10_lpi_1_dfm_5);
  assign cvt_if_mux_145_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_9_nl),
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_3_lpi_1_dfm_5_1_reg[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2317_nl = MUX_s_1_2_2((cvt_if_mux_145_nl), (chn_idata_data_sva_3_303_287_1[1]),
      cfg_mode_eql_1_sva_6);
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_9_nl = (cvt_9_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_1_itm_1
      & (~ cvt_10_IntSaturation_17U_8U_else_if_acc_2_itm_10)) | FpFloatToInt_16U_5U_10U_internal_int_0_1_sva_2;
  assign cvt_else_mux1h_181_nl = MUX1HOT_s_1_3_2((FpIntToFloat_17U_5U_10U_o_mant_10_lpi_1_dfm_1[0]),
      cvt_6_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1,
      (IntSaturation_17U_8U_IntSaturation_17U_8U_or_9_nl), {cvt_else_nor_dfs_9_mx1
      , cvt_else_equal_tmp_27_mx0 , cvt_else_equal_tmp_28_mx1});
  assign cvt_mux_2316_nl = MUX_s_1_2_2((cvt_else_mux1h_181_nl), (chn_idata_data_sva_3_303_287_1[1]),
      cfg_mode_eql_1_sva_6);
  assign cvt_else_mux1h_179_nl = MUX1HOT_s_1_3_2(IntShiftRightSat_49U_6U_17U_o_16_10_sva_3,
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_reg[4]), (IntSaturation_17U_8U_o_7_1_10_lpi_1_dfm_1[6]),
      {cvt_else_nor_dfs_9_mx1 , cvt_else_equal_tmp_27_mx0 , cvt_else_equal_tmp_28_mx1});
  assign cvt_if_mux_143_nl = MUX_s_1_2_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_10_lpi_1_dfm_5_reg[4]),
      (chn_idata_data_sva_3_335_319_1[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2364_nl = MUX_s_1_2_2((cvt_if_mux_143_nl), (cvt_else_mux1h_179_nl),
      cvt_and_tmp_1);
  assign FpFloatToInt_16U_5U_10U_else_mux_32_nl = MUX_s_1_2_2(FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_2,
      cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1,
      chn_idata_data_sva_3_367_351_1[0]);
  assign FpFloatToInt_16U_5U_10U_mux_74_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_else_mux_32_nl),
      cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1,
      cvt_11_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_10_nl = (FpFloatToInt_16U_5U_10U_mux_74_nl)
      & (~ IsNaN_5U_10U_land_11_lpi_1_dfm_5);
  assign cvt_if_mux_160_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_10_nl),
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_5_lpi_1_dfm_5_1_reg[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2321_nl = MUX_s_1_2_2((cvt_if_mux_160_nl), (chn_idata_data_sva_3_335_319_1[1]),
      cfg_mode_eql_1_sva_6);
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_10_nl = (IntShiftRightSat_49U_6U_17U_o_0_11_sva_3
      & (~ cvt_11_IntSaturation_17U_8U_else_if_acc_2_itm_10)) | FpFloatToInt_16U_5U_10U_internal_int_0_10_sva_2;
  assign cvt_else_mux1h_200_nl = MUX1HOT_s_1_3_2((FpIntToFloat_17U_5U_10U_o_mant_11_lpi_1_dfm_1[0]),
      cvt_10_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1,
      (IntSaturation_17U_8U_IntSaturation_17U_8U_or_10_nl), {cvt_else_nor_dfs_10_mx1
      , cvt_else_equal_tmp_30_mx0 , cvt_else_equal_tmp_31_mx0});
  assign cvt_mux_2320_nl = MUX_s_1_2_2((cvt_else_mux1h_200_nl), (chn_idata_data_sva_3_335_319_1[1]),
      cfg_mode_eql_1_sva_6);
  assign cvt_else_mux1h_198_nl = MUX1HOT_s_1_3_2(IntShiftRightSat_49U_6U_17U_o_16_11_sva_3,
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_reg[4]), (IntSaturation_17U_8U_o_7_1_11_lpi_1_dfm_1[6]),
      {cvt_else_nor_dfs_10_mx1 , cvt_else_equal_tmp_30_mx0 , cvt_else_equal_tmp_31_mx0});
  assign cvt_if_mux_158_nl = MUX_s_1_2_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_11_lpi_1_dfm_5_reg[4]),
      (chn_idata_data_sva_3_367_351_1[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2366_nl = MUX_s_1_2_2((cvt_if_mux_158_nl), (cvt_else_mux1h_198_nl),
      cvt_and_tmp_1);
  assign FpFloatToInt_16U_5U_10U_else_mux_35_nl = MUX_s_1_2_2(FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_2,
      cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1,
      chn_idata_data_sva_3_399_383_1[0]);
  assign FpFloatToInt_16U_5U_10U_mux_81_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_else_mux_35_nl),
      cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1,
      cvt_12_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_11_nl = (FpFloatToInt_16U_5U_10U_mux_81_nl)
      & (~ IsNaN_5U_10U_land_12_lpi_1_dfm_5);
  assign cvt_if_mux_175_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_11_nl),
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_6_lpi_1_dfm_5_1_reg[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2325_nl = MUX_s_1_2_2((cvt_if_mux_175_nl), (chn_idata_data_sva_3_367_351_1[1]),
      cfg_mode_eql_1_sva_6);
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_11_nl = (IntShiftRightSat_49U_6U_17U_o_0_12_sva_3
      & (~ cvt_12_IntSaturation_17U_8U_else_if_acc_3_itm_10)) | FpFloatToInt_16U_5U_10U_internal_int_0_11_sva_2;
  assign cvt_else_mux1h_219_nl = MUX1HOT_s_1_3_2((FpIntToFloat_17U_5U_10U_o_mant_12_lpi_1_dfm_1[0]),
      cvt_11_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1,
      (IntSaturation_17U_8U_IntSaturation_17U_8U_or_11_nl), {cvt_else_nor_dfs_11_mx1
      , cvt_else_equal_tmp_33_mx1 , cvt_else_equal_tmp_34_mx1});
  assign cvt_mux_2324_nl = MUX_s_1_2_2((cvt_else_mux1h_219_nl), (chn_idata_data_sva_3_367_351_1[1]),
      cfg_mode_eql_1_sva_6);
  assign cvt_else_mux1h_217_nl = MUX1HOT_s_1_3_2(IntShiftRightSat_49U_6U_17U_o_16_12_sva_3,
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_reg[4]), (IntSaturation_17U_8U_o_7_1_12_lpi_1_dfm_1[6]),
      {cvt_else_nor_dfs_11_mx1 , cvt_else_equal_tmp_33_mx1 , cvt_else_equal_tmp_34_mx1});
  assign cvt_if_mux_173_nl = MUX_s_1_2_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_12_lpi_1_dfm_5_reg[4]),
      (chn_idata_data_sva_3_399_383_1[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2370_nl = MUX_s_1_2_2((cvt_if_mux_173_nl), (cvt_else_mux1h_217_nl),
      cvt_and_tmp_1);
  assign FpFloatToInt_16U_5U_10U_else_mux_38_nl = MUX_s_1_2_2(FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_2,
      cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1,
      chn_idata_data_sva_3_431_415_1[0]);
  assign FpFloatToInt_16U_5U_10U_mux_88_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_else_mux_38_nl),
      cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1,
      cvt_13_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_12_nl = (FpFloatToInt_16U_5U_10U_mux_88_nl)
      & (~ IsNaN_5U_10U_land_13_lpi_1_dfm_5);
  assign cvt_if_mux_190_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_12_nl),
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_7_lpi_1_dfm_5_1_reg[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2329_nl = MUX_s_1_2_2((cvt_if_mux_190_nl), (chn_idata_data_sva_3_399_383_1[1]),
      cfg_mode_eql_1_sva_6);
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_12_nl = (IntShiftRightSat_49U_6U_17U_o_0_13_sva_3
      & (~ cvt_13_IntSaturation_17U_8U_else_if_acc_2_itm_10)) | FpFloatToInt_16U_5U_10U_internal_int_0_12_sva_2;
  assign cvt_else_mux1h_238_nl = MUX1HOT_s_1_3_2((FpIntToFloat_17U_5U_10U_o_mant_13_lpi_1_dfm_1[0]),
      cvt_12_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1,
      (IntSaturation_17U_8U_IntSaturation_17U_8U_or_12_nl), {cvt_else_nor_dfs_9_mx1
      , cvt_else_equal_tmp_36_mx0 , cvt_else_equal_tmp_37_mx0});
  assign cvt_mux_2328_nl = MUX_s_1_2_2((cvt_else_mux1h_238_nl), (chn_idata_data_sva_3_399_383_1[1]),
      cfg_mode_eql_1_sva_6);
  assign cvt_else_mux1h_236_nl = MUX1HOT_s_1_3_2(IntShiftRightSat_49U_6U_17U_o_16_13_sva_3,
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_reg[4]), (IntSaturation_17U_8U_o_7_1_13_lpi_1_dfm_1[6]),
      {cvt_else_nor_dfs_9_mx1 , cvt_else_equal_tmp_36_mx0 , cvt_else_equal_tmp_37_mx0});
  assign cvt_if_mux_188_nl = MUX_s_1_2_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_13_lpi_1_dfm_5_reg[4]),
      (chn_idata_data_sva_3_431_415_1[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2372_nl = MUX_s_1_2_2((cvt_if_mux_188_nl), (cvt_else_mux1h_236_nl),
      cvt_and_tmp_1);
  assign FpFloatToInt_16U_5U_10U_else_mux_41_nl = MUX_s_1_2_2(FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_2,
      cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1,
      chn_idata_data_sva_3_463_447_1[0]);
  assign FpFloatToInt_16U_5U_10U_mux_95_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_else_mux_41_nl),
      cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1,
      cvt_14_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_13_nl = (FpFloatToInt_16U_5U_10U_mux_95_nl)
      & (~ IsNaN_5U_10U_land_14_lpi_1_dfm_6);
  assign cvt_if_mux_205_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_13_nl),
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_8_lpi_1_dfm_5_1_reg[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2333_nl = MUX_s_1_2_2((cvt_if_mux_205_nl), (chn_idata_data_sva_3_431_415_1[1]),
      cfg_mode_eql_1_sva_6);
  assign chn_odata_data_mux_1_nl = MUX_s_1_2_2(chn_odata_data_13_0_lpi_1_dfm_1_mx0w0,
      chn_odata_data_13_0_lpi_1_dfm_1, or_dcpl_195);
  assign cvt_mux_2332_nl = MUX_s_1_2_2((chn_odata_data_mux_1_nl), (chn_idata_data_sva_3_431_415_1[1]),
      cfg_mode_eql_1_sva_6);
  assign cvt_else_mux1h_255_nl = MUX1HOT_s_1_3_2(IntShiftRightSat_49U_6U_17U_o_16_14_sva_3,
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_reg[4]), (IntSaturation_17U_8U_o_7_1_14_lpi_1_dfm_1[6]),
      {cvt_else_nor_dfs_13_mx1 , cvt_else_equal_tmp_39_mx1 , cvt_else_equal_tmp_40_mx1});
  assign cvt_if_mux_203_nl = MUX_s_1_2_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_reg[4]),
      (chn_idata_data_sva_3_463_447_1[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2368_nl = MUX_s_1_2_2((cvt_if_mux_203_nl), (cvt_else_mux1h_255_nl),
      cvt_and_tmp_1);
  assign FpFloatToInt_16U_5U_10U_else_mux_44_nl = MUX_s_1_2_2(FpFloatToInt_16U_5U_10U_internal_int_0_15_sva_2,
      cvt_15_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_2,
      chn_idata_data_sva_3_495_479_1[0]);
  assign FpFloatToInt_16U_5U_10U_mux_102_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_else_mux_44_nl),
      cvt_15_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_2,
      cvt_15_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_14_nl = (FpFloatToInt_16U_5U_10U_mux_102_nl)
      & (~ IsNaN_5U_10U_land_15_lpi_1_dfm_3);
  assign cvt_if_mux_220_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_14_nl),
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_9_lpi_1_dfm_5_1_reg[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2337_nl = MUX_s_1_2_2((cvt_if_mux_220_nl), (chn_idata_data_sva_3_463_447_1[1]),
      cfg_mode_eql_1_sva_6);
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_14_nl = (IntShiftRightSat_49U_6U_17U_o_0_15_sva_3
      & (~ cvt_15_IntSaturation_17U_8U_else_if_acc_3_itm_10)) | FpFloatToInt_16U_5U_10U_internal_int_0_13_sva_2;
  assign cvt_else_mux1h_276_nl = MUX1HOT_s_1_3_2((FpIntToFloat_17U_5U_10U_o_mant_15_lpi_1_dfm_1[0]),
      cvt_13_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_2_itm_1,
      (IntSaturation_17U_8U_IntSaturation_17U_8U_or_14_nl), {cvt_else_nor_dfs_14_mx1
      , cvt_else_equal_tmp_42_mx0 , cvt_else_equal_tmp_43_mx0});
  assign cvt_mux_2336_nl = MUX_s_1_2_2((cvt_else_mux1h_276_nl), (chn_idata_data_sva_3_463_447_1[1]),
      cfg_mode_eql_1_sva_6);
  assign cvt_else_mux1h_274_nl = MUX1HOT_s_1_3_2(IntShiftRightSat_49U_6U_17U_o_16_15_sva_3,
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_reg[4]), (IntSaturation_17U_8U_o_7_1_15_lpi_1_dfm_1[6]),
      {cvt_else_nor_dfs_14_mx1 , cvt_else_equal_tmp_42_mx0 , cvt_else_equal_tmp_43_mx0});
  assign cvt_if_mux_218_nl = MUX_s_1_2_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_15_lpi_1_dfm_5_reg[4]),
      (chn_idata_data_sva_3_495_479_1[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2356_nl = MUX_s_1_2_2((cvt_if_mux_218_nl), (cvt_else_mux1h_274_nl),
      cvt_and_tmp_1);
  assign IntSaturation_17U_8U_IntSaturation_17U_8U_or_15_nl = (IntShiftRightSat_49U_6U_17U_o_0_sva_3
      & (~ cvt_16_IntSaturation_17U_8U_else_if_acc_4_itm_10)) | FpFloatToInt_16U_5U_10U_internal_int_0_14_sva_2;
  assign cvt_else_mux1h_295_nl = MUX1HOT_s_1_3_2((FpIntToFloat_17U_5U_10U_o_mant_lpi_1_dfm_1[0]),
      cvt_14_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_3_itm_1,
      (IntSaturation_17U_8U_IntSaturation_17U_8U_or_15_nl), {cvt_else_nor_dfs_15_mx1
      , cvt_else_equal_tmp_45_mx1 , cvt_else_equal_tmp_46_mx1});
  assign FpFloatToInt_16U_5U_10U_else_mux_47_nl = MUX_s_1_2_2(FpFloatToInt_16U_5U_10U_internal_int_0_sva_3,
      cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1,
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_1_itm_3);
  assign FpFloatToInt_16U_5U_10U_mux_109_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_else_mux_47_nl),
      cvt_16_FpFloatToInt_16U_5U_10U_else_if_slc_FpFloatToInt_16U_5U_10U_else_if_ac_int_cctor_0_4_itm_1,
      cvt_16_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_4_svs_2);
  assign FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_15_nl = (FpFloatToInt_16U_5U_10U_mux_109_nl)
      & (~ IsNaN_5U_10U_land_lpi_1_dfm_5);
  assign cvt_if_mux_235_nl = MUX_s_1_2_2((FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_and_15_nl),
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_14_lpi_1_dfm_5_1_reg[0]), cvt_if_unequal_tmp);
  assign cvt_mux_2340_nl = MUX_s_1_2_2((cvt_if_mux_235_nl), (cvt_else_mux1h_295_nl),
      cvt_unequal_tmp_21);
  assign cvt_else_mux1h_292_nl = MUX1HOT_s_1_3_2(IntShiftRightSat_49U_6U_17U_o_16_sva_3,
      (reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_reg[4]), (IntSaturation_17U_8U_o_7_1_lpi_1_dfm_1[6]),
      {cvt_else_nor_dfs_15_mx1 , cvt_else_equal_tmp_45_mx1 , cvt_else_equal_tmp_46_mx1});
  assign cvt_if_mux_232_nl = MUX_s_1_2_2((reg_FpFloatToInt_16U_5U_10U_o_int_15_1_lpi_1_dfm_5_reg[4]),
      IntSaturation_17U_16U_IntSaturation_17U_16U_or_1_itm_3, cvt_if_unequal_tmp);
  assign cvt_mux_2341_nl = MUX_s_1_2_2((cvt_if_mux_232_nl), (cvt_else_mux1h_292_nl),
      cvt_unequal_tmp_21);
  assign nor_2081_nl = ~(cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_itm_8_1
      | cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1 | (~ cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt));
  assign nor_2082_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | (~ cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_st_2
      | cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_2);
  assign mux_nl = MUX_s_1_2_2((nor_2082_nl), (nor_2081_nl), or_5189_cse);
  assign or_9_nl = (~((cfg_proc_precision_rsci_d!=2'b10))) | cfg_mode_eql_rsci_d;
  assign or_11_nl = (~((cvt_1_FpMantRNE_24U_11U_else_and_tmp & cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_itm_8_1
      & (cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_tmp==5'b11111))
      | (cfg_proc_precision_rsci_d!=2'b10))) | cfg_mode_eql_rsci_d;
  assign or_13_nl = (~(cvt_1_FpMantRNE_24U_11U_else_and_svs | (cfg_proc_precision_rsci_d!=2'b10)))
      | cfg_mode_eql_rsci_d;
  assign nor_2080_nl = ~(cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1
      | (~ cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_itm_8_1));
  assign mux_1_nl = MUX_s_1_2_2((or_13_nl), (or_11_nl), nor_2080_nl);
  assign mux_2_nl = MUX_s_1_2_2((mux_1_nl), (or_9_nl), IsNaN_8U_23U_IsNaN_8U_23U_nor_tmp);
  assign and_98_nl = chn_in_rsci_bawt & (mux_2_nl);
  assign and_2240_nl = ((~(((~(cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_2
      & (~ FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_2)
      & cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_2
      & FpWidthDec_8U_23U_5U_10U_1U_1U_nand_itm_2)) & cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_2)
      | (cfg_proc_precision_1_sva_st_64!=2'b10))) | cfg_mode_eql_1_sva_4) & main_stage_v_1;
  assign or_14_nl = (~ cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_st_2;
  assign mux_3_nl = MUX_s_1_2_2((and_2240_nl), and_2239_cse, or_14_nl);
  assign and_2242_nl = (nor_8_cse | cfg_mode_eql_1_sva_4) & main_stage_v_1;
  assign nor_2_nl = ~(IsNaN_8U_23U_land_1_lpi_1_dfm_3 | (~ cvt_1_FpMantRNE_24U_11U_else_and_svs_2));
  assign mux_4_nl = MUX_s_1_2_2((and_2242_nl), (mux_3_nl), nor_2_nl);
  assign mux_5_nl = MUX_s_1_2_2((mux_4_nl), (and_98_nl), or_5189_cse);
  assign or_19_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_st_2
      | (~ cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_2)
      | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~ main_stage_v_1)
      | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign nor_10_nl = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_st_2
      | (~ cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_2));
  assign mux_7_nl = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, nor_10_nl);
  assign or_17_nl = (~ cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_itm_8_1) | cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1;
  assign mux_8_nl = MUX_s_1_2_2((mux_7_nl), (or_19_nl), or_17_nl);
  assign mux_9_nl = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_2);
  assign or_28_nl = (~ cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_svs_st_2)
      | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~ main_stage_v_1)
      | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_10_nl = MUX_s_1_2_2((or_28_nl), (mux_9_nl), cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_itm_8_1);
  assign nor_2075_nl = ~(cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1
      | cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1 | (~ cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt));
  assign nor_2076_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | (~ cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_st_2
      | cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2);
  assign mux_11_nl = MUX_s_1_2_2((nor_2076_nl), (nor_2075_nl), or_5189_cse);
  assign nor_12_nl = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_st_2
      | (~ cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2));
  assign mux_13_nl = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, nor_12_nl);
  assign or_35_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_st_2
      | (~ cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2)
      | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~ main_stage_v_1)
      | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign nor_11_nl = ~(cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1
      | (~ cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1));
  assign mux_14_nl = MUX_s_1_2_2((or_35_nl), (mux_13_nl), nor_11_nl);
  assign mux_15_nl = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2);
  assign or_37_nl = (~ cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2)
      | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~ main_stage_v_1)
      | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_16_nl = MUX_s_1_2_2((or_37_nl), (mux_15_nl), cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1);
  assign nor_2073_nl = ~(cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1
      | cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1 | (~ cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt));
  assign nor_2074_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | (~ cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_st_2
      | cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2);
  assign mux_17_nl = MUX_s_1_2_2((nor_2074_nl), (nor_2073_nl), or_5189_cse);
  assign nor_14_nl = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_st_2
      | (~ cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2));
  assign mux_18_nl = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, nor_14_nl);
  assign or_43_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_st_2
      | (~ cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2)
      | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~ main_stage_v_1)
      | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign nor_13_nl = ~(cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1
      | (~ cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1));
  assign mux_19_nl = MUX_s_1_2_2((or_43_nl), (mux_18_nl), nor_13_nl);
  assign mux_20_nl = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2);
  assign or_45_nl = (~ cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2)
      | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~ main_stage_v_1)
      | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_21_nl = MUX_s_1_2_2((or_45_nl), (mux_20_nl), cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1);
  assign nor_2071_nl = ~(cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1
      | cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt));
  assign nor_2072_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | (~ cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_st_2
      | cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2);
  assign mux_22_nl = MUX_s_1_2_2((nor_2072_nl), (nor_2071_nl), or_5189_cse);
  assign nor_16_nl = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_st_2
      | (~ cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2));
  assign mux_23_nl = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, nor_16_nl);
  assign or_51_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_st_2
      | (~ cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2)
      | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~ main_stage_v_1)
      | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign nor_15_nl = ~(cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1
      | (~ cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1));
  assign mux_24_nl = MUX_s_1_2_2((or_51_nl), (mux_23_nl), nor_15_nl);
  assign mux_25_nl = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2);
  assign or_53_nl = (~ cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2)
      | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~ main_stage_v_1)
      | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_26_nl = MUX_s_1_2_2((or_53_nl), (mux_25_nl), cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1);
  assign or_56_nl = cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_st_2
      | (~ cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2)
      | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_27_nl = MUX_s_1_2_2((or_56_nl), or_tmp_19, or_5189_cse);
  assign or_58_nl = (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_st_2
      | (~ cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2)
      | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign nor_17_nl = ~(cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1
      | cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1 | (~ cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1));
  assign mux_28_nl = MUX_s_1_2_2((or_58_nl), (mux_27_nl), nor_17_nl);
  assign or_61_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_st_2
      | (~ cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2)
      | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_29_nl = MUX_s_1_2_2((or_61_nl), or_tmp_19, or_5189_cse);
  assign or_63_nl = (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_st_2
      | (~ cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2)
      | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign nor_18_nl = ~(cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1
      | (~ cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1));
  assign mux_30_nl = MUX_s_1_2_2((or_63_nl), (mux_29_nl), nor_18_nl);
  assign nand_235_nl = ~(cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2
      & main_stage_v_1 & (cfg_proc_precision_1_sva_st_64==2'b10));
  assign mux_31_nl = MUX_s_1_2_2((nand_235_nl), or_tmp_19, or_5189_cse);
  assign or_68_nl = (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~
      cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2)
      | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_32_nl = MUX_s_1_2_2((or_68_nl), (mux_31_nl), cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1);
  assign or_71_nl = cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_st_2
      | (~ cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2)
      | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_33_nl = MUX_s_1_2_2((or_71_nl), or_tmp_19, or_5189_cse);
  assign or_73_nl = (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_st_2
      | (~ cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2)
      | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign nor_19_nl = ~(cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1
      | cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1));
  assign mux_34_nl = MUX_s_1_2_2((or_73_nl), (mux_33_nl), nor_19_nl);
  assign or_76_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_st_2
      | (~ cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2)
      | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_35_nl = MUX_s_1_2_2((or_76_nl), or_tmp_19, or_5189_cse);
  assign or_78_nl = (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_st_2
      | (~ cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2)
      | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign nor_20_nl = ~(cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1
      | (~ cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1));
  assign mux_36_nl = MUX_s_1_2_2((or_78_nl), (mux_35_nl), nor_20_nl);
  assign nand_234_nl = ~(cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
      & main_stage_v_1 & (cfg_proc_precision_1_sva_st_64==2'b10));
  assign mux_37_nl = MUX_s_1_2_2((nand_234_nl), or_tmp_19, or_5189_cse);
  assign or_83_nl = (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~
      cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2)
      | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_38_nl = MUX_s_1_2_2((or_83_nl), (mux_37_nl), cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1);
  assign mux_40_nl = MUX_s_1_2_2(mux_tmp_39, or_tmp_24, cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2);
  assign or_88_nl = cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2
      | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~ cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_st_2
      | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign nor_21_nl = ~(cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1
      | cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1));
  assign mux_41_nl = MUX_s_1_2_2((or_88_nl), (mux_40_nl), nor_21_nl);
  assign or_90_nl = (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~
      cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_st_2
      | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign nor_22_nl = ~(cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1
      | (~ cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1));
  assign mux_42_nl = MUX_s_1_2_2((or_90_nl), mux_tmp_39, nor_22_nl);
  assign nand_233_nl = ~(cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
      & main_stage_v_1 & (cfg_proc_precision_1_sva_st_64==2'b10));
  assign mux_43_nl = MUX_s_1_2_2((nand_233_nl), or_tmp_19, or_5189_cse);
  assign or_95_nl = (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~
      cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2)
      | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_44_nl = MUX_s_1_2_2((or_95_nl), (mux_43_nl), cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1);
  assign nor_2069_nl = ~(cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1
      | cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 | (~ cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt));
  assign nor_2070_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | (~ cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_st_2
      | cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2);
  assign mux_45_nl = MUX_s_1_2_2((nor_2070_nl), (nor_2069_nl), or_5189_cse);
  assign nor_24_nl = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_st_2
      | (~ cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2));
  assign mux_46_nl = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, nor_24_nl);
  assign or_101_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_st_2
      | (~ cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2)
      | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~ main_stage_v_1)
      | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign nor_23_nl = ~(cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1
      | (~ cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1));
  assign mux_47_nl = MUX_s_1_2_2((or_101_nl), (mux_46_nl), nor_23_nl);
  assign mux_48_nl = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2);
  assign or_103_nl = (~ cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2)
      | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~ main_stage_v_1)
      | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_49_nl = MUX_s_1_2_2((or_103_nl), (mux_48_nl), cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1);
  assign nor_2067_nl = ~(cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1
      | cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1 | (~ cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt));
  assign nor_2068_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | (~ cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_st_2
      | cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2);
  assign mux_50_nl = MUX_s_1_2_2((nor_2068_nl), (nor_2067_nl), or_5189_cse);
  assign nor_26_nl = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_st_2
      | (~ cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2));
  assign mux_51_nl = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, nor_26_nl);
  assign or_109_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_st_2
      | (~ cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2)
      | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~ main_stage_v_1)
      | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign nor_25_nl = ~(cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1
      | (~ cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1));
  assign mux_52_nl = MUX_s_1_2_2((or_109_nl), (mux_51_nl), nor_25_nl);
  assign mux_53_nl = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2);
  assign or_111_nl = (~ cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_1_svs_st_2)
      | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~ main_stage_v_1)
      | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_54_nl = MUX_s_1_2_2((or_111_nl), (mux_53_nl), cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1);
  assign or_114_nl = cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_st_2
      | (~ cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2)
      | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_55_nl = MUX_s_1_2_2((or_114_nl), or_tmp_19, or_5189_cse);
  assign or_116_nl = (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt |
      cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_st_2
      | (~ cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2)
      | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign nor_27_nl = ~(cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1
      | cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1));
  assign mux_56_nl = MUX_s_1_2_2((or_116_nl), (mux_55_nl), nor_27_nl);
  assign or_119_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_st_2
      | (~ cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2)
      | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_57_nl = MUX_s_1_2_2((or_119_nl), or_tmp_19, or_5189_cse);
  assign or_121_nl = (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt |
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_st_2
      | (~ cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2)
      | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign nor_28_nl = ~(cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1
      | (~ cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1));
  assign mux_58_nl = MUX_s_1_2_2((or_121_nl), (mux_57_nl), nor_28_nl);
  assign nand_232_nl = ~(cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
      & main_stage_v_1 & (cfg_proc_precision_1_sva_st_64==2'b10));
  assign mux_59_nl = MUX_s_1_2_2((nand_232_nl), or_tmp_19, or_5189_cse);
  assign or_126_nl = (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt |
      (~ cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2)
      | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_60_nl = MUX_s_1_2_2((or_126_nl), (mux_59_nl), cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1);
  assign nor_2065_nl = ~(cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1
      | cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt));
  assign nor_2066_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | (~ cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_st_2
      | cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2);
  assign mux_61_nl = MUX_s_1_2_2((nor_2066_nl), (nor_2065_nl), or_5189_cse);
  assign nor_30_nl = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_st_2
      | (~ cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2));
  assign mux_62_nl = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, nor_30_nl);
  assign or_132_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_st_2
      | (~ cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2)
      | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~ main_stage_v_1)
      | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign nor_29_nl = ~(cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1
      | (~ cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1));
  assign mux_63_nl = MUX_s_1_2_2((or_132_nl), (mux_62_nl), nor_29_nl);
  assign mux_64_nl = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2);
  assign or_134_nl = (~ cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2)
      | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~ main_stage_v_1)
      | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_65_nl = MUX_s_1_2_2((or_134_nl), (mux_64_nl), cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1);
  assign nor_2063_nl = ~(cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1
      | cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 | (~ cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt));
  assign nor_2064_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | (~ cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_st_2
      | cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2);
  assign mux_66_nl = MUX_s_1_2_2((nor_2064_nl), (nor_2063_nl), or_5189_cse);
  assign nor_32_nl = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_st_2
      | (~ cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2));
  assign mux_67_nl = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, nor_32_nl);
  assign or_140_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_st_2
      | (~ cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2)
      | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~ main_stage_v_1)
      | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign nor_31_nl = ~(cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1
      | (~ cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1));
  assign mux_68_nl = MUX_s_1_2_2((or_140_nl), (mux_67_nl), nor_31_nl);
  assign mux_69_nl = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2);
  assign or_142_nl = (~ cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2)
      | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~ main_stage_v_1)
      | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_70_nl = MUX_s_1_2_2((or_142_nl), (mux_69_nl), cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1);
  assign or_145_nl = cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_st_2
      | (~ cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2)
      | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_71_nl = MUX_s_1_2_2((or_145_nl), or_tmp_19, or_5189_cse);
  assign or_147_nl = (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt |
      cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_st_2
      | (~ cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2)
      | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign nor_33_nl = ~(cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1
      | cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1));
  assign mux_72_nl = MUX_s_1_2_2((or_147_nl), (mux_71_nl), nor_33_nl);
  assign or_150_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_st_2
      | (~ cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2)
      | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_73_nl = MUX_s_1_2_2((or_150_nl), or_tmp_19, or_5189_cse);
  assign or_152_nl = (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt |
      FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_st_2
      | (~ cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2)
      | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign nor_34_nl = ~(cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1
      | (~ cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1));
  assign mux_74_nl = MUX_s_1_2_2((or_152_nl), (mux_73_nl), nor_34_nl);
  assign nand_231_nl = ~(cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2
      & main_stage_v_1 & (cfg_proc_precision_1_sva_st_64==2'b10));
  assign mux_75_nl = MUX_s_1_2_2((nand_231_nl), or_tmp_19, or_5189_cse);
  assign or_157_nl = (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt |
      (~ cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_2_svs_st_2)
      | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_76_nl = MUX_s_1_2_2((or_157_nl), (mux_75_nl), cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1);
  assign nor_2061_nl = ~(cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1
      | cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 | (~ cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt));
  assign nor_2062_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | (~ cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_st_2
      | cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2);
  assign mux_77_nl = MUX_s_1_2_2((nor_2062_nl), (nor_2061_nl), or_5189_cse);
  assign nor_36_nl = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_st_2
      | (~ cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2));
  assign mux_78_nl = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, nor_36_nl);
  assign or_163_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_st_2
      | (~ cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2)
      | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~ main_stage_v_1)
      | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign nor_35_nl = ~(cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1
      | (~ cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1));
  assign mux_79_nl = MUX_s_1_2_2((or_163_nl), (mux_78_nl), nor_35_nl);
  assign mux_80_nl = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2);
  assign or_165_nl = (~ cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2)
      | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~ main_stage_v_1)
      | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_81_nl = MUX_s_1_2_2((or_165_nl), (mux_80_nl), cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1);
  assign nor_2059_nl = ~(cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1
      | cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 | (~ cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt));
  assign nor_2060_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | (~ cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_st_2
      | cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2);
  assign mux_82_nl = MUX_s_1_2_2((nor_2060_nl), (nor_2059_nl), or_5189_cse);
  assign nor_38_nl = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_st_2
      | (~ cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2));
  assign mux_83_nl = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, nor_38_nl);
  assign or_171_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_st_2
      | (~ cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2)
      | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~ main_stage_v_1)
      | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign nor_37_nl = ~(cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1
      | (~ cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1));
  assign mux_84_nl = MUX_s_1_2_2((or_171_nl), (mux_83_nl), nor_37_nl);
  assign mux_85_nl = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2);
  assign or_173_nl = (~ cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_3_svs_st_2)
      | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~ main_stage_v_1)
      | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_86_nl = MUX_s_1_2_2((or_173_nl), (mux_85_nl), cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1);
  assign nor_2057_nl = ~(cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_itm_8_1
      | cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_itm_7_1 | (~ cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt));
  assign nor_2058_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | (~ cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_4_svs_st_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_2
      | cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_st_2);
  assign mux_87_nl = MUX_s_1_2_2((nor_2058_nl), (nor_2057_nl), or_5189_cse);
  assign nor_40_nl = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_2
      | (~ cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_4_svs_st_2));
  assign mux_88_nl = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, nor_40_nl);
  assign or_179_nl = FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_2
      | (~ cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_4_svs_st_2)
      | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~ main_stage_v_1)
      | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign nor_39_nl = ~(cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_itm_7_1
      | (~ cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_itm_8_1));
  assign mux_89_nl = MUX_s_1_2_2((or_179_nl), (mux_88_nl), nor_39_nl);
  assign mux_90_nl = MUX_s_1_2_2(or_tmp_24, mux_tmp_6, cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_4_svs_st_2);
  assign or_181_nl = (~ cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_8_4_svs_st_2)
      | (~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt | (~ main_stage_v_1)
      | (cfg_proc_precision_1_sva_st_64!=2'b10);
  assign mux_91_nl = MUX_s_1_2_2((or_181_nl), (mux_90_nl), cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_itm_8_1);
  assign FpMantRNE_24U_11U_else_mux_31_nl = MUX_s_1_2_2(cvt_16_FpMantRNE_24U_11U_else_and_4_tmp,
      cvt_16_FpMantRNE_24U_11U_else_and_4_svs, or_dcpl_320);
  assign FpMantRNE_24U_11U_else_mux_29_nl = MUX_s_1_2_2(cvt_15_FpMantRNE_24U_11U_else_and_3_tmp,
      cvt_15_FpMantRNE_24U_11U_else_and_3_svs, or_dcpl_322);
  assign FpMantRNE_24U_11U_else_mux_27_nl = MUX_s_1_2_2(cvt_14_FpMantRNE_24U_11U_else_and_3_tmp,
      cvt_14_FpMantRNE_24U_11U_else_and_3_svs, or_dcpl_324);
  assign FpMantRNE_24U_11U_else_mux_25_nl = MUX_s_1_2_2(cvt_13_FpMantRNE_24U_11U_else_and_2_tmp,
      cvt_13_FpMantRNE_24U_11U_else_and_2_svs, or_dcpl_326);
  assign FpMantRNE_24U_11U_else_mux_23_nl = MUX_s_1_2_2(cvt_12_FpMantRNE_24U_11U_else_and_3_tmp,
      cvt_12_FpMantRNE_24U_11U_else_and_3_svs, or_dcpl_328);
  assign FpMantRNE_24U_11U_else_mux_21_nl = MUX_s_1_2_2(cvt_11_FpMantRNE_24U_11U_else_and_2_tmp,
      cvt_11_FpMantRNE_24U_11U_else_and_2_svs, or_dcpl_330);
  assign FpMantRNE_24U_11U_else_mux_19_nl = MUX_s_1_2_2(cvt_10_FpMantRNE_24U_11U_else_and_2_tmp,
      cvt_10_FpMantRNE_24U_11U_else_and_2_svs, or_dcpl_332);
  assign FpMantRNE_24U_11U_else_mux_17_nl = MUX_s_1_2_2(cvt_9_FpMantRNE_24U_11U_else_and_1_tmp,
      cvt_9_FpMantRNE_24U_11U_else_and_1_svs, or_dcpl_334);
  assign FpMantRNE_24U_11U_else_mux_15_nl = MUX_s_1_2_2(cvt_8_FpMantRNE_24U_11U_else_and_3_tmp,
      cvt_8_FpMantRNE_24U_11U_else_and_3_svs, or_dcpl_336);
  assign FpMantRNE_24U_11U_else_mux_13_nl = MUX_s_1_2_2(cvt_7_FpMantRNE_24U_11U_else_and_2_tmp,
      cvt_7_FpMantRNE_24U_11U_else_and_2_svs, or_dcpl_338);
  assign FpMantRNE_24U_11U_else_mux_11_nl = MUX_s_1_2_2(cvt_6_FpMantRNE_24U_11U_else_and_2_tmp,
      cvt_6_FpMantRNE_24U_11U_else_and_2_svs, or_dcpl_340);
  assign FpMantRNE_24U_11U_else_mux_9_nl = MUX_s_1_2_2(cvt_5_FpMantRNE_24U_11U_else_and_1_tmp,
      cvt_5_FpMantRNE_24U_11U_else_and_1_svs, or_dcpl_342);
  assign FpMantRNE_24U_11U_else_mux_7_nl = MUX_s_1_2_2(cvt_4_FpMantRNE_24U_11U_else_and_2_tmp,
      cvt_4_FpMantRNE_24U_11U_else_and_2_svs, or_dcpl_344);
  assign FpMantRNE_24U_11U_else_mux_5_nl = MUX_s_1_2_2(cvt_3_FpMantRNE_24U_11U_else_and_1_tmp,
      cvt_3_FpMantRNE_24U_11U_else_and_1_svs, or_dcpl_346);
  assign FpMantRNE_24U_11U_else_mux_3_nl = MUX_s_1_2_2(cvt_2_FpMantRNE_24U_11U_else_and_1_tmp,
      cvt_2_FpMantRNE_24U_11U_else_and_1_svs, or_dcpl_348);
  assign FpMantRNE_24U_11U_else_mux_1_nl = MUX_s_1_2_2(cvt_1_FpMantRNE_24U_11U_else_and_tmp,
      cvt_1_FpMantRNE_24U_11U_else_and_svs, or_dcpl_350);
  assign nl_cvt_2_IntSubExt_32U_32U_33U_o_acc_1_nl = conv_s2s_32_33(chn_in_rsci_d_mxwt[63:32])
      - conv_s2s_32_33(cfg_offset_rsci_d);
  assign cvt_2_IntSubExt_32U_32U_33U_o_acc_1_nl = nl_cvt_2_IntSubExt_32U_32U_33U_o_acc_1_nl[32:0];
  assign nl_cvt_3_IntSubExt_32U_32U_33U_o_acc_1_nl = conv_s2s_32_33(chn_in_rsci_d_mxwt[95:64])
      - conv_s2s_32_33(cfg_offset_rsci_d);
  assign cvt_3_IntSubExt_32U_32U_33U_o_acc_1_nl = nl_cvt_3_IntSubExt_32U_32U_33U_o_acc_1_nl[32:0];
  assign nl_cvt_9_IntSubExt_32U_32U_33U_o_acc_1_nl = conv_s2s_32_33(chn_in_rsci_d_mxwt[287:256])
      - conv_s2s_32_33(cfg_offset_rsci_d);
  assign cvt_9_IntSubExt_32U_32U_33U_o_acc_1_nl = nl_cvt_9_IntSubExt_32U_32U_33U_o_acc_1_nl[32:0];
  assign nl_cvt_4_IntSubExt_32U_32U_33U_o_acc_2_nl = conv_s2s_32_33(chn_in_rsci_d_mxwt[127:96])
      - conv_s2s_32_33(cfg_offset_rsci_d);
  assign cvt_4_IntSubExt_32U_32U_33U_o_acc_2_nl = nl_cvt_4_IntSubExt_32U_32U_33U_o_acc_2_nl[32:0];
  assign cvt_4_IntMulExt_33U_16U_49U_o_mul_2_nl = conv_s2u_49_49($signed((cvt_4_IntSubExt_32U_32U_33U_o_acc_2_nl))
      * $signed((cfg_scale_rsci_d)));
  assign nl_cvt_6_IntSubExt_32U_32U_33U_o_acc_2_nl = conv_s2s_32_33(chn_in_rsci_d_mxwt[191:160])
      - conv_s2s_32_33(cfg_offset_rsci_d);
  assign cvt_6_IntSubExt_32U_32U_33U_o_acc_2_nl = nl_cvt_6_IntSubExt_32U_32U_33U_o_acc_2_nl[32:0];
  assign cvt_6_IntMulExt_33U_16U_49U_o_mul_2_nl = conv_s2u_49_49($signed((cvt_6_IntSubExt_32U_32U_33U_o_acc_2_nl))
      * $signed((cfg_scale_rsci_d)));
  assign nl_cvt_8_IntSubExt_32U_32U_33U_o_acc_3_nl = conv_s2s_32_33(chn_in_rsci_d_mxwt[255:224])
      - conv_s2s_32_33(cfg_offset_rsci_d);
  assign cvt_8_IntSubExt_32U_32U_33U_o_acc_3_nl = nl_cvt_8_IntSubExt_32U_32U_33U_o_acc_3_nl[32:0];
  assign cvt_8_IntMulExt_33U_16U_49U_o_mul_3_nl = conv_s2u_49_49($signed((cvt_8_IntSubExt_32U_32U_33U_o_acc_3_nl))
      * $signed((cfg_scale_rsci_d)));
  assign nl_cvt_7_IntSubExt_32U_32U_33U_o_acc_2_nl = conv_s2s_32_33(chn_in_rsci_d_mxwt[223:192])
      - conv_s2s_32_33(cfg_offset_rsci_d);
  assign cvt_7_IntSubExt_32U_32U_33U_o_acc_2_nl = nl_cvt_7_IntSubExt_32U_32U_33U_o_acc_2_nl[32:0];
  assign cvt_7_IntMulExt_33U_16U_49U_o_mul_2_nl = conv_s2u_49_49($signed((cvt_7_IntSubExt_32U_32U_33U_o_acc_2_nl))
      * $signed((cfg_scale_rsci_d)));
  assign nl_cvt_10_IntSubExt_32U_32U_33U_o_acc_2_nl = conv_s2s_32_33(chn_in_rsci_d_mxwt[319:288])
      - conv_s2s_32_33(cfg_offset_rsci_d);
  assign cvt_10_IntSubExt_32U_32U_33U_o_acc_2_nl = nl_cvt_10_IntSubExt_32U_32U_33U_o_acc_2_nl[32:0];
  assign cvt_10_IntMulExt_33U_16U_49U_o_mul_2_nl = conv_s2u_49_49($signed((cvt_10_IntSubExt_32U_32U_33U_o_acc_2_nl))
      * $signed((cfg_scale_rsci_d)));
  assign nl_cvt_12_IntSubExt_32U_32U_33U_o_acc_3_nl = conv_s2s_32_33(chn_in_rsci_d_mxwt[383:352])
      - conv_s2s_32_33(cfg_offset_rsci_d);
  assign cvt_12_IntSubExt_32U_32U_33U_o_acc_3_nl = nl_cvt_12_IntSubExt_32U_32U_33U_o_acc_3_nl[32:0];
  assign cvt_12_IntMulExt_33U_16U_49U_o_mul_3_nl = conv_s2u_49_49($signed((cvt_12_IntSubExt_32U_32U_33U_o_acc_3_nl))
      * $signed((cfg_scale_rsci_d)));
  assign nl_cvt_11_IntSubExt_32U_32U_33U_o_acc_2_nl = conv_s2s_32_33(chn_in_rsci_d_mxwt[351:320])
      - conv_s2s_32_33(cfg_offset_rsci_d);
  assign cvt_11_IntSubExt_32U_32U_33U_o_acc_2_nl = nl_cvt_11_IntSubExt_32U_32U_33U_o_acc_2_nl[32:0];
  assign cvt_11_IntMulExt_33U_16U_49U_o_mul_2_nl = conv_s2u_49_49($signed((cvt_11_IntSubExt_32U_32U_33U_o_acc_2_nl))
      * $signed((cfg_scale_rsci_d)));
  assign nl_cvt_14_IntSubExt_32U_32U_33U_o_acc_3_nl = conv_s2s_32_33(chn_in_rsci_d_mxwt[447:416])
      - conv_s2s_32_33(cfg_offset_rsci_d);
  assign cvt_14_IntSubExt_32U_32U_33U_o_acc_3_nl = nl_cvt_14_IntSubExt_32U_32U_33U_o_acc_3_nl[32:0];
  assign cvt_14_IntMulExt_33U_16U_49U_o_mul_3_nl = conv_s2u_49_49($signed((cvt_14_IntSubExt_32U_32U_33U_o_acc_3_nl))
      * $signed((cfg_scale_rsci_d)));
  assign nl_cvt_16_IntSubExt_32U_32U_33U_o_acc_4_nl = conv_s2s_32_33(chn_in_rsci_d_mxwt[511:480])
      - conv_s2s_32_33(cfg_offset_rsci_d);
  assign cvt_16_IntSubExt_32U_32U_33U_o_acc_4_nl = nl_cvt_16_IntSubExt_32U_32U_33U_o_acc_4_nl[32:0];
  assign cvt_16_IntMulExt_33U_16U_49U_o_mul_4_nl = conv_s2u_49_49($signed((cvt_16_IntSubExt_32U_32U_33U_o_acc_4_nl))
      * $signed((cfg_scale_rsci_d)));
  assign nl_cvt_15_IntSubExt_32U_32U_33U_o_acc_3_nl = conv_s2s_32_33(chn_in_rsci_d_mxwt[479:448])
      - conv_s2s_32_33(cfg_offset_rsci_d);
  assign cvt_15_IntSubExt_32U_32U_33U_o_acc_3_nl = nl_cvt_15_IntSubExt_32U_32U_33U_o_acc_3_nl[32:0];
  assign cvt_15_IntMulExt_33U_16U_49U_o_mul_3_nl = conv_s2u_49_49($signed((cvt_15_IntSubExt_32U_32U_33U_o_acc_3_nl))
      * $signed((cfg_scale_rsci_d)));
  assign nl_cvt_13_IntSubExt_32U_32U_33U_o_acc_2_nl = conv_s2s_32_33(chn_in_rsci_d_mxwt[415:384])
      - conv_s2s_32_33(cfg_offset_rsci_d);
  assign cvt_13_IntSubExt_32U_32U_33U_o_acc_2_nl = nl_cvt_13_IntSubExt_32U_32U_33U_o_acc_2_nl[32:0];
  assign cvt_13_IntMulExt_33U_16U_49U_o_mul_2_nl = conv_s2u_49_49($signed((cvt_13_IntSubExt_32U_32U_33U_o_acc_2_nl))
      * $signed((cfg_scale_rsci_d)));
  assign nl_cvt_5_IntSubExt_32U_32U_33U_o_acc_1_nl = conv_s2s_32_33(chn_in_rsci_d_mxwt[159:128])
      - conv_s2s_32_33(cfg_offset_rsci_d);
  assign cvt_5_IntSubExt_32U_32U_33U_o_acc_1_nl = nl_cvt_5_IntSubExt_32U_32U_33U_o_acc_1_nl[32:0];
  assign mux_154_nl = MUX_s_1_2_2(mux_110_cse, (~ or_4550_cse), reg_cfg_proc_precision_1_sva_st_40_cse[1]);
  assign mux_155_nl = MUX_s_1_2_2((mux_154_nl), mux_110_cse, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign and_132_nl = main_stage_v_1 & (mux_155_nl);
  assign mux_159_nl = MUX_s_1_2_2((and_132_nl), chn_in_rsci_bawt, or_5189_cse);
  assign nl_cvt_1_IntSubExt_32U_32U_33U_o_acc_nl = conv_s2s_32_33(chn_in_rsci_d_mxwt[31:0])
      - conv_s2s_32_33(cfg_offset_rsci_d);
  assign cvt_1_IntSubExt_32U_32U_33U_o_acc_nl = nl_cvt_1_IntSubExt_32U_32U_33U_o_acc_nl[32:0];
  assign nl_cvt_1_FpFloatToInt_16U_5U_10U_shift_acc_itm_2 = conv_u2u_4_5({(~ FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_7_4_mx0w0)
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_7_3_0_mx0w0[3:1]))})
      + 5'b11101;
  assign nor_2048_nl = ~((~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149[1])
      | (cfg_proc_precision_1_sva_st_65[0]) | nand_219_cse);
  assign mux_162_nl = MUX_s_1_2_2((nor_2048_nl), nor_2047_cse, or_5189_cse);
  assign nl_cvt_2_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2 = conv_u2u_4_5({(~ FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_7_4_mx0w0)
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_7_3_0_mx0w0[3:1]))})
      + 5'b11101;
  assign nl_cvt_3_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2 = conv_u2u_4_5({(~ FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_7_4_mx0w0)
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_3_lpi_1_dfm_7_3_0_mx0w0[3:1]))})
      + 5'b11101;
  assign nl_cvt_4_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 = conv_u2u_4_5({(~ FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_7_4_mx0w0)
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_4_lpi_1_dfm_7_3_0_mx0w0[3:1]))})
      + 5'b11101;
  assign nl_cvt_5_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2 = conv_u2u_4_5({(~ FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_7_4_mx0w0)
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_5_lpi_1_dfm_7_3_0_mx0w0[3:1]))})
      + 5'b11101;
  assign mux_167_nl = MUX_s_1_2_2(mux_166_cse, or_303_cse, or_300_cse);
  assign nl_cvt_6_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 = conv_u2u_4_5({(~ FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_7_4_mx0w0)
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_6_lpi_1_dfm_7_3_0_mx0w0[3:1]))})
      + 5'b11101;
  assign nl_cvt_7_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 = conv_u2u_4_5({(~ FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_7_4_mx0w0)
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_7_lpi_1_dfm_7_3_0_mx0w0[3:1]))})
      + 5'b11101;
  assign nl_cvt_8_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2 = conv_u2u_4_5({(~ FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_7_4_mx0w0)
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_8_lpi_1_dfm_7_3_0_mx0w0[3:1]))})
      + 5'b11101;
  assign nl_cvt_10_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 = conv_u2u_4_5({(~
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_7_4_mx0w0) , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_10_lpi_1_dfm_7_3_0_mx0w0[3:1]))})
      + 5'b11101;
  assign nl_cvt_11_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 = conv_u2u_4_5({(~
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_7_4_mx0w0) , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_11_lpi_1_dfm_7_3_0_mx0w0[3:1]))})
      + 5'b11101;
  assign nl_cvt_13_FpFloatToInt_16U_5U_10U_shift_acc_2_itm_2 = conv_u2u_4_5({(~
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_7_4_mx0w0) , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_13_lpi_1_dfm_7_3_0_mx0w0[3:1]))})
      + 5'b11101;
  assign nl_cvt_15_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2 = conv_u2u_4_5({(~
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_7_4_mx0w0) , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_7_3_0_mx0w0[3:1]))})
      + 5'b11101;
  assign nl_cvt_9_FpFloatToInt_16U_5U_10U_shift_acc_1_itm_2 = conv_u2u_4_5({(~ FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_7_4_mx0w0)
      , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_9_lpi_1_dfm_7_3_0_mx0w0[3:1]))})
      + 5'b11101;
  assign nl_cvt_12_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2 = conv_u2u_4_5({(~
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_7_4_mx0w0) , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_12_lpi_1_dfm_7_3_0_mx0w0[3:1]))})
      + 5'b11101;
  assign nl_cvt_14_FpFloatToInt_16U_5U_10U_shift_acc_3_itm_2 = conv_u2u_4_5({(~
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_7_4_mx0w0) , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_14_lpi_1_dfm_7_3_0_mx0w0[3:1]))})
      + 5'b11101;
  assign mux_190_nl = MUX_s_1_2_2((~ main_stage_v_2), or_tmp_378, cfg_mode_eql_1_sva_5);
  assign mux_191_nl = MUX_s_1_2_2((mux_190_nl), mux_tmp_189, or_5189_cse);
  assign nl_cvt_16_FpFloatToInt_16U_5U_10U_shift_acc_4_itm_2 = conv_u2u_4_5({(~
      FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_7_4_mx0w0) , (~ (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_lpi_1_dfm_7_3_0_mx0w0[3:1]))})
      + 5'b11101;
  assign mux_192_nl = MUX_s_1_2_2(or_tmp_378, or_306_cse, or_5189_cse);
  assign and_143_nl = main_stage_v_1 & cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_tmp
      & or_4550_cse;
  assign mux_232_nl = MUX_s_1_2_2(and_2237_cse, (and_143_nl), or_5189_cse);
  assign and_145_nl = or_5189_cse & main_stage_v_1 & cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_tmp
      & or_4550_cse;
  assign mux_235_nl = MUX_s_1_2_2((and_145_nl), (mux_232_nl), cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_svs_2);
  assign nor_2020_nl = ~((cfg_out_precision_1_sva_st_154!=2'b00) | (~ mux_tmp_236));
  assign mux_237_nl = MUX_s_1_2_2((nor_2020_nl), mux_tmp_236, cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_tmp);
  assign mux_238_nl = MUX_s_1_2_2(main_stage_v_1, (mux_237_nl), or_419_cse);
  assign and_2857_nl = mux_tmp_239 & (~ or_425_cse);
  assign mux_241_nl = MUX_s_1_2_2((and_2857_nl), mux_tmp_239, cvt_1_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_svs_2);
  assign mux_242_nl = MUX_s_1_2_2(main_stage_v_2, (mux_241_nl), or_423_cse);
  assign mux_243_nl = MUX_s_1_2_2((mux_242_nl), (mux_238_nl), or_5189_cse);
  assign nor_2016_nl = ~((cfg_out_precision_1_sva_st_154!=2'b10) | (~ and_tmp_11));
  assign mux_246_nl = MUX_s_1_2_2(and_2237_cse, (nor_2016_nl), or_5189_cse);
  assign nor_2017_nl = ~(nor_2040_cse | (cfg_out_precision_1_sva_st_154!=2'b10) |
      (~ and_tmp_11));
  assign mux_247_nl = MUX_s_1_2_2((nor_2017_nl), (mux_246_nl), nor_57_cse);
  assign and_147_nl = main_stage_v_1 & cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp
      & and_tmp_12;
  assign mux_248_nl = MUX_s_1_2_2(and_tmp_52, (and_147_nl), or_5189_cse);
  assign mux_254_nl = MUX_s_1_2_2(main_stage_v_2, and_1078_cse, or_451_cse);
  assign mux_255_nl = MUX_s_1_2_2((mux_254_nl), mux_tmp_251, or_5189_cse);
  assign and_2234_nl = (cfg_out_precision_1_sva_st_149[1]) & cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign mux_256_nl = MUX_s_1_2_2((mux_255_nl), mux_tmp_253, and_2234_nl);
  assign mux_257_nl = MUX_s_1_2_2((mux_256_nl), mux_tmp_253, cfg_out_precision_1_sva_st_149[0]);
  assign mux_260_nl = MUX_s_1_2_2(nor_2011_cse, mux_tmp_259, cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp);
  assign mux_261_nl = MUX_s_1_2_2(main_stage_v_1, (mux_260_nl), or_419_cse);
  assign and_2233_nl = IntShiftRightSat_49U_6U_17U_lor_3_lpi_1_dfm & mux_tmp_263;
  assign mux_264_nl = MUX_s_1_2_2(mux_tmp_263, (and_2233_nl), or_461_cse);
  assign mux_265_nl = MUX_s_1_2_2((mux_264_nl), mux_tmp_263, cvt_2_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2);
  assign mux_266_nl = MUX_s_1_2_2(main_stage_v_2, (mux_265_nl), or_423_cse);
  assign mux_267_nl = MUX_s_1_2_2((mux_266_nl), (mux_261_nl), or_5189_cse);
  assign mux_270_nl = MUX_s_1_2_2(and_1078_cse, nor_2004_cse, or_5189_cse);
  assign mux_271_nl = MUX_s_1_2_2(nor_2005_cse, (mux_270_nl), nor_63_cse);
  assign and_156_nl = main_stage_v_1 & cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp
      & and_tmp_12;
  assign and_160_nl = main_stage_v_2 & cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2
      & and_tmp_50;
  assign mux_275_nl = MUX_s_1_2_2((and_160_nl), (and_156_nl), or_5189_cse);
  assign mux_279_nl = MUX_s_1_2_2(nor_2011_cse, mux_tmp_259, cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp);
  assign mux_280_nl = MUX_s_1_2_2(main_stage_v_1, (mux_279_nl), or_419_cse);
  assign and_161_nl = (IntShiftRightSat_49U_6U_17U_lor_4_lpi_1_dfm | cvt_3_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2)
      & mux_tmp_263;
  assign mux_283_nl = MUX_s_1_2_2(mux_tmp_263, (and_161_nl), or_461_cse);
  assign mux_284_nl = MUX_s_1_2_2(main_stage_v_2, (mux_283_nl), or_423_cse);
  assign mux_285_nl = MUX_s_1_2_2((mux_284_nl), (mux_280_nl), or_5189_cse);
  assign nor_1992_nl = ~((cfg_out_precision_1_sva_st_154[0]) | not_tmp_270);
  assign mux_288_nl = MUX_s_1_2_2(and_1078_cse, (nor_1992_nl), or_5189_cse);
  assign nor_1993_nl = ~(nor_2040_cse | (cfg_out_precision_1_sva_st_154[0]) | not_tmp_270);
  assign mux_289_nl = MUX_s_1_2_2((nor_1993_nl), (mux_288_nl), nor_63_cse);
  assign and_164_nl = main_stage_v_1 & cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp
      & mux_tmp_117;
  assign nor_1991_nl = ~((cfg_proc_precision_1_sva_st_101[1]) | (~ and_tmp_67));
  assign mux_290_nl = MUX_s_1_2_2((nor_1991_nl), and_tmp_67, cfg_proc_precision_1_sva_st_101[0]);
  assign and_166_nl = main_stage_v_2 & (mux_290_nl);
  assign mux_291_nl = MUX_s_1_2_2((and_166_nl), (and_164_nl), or_5189_cse);
  assign nor_1984_nl = ~((reg_cfg_proc_precision_1_sva_st_40_cse[1]) | (~ mux_tmp_294));
  assign mux_295_nl = MUX_s_1_2_2((nor_1984_nl), mux_tmp_294, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign mux_296_nl = MUX_s_1_2_2(main_stage_v_1, (mux_295_nl), or_513_cse);
  assign nor_1985_nl = ~((cfg_proc_precision_1_sva_st_89[1]) | (~ mux_tmp_299));
  assign mux_300_nl = MUX_s_1_2_2((nor_1985_nl), mux_tmp_299, cfg_proc_precision_1_sva_st_89[0]);
  assign mux_301_nl = MUX_s_1_2_2(main_stage_v_2, (mux_300_nl), or_451_cse);
  assign mux_302_nl = MUX_s_1_2_2((mux_301_nl), (mux_296_nl), or_5189_cse);
  assign mux_306_nl = MUX_s_1_2_2(nor_1980_cse, mux_tmp_305, cvt_4_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp);
  assign mux_307_nl = MUX_s_1_2_2(main_stage_v_1, (mux_306_nl), or_419_cse);
  assign mux_314_nl = MUX_s_1_2_2(mux_tmp_313, (~ or_tmp_533), cfg_proc_precision_1_sva_st_89[1]);
  assign mux_315_nl = MUX_s_1_2_2((mux_314_nl), mux_tmp_313, cfg_proc_precision_1_sva_st_89[0]);
  assign mux_316_nl = MUX_s_1_2_2((mux_315_nl), (mux_307_nl), or_5189_cse);
  assign and_168_nl = main_stage_v_2 & mux_tmp_321;
  assign mux_322_nl = MUX_s_1_2_2((and_168_nl), and_tmp_16, or_5189_cse);
  assign mux_327_nl = MUX_s_1_2_2(and_2230_cse, and_tmp_71, or_5189_cse);
  assign and_171_nl = cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2
      & main_stage_v_2 & mux_1126_cse;
  assign mux_328_nl = MUX_s_1_2_2((and_171_nl), and_tmp_71, or_5189_cse);
  assign mux_329_nl = MUX_s_1_2_2((mux_328_nl), (mux_327_nl), IntShiftRightSat_49U_6U_17U_lor_6_lpi_1_dfm);
  assign mux_332_nl = MUX_s_1_2_2(nor_2011_cse, mux_tmp_259, cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp);
  assign mux_333_nl = MUX_s_1_2_2(main_stage_v_1, (mux_332_nl), or_419_cse);
  assign and_172_nl = (IntShiftRightSat_49U_6U_17U_lor_6_lpi_1_dfm | cvt_5_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_st_2)
      & mux_tmp_263;
  assign mux_336_nl = MUX_s_1_2_2(mux_tmp_263, (and_172_nl), or_461_cse);
  assign mux_337_nl = MUX_s_1_2_2(main_stage_v_2, (mux_336_nl), or_423_cse);
  assign mux_338_nl = MUX_s_1_2_2((mux_337_nl), (mux_333_nl), or_5189_cse);
  assign and_2265_nl = (nor_2150_cse | (cfg_out_precision_1_sva_st_154!=2'b10)) &
      or_tmp_3768;
  assign mux_2175_nl = MUX_s_1_2_2((and_2265_nl), or_tmp_3768, nor_8_cse);
  assign or_4569_nl = nor_8_cse | nor_2150_cse | (cfg_out_precision_1_sva_st_154!=2'b10);
  assign mux_2176_nl = MUX_s_1_2_2((or_4569_nl), (mux_2175_nl), main_stage_v_2);
  assign nor_1962_nl = ~(nor_2040_cse | (cfg_out_precision_1_sva_st_154[0]) | not_tmp_119);
  assign mux_341_nl = MUX_s_1_2_2(and_2230_cse, (~ or_tmp_218), or_5189_cse);
  assign mux_342_nl = MUX_s_1_2_2((mux_341_nl), (nor_1962_nl), or_578_cse);
  assign and_173_nl = main_stage_v_1 & cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp
      & mux_344_cse;
  assign and_2229_nl = IntShiftRightSat_49U_6U_17U_lor_7_lpi_1_dfm & main_stage_v_2
      & mux_382_cse;
  assign mux_347_nl = MUX_s_1_2_2((and_2229_nl), and_174_cse, cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_svs_st_2);
  assign mux_348_nl = MUX_s_1_2_2((mux_347_nl), (and_173_nl), or_5189_cse);
  assign nor_1951_nl = ~((reg_cfg_proc_precision_1_sva_st_40_cse[1]) | (~ mux_tmp_351));
  assign mux_352_nl = MUX_s_1_2_2((nor_1951_nl), mux_tmp_351, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign mux_353_nl = MUX_s_1_2_2(main_stage_v_1, (mux_352_nl), or_513_cse);
  assign nor_1952_nl = ~((cfg_proc_precision_1_sva_st_89[1]) | (~ mux_tmp_356));
  assign mux_357_nl = MUX_s_1_2_2((nor_1952_nl), mux_tmp_356, cfg_proc_precision_1_sva_st_89[0]);
  assign mux_358_nl = MUX_s_1_2_2(main_stage_v_2, (mux_357_nl), or_451_cse);
  assign mux_359_nl = MUX_s_1_2_2((mux_358_nl), (mux_353_nl), or_5189_cse);
  assign mux_363_nl = MUX_s_1_2_2(nor_1980_cse, mux_tmp_305, cvt_6_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp);
  assign mux_364_nl = MUX_s_1_2_2(main_stage_v_1, (mux_363_nl), or_419_cse);
  assign mux_371_nl = MUX_s_1_2_2(mux_tmp_370, (~ or_tmp_533), cfg_proc_precision_1_sva_st_89[1]);
  assign mux_372_nl = MUX_s_1_2_2((mux_371_nl), mux_tmp_370, cfg_proc_precision_1_sva_st_89[0]);
  assign mux_373_nl = MUX_s_1_2_2((mux_372_nl), (mux_364_nl), or_5189_cse);
  assign and_179_nl = main_stage_v_1 & cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp
      & mux_344_cse;
  assign and_180_nl = or_4536_cse & main_stage_v_2 & mux_382_cse;
  assign mux_383_nl = MUX_s_1_2_2((and_180_nl), (and_179_nl), or_5189_cse);
  assign nor_1931_nl = ~((reg_cfg_proc_precision_1_sva_st_40_cse[1]) | (~ mux_tmp_386));
  assign mux_387_nl = MUX_s_1_2_2((nor_1931_nl), mux_tmp_386, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign mux_388_nl = MUX_s_1_2_2(main_stage_v_1, (mux_387_nl), or_513_cse);
  assign nor_1932_nl = ~((cfg_proc_precision_1_sva_st_89[1]) | (~ mux_tmp_391));
  assign mux_392_nl = MUX_s_1_2_2((nor_1932_nl), mux_tmp_391, cfg_proc_precision_1_sva_st_89[0]);
  assign mux_393_nl = MUX_s_1_2_2(main_stage_v_2, (mux_392_nl), or_451_cse);
  assign mux_394_nl = MUX_s_1_2_2((mux_393_nl), (mux_388_nl), or_5189_cse);
  assign mux_398_nl = MUX_s_1_2_2(nor_1980_cse, mux_tmp_305, cvt_7_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp);
  assign mux_399_nl = MUX_s_1_2_2(main_stage_v_1, (mux_398_nl), or_419_cse);
  assign mux_406_nl = MUX_s_1_2_2(mux_tmp_405, (~ or_tmp_533), cfg_proc_precision_1_sva_st_89[1]);
  assign mux_407_nl = MUX_s_1_2_2((mux_406_nl), mux_tmp_405, cfg_proc_precision_1_sva_st_89[0]);
  assign mux_408_nl = MUX_s_1_2_2((mux_407_nl), (mux_399_nl), or_5189_cse);
  assign and_182_nl = main_stage_v_1 & cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp
      & mux_344_cse;
  assign and_183_nl = or_4535_cse & main_stage_v_2 & mux_417_cse;
  assign mux_418_nl = MUX_s_1_2_2((and_183_nl), (and_182_nl), or_5189_cse);
  assign nor_1907_nl = ~((reg_cfg_proc_precision_1_sva_st_40_cse[1]) | (~ mux_tmp_422));
  assign mux_423_nl = MUX_s_1_2_2((nor_1907_nl), mux_tmp_422, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign mux_424_nl = MUX_s_1_2_2(main_stage_v_1, (mux_423_nl), or_513_cse);
  assign nor_1908_nl = ~((cfg_proc_precision_1_sva_st_89[1]) | (~ mux_tmp_428));
  assign mux_429_nl = MUX_s_1_2_2((nor_1908_nl), mux_tmp_428, cfg_proc_precision_1_sva_st_89[0]);
  assign mux_430_nl = MUX_s_1_2_2(main_stage_v_2, (mux_429_nl), or_451_cse);
  assign mux_431_nl = MUX_s_1_2_2((mux_430_nl), (mux_424_nl), or_5189_cse);
  assign mux_436_nl = MUX_s_1_2_2(nor_1898_cse, mux_tmp_435, cvt_8_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp);
  assign mux_437_nl = MUX_s_1_2_2(main_stage_v_1, (mux_436_nl), or_419_cse);
  assign and_185_nl = or_4535_cse & mux_tmp_441;
  assign mux_442_nl = MUX_s_1_2_2(mux_tmp_441, (and_185_nl), or_461_cse);
  assign mux_443_nl = MUX_s_1_2_2(main_stage_v_2, (mux_442_nl), or_423_cse);
  assign mux_444_nl = MUX_s_1_2_2((mux_443_nl), (mux_437_nl), or_5189_cse);
  assign mux_2183_nl = MUX_s_1_2_2(nor_2326_cse, or_tmp_3763, or_4559_cse);
  assign mux_2185_nl = MUX_s_1_2_2((mux_2183_nl), or_tmp_3763, nor_2150_cse);
  assign mux_2186_nl = MUX_s_1_2_2((mux_2185_nl), or_tmp_3763, nor_8_cse);
  assign mux_450_nl = MUX_s_1_2_2(and_178_itm, mux_tmp_129, or_5189_cse);
  assign mux_453_nl = MUX_s_1_2_2(and_2230_cse, and_tmp_18, or_5189_cse);
  assign mux_456_nl = MUX_s_1_2_2(and_tmp_94, and_tmp_93, or_5189_cse);
  assign and_2856_nl = and_tmp_93 & or_5189_cse;
  assign mux_458_nl = MUX_s_1_2_2((and_2856_nl), (mux_456_nl), cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_2);
  assign mux_461_nl = MUX_s_1_2_2(nor_2011_cse, mux_tmp_259, cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_tmp);
  assign mux_462_nl = MUX_s_1_2_2(main_stage_v_1, (mux_461_nl), or_419_cse);
  assign and_194_nl = cvt_9_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_1_svs_2
      & mux_tmp_263;
  assign mux_465_nl = MUX_s_1_2_2(mux_tmp_263, (and_194_nl), or_461_cse);
  assign mux_466_nl = MUX_s_1_2_2(main_stage_v_2, (mux_465_nl), or_423_cse);
  assign mux_467_nl = MUX_s_1_2_2((mux_466_nl), (mux_462_nl), or_5189_cse);
  assign mux_471_nl = MUX_s_1_2_2(and_tmp_94, nor_2004_cse, or_5189_cse);
  assign mux_472_nl = MUX_s_1_2_2(nor_2005_cse, (mux_471_nl), nor_63_cse);
  assign and_195_nl = main_stage_v_1 & cvt_10_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp
      & mux_474_cse;
  assign and_2221_nl = IntShiftRightSat_49U_6U_17U_lor_10_lpi_1_dfm & main_stage_v_2
      & mux_382_cse;
  assign mux_477_nl = MUX_s_1_2_2((and_2221_nl), and_174_cse, IntShiftRightSat_49U_6U_17U_lor_11_lpi_1_dfm);
  assign mux_478_nl = MUX_s_1_2_2((mux_477_nl), (and_195_nl), or_5189_cse);
  assign nor_1868_nl = ~((reg_cfg_proc_precision_1_sva_st_40_cse[1]) | (~ mux_tmp_481));
  assign mux_482_nl = MUX_s_1_2_2((nor_1868_nl), mux_tmp_481, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign mux_483_nl = MUX_s_1_2_2(main_stage_v_1, (mux_482_nl), or_513_cse);
  assign nor_1869_nl = ~((cfg_proc_precision_1_sva_st_89[1]) | (~ mux_tmp_487));
  assign mux_488_nl = MUX_s_1_2_2((nor_1869_nl), mux_tmp_487, cfg_proc_precision_1_sva_st_89[0]);
  assign mux_489_nl = MUX_s_1_2_2(main_stage_v_2, (mux_488_nl), or_451_cse);
  assign mux_490_nl = MUX_s_1_2_2((mux_489_nl), (mux_483_nl), or_5189_cse);
  assign mux_494_nl = MUX_s_1_2_2(nor_1980_cse, mux_tmp_305, cvt_10_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp);
  assign mux_495_nl = MUX_s_1_2_2(main_stage_v_1, (mux_494_nl), or_419_cse);
  assign mux_503_nl = MUX_s_1_2_2(mux_tmp_502, (~ or_tmp_533), cfg_proc_precision_1_sva_st_89[1]);
  assign mux_504_nl = MUX_s_1_2_2((mux_503_nl), mux_tmp_502, cfg_proc_precision_1_sva_st_89[0]);
  assign mux_505_nl = MUX_s_1_2_2((mux_504_nl), (mux_495_nl), or_5189_cse);
  assign and_199_nl = main_stage_v_1 & cvt_11_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp
      & mux_474_cse;
  assign and_2217_nl = IntShiftRightSat_49U_6U_17U_lor_12_lpi_1_dfm & main_stage_v_2
      & mux_382_cse;
  assign mux_515_nl = MUX_s_1_2_2((and_2217_nl), and_174_cse, IntShiftRightSat_49U_6U_17U_lor_2_lpi_1_dfm);
  assign mux_516_nl = MUX_s_1_2_2((mux_515_nl), (and_199_nl), or_5189_cse);
  assign nor_1847_nl = ~((reg_cfg_proc_precision_1_sva_st_40_cse[1]) | (~ mux_tmp_519));
  assign mux_520_nl = MUX_s_1_2_2((nor_1847_nl), mux_tmp_519, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign mux_521_nl = MUX_s_1_2_2(main_stage_v_1, (mux_520_nl), or_513_cse);
  assign nor_1848_nl = ~((cfg_proc_precision_1_sva_st_89[1]) | (~ mux_tmp_525));
  assign mux_526_nl = MUX_s_1_2_2((nor_1848_nl), mux_tmp_525, cfg_proc_precision_1_sva_st_89[0]);
  assign mux_527_nl = MUX_s_1_2_2(main_stage_v_2, (mux_526_nl), or_451_cse);
  assign mux_528_nl = MUX_s_1_2_2((mux_527_nl), (mux_521_nl), or_5189_cse);
  assign mux_532_nl = MUX_s_1_2_2(nor_1980_cse, mux_tmp_305, cvt_11_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp);
  assign mux_533_nl = MUX_s_1_2_2(main_stage_v_1, (mux_532_nl), or_419_cse);
  assign mux_542_nl = MUX_s_1_2_2(mux_tmp_541, (~ or_tmp_533), cfg_proc_precision_1_sva_st_89[1]);
  assign mux_543_nl = MUX_s_1_2_2((mux_542_nl), mux_tmp_541, cfg_proc_precision_1_sva_st_89[0]);
  assign mux_544_nl = MUX_s_1_2_2((mux_543_nl), (mux_533_nl), or_5189_cse);
  assign and_203_nl = main_stage_v_1 & cvt_12_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp
      & mux_474_cse;
  assign and_2213_nl = IntShiftRightSat_49U_6U_17U_lor_13_lpi_1_dfm & mux_417_cse;
  assign mux_555_nl = MUX_s_1_2_2((and_2213_nl), mux_417_cse, IsNaN_5U_10U_IsNaN_5U_10U_nand_14_itm_2);
  assign and_205_nl = main_stage_v_2 & (mux_555_nl);
  assign mux_556_nl = MUX_s_1_2_2((and_205_nl), (and_203_nl), or_5189_cse);
  assign nor_1822_nl = ~((reg_cfg_proc_precision_1_sva_st_40_cse[1]) | (~ mux_tmp_560));
  assign mux_561_nl = MUX_s_1_2_2((nor_1822_nl), mux_tmp_560, reg_cfg_proc_precision_1_sva_st_40_cse[0]);
  assign mux_562_nl = MUX_s_1_2_2(main_stage_v_1, (mux_561_nl), or_513_cse);
  assign nor_1823_nl = ~((cfg_proc_precision_1_sva_st_89[1]) | (~ mux_tmp_566));
  assign mux_567_nl = MUX_s_1_2_2((nor_1823_nl), mux_tmp_566, cfg_proc_precision_1_sva_st_89[0]);
  assign mux_568_nl = MUX_s_1_2_2(main_stage_v_2, (mux_567_nl), or_451_cse);
  assign mux_569_nl = MUX_s_1_2_2((mux_568_nl), (mux_562_nl), or_5189_cse);
  assign mux_574_nl = MUX_s_1_2_2(nor_1898_cse, mux_tmp_435, cvt_12_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp);
  assign mux_575_nl = MUX_s_1_2_2(main_stage_v_1, (mux_574_nl), or_419_cse);
  assign nor_1814_nl = ~((cfg_proc_precision_1_sva_st_89[1]) | (~ mux_tmp_580));
  assign mux_581_nl = MUX_s_1_2_2((nor_1814_nl), mux_tmp_580, cfg_proc_precision_1_sva_st_89[0]);
  assign mux_582_nl = MUX_s_1_2_2(main_stage_v_2, (mux_581_nl), or_423_cse);
  assign mux_583_nl = MUX_s_1_2_2((mux_582_nl), (mux_575_nl), or_5189_cse);
  assign and_210_nl = main_stage_v_1 & cvt_13_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp
      & mux_474_cse;
  assign nor_1809_nl = ~((cfg_proc_precision_1_sva_st_65[1]) | (~ mux_tmp_592));
  assign mux_593_nl = MUX_s_1_2_2((nor_1809_nl), mux_tmp_592, cfg_proc_precision_1_sva_st_65[0]);
  assign and_212_nl = main_stage_v_2 & (mux_593_nl);
  assign mux_594_nl = MUX_s_1_2_2((and_212_nl), (and_210_nl), or_5189_cse);
  assign nor_1800_nl = ~(((cfg_out_precision_1_sva_st_154[1]) & cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp)
      | (cfg_out_precision_1_sva_st_154[0]) | (~ mux_tmp_597));
  assign mux_598_nl = MUX_s_1_2_2((nor_1800_nl), mux_tmp_597, cvt_13_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp);
  assign mux_599_nl = MUX_s_1_2_2(main_stage_v_1, (mux_598_nl), or_513_cse);
  assign nor_1801_nl = ~((cfg_proc_precision_1_sva_st_65[1]) | (~ mux_tmp_602));
  assign mux_603_nl = MUX_s_1_2_2((nor_1801_nl), mux_tmp_602, cfg_proc_precision_1_sva_st_65[0]);
  assign mux_604_nl = MUX_s_1_2_2(main_stage_v_2, (mux_603_nl), or_451_cse);
  assign mux_605_nl = MUX_s_1_2_2((mux_604_nl), (mux_599_nl), or_5189_cse);
  assign nor_1793_nl = ~((cfg_out_precision_1_sva_st_154!=2'b00) | (~ mux_tmp_597));
  assign mux_609_nl = MUX_s_1_2_2((nor_1793_nl), mux_tmp_597, cvt_13_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_2_tmp);
  assign mux_610_nl = MUX_s_1_2_2(main_stage_v_1, (mux_609_nl), or_419_cse);
  assign nor_1794_nl = ~((cfg_proc_precision_1_sva_st_65[1]) | (~ mux_tmp_614));
  assign mux_615_nl = MUX_s_1_2_2((nor_1794_nl), mux_tmp_614, cfg_proc_precision_1_sva_st_65[0]);
  assign mux_616_nl = MUX_s_1_2_2(main_stage_v_2, (mux_615_nl), or_423_cse);
  assign mux_617_nl = MUX_s_1_2_2((mux_616_nl), (mux_610_nl), or_5189_cse);
  assign and_213_nl = main_stage_v_1 & cvt_14_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp
      & mux_474_cse;
  assign and_2203_nl = IntShiftRightSat_49U_6U_17U_lor_15_lpi_1_dfm & mux_417_cse;
  assign mux_629_nl = MUX_s_1_2_2((and_2203_nl), mux_417_cse, IsNaN_5U_10U_nor_1_itm_2);
  assign and_215_nl = main_stage_v_2 & (mux_629_nl);
  assign mux_630_nl = MUX_s_1_2_2((and_215_nl), (and_213_nl), or_5189_cse);
  assign mux_635_nl = MUX_s_1_2_2(nor_1772_cse, mux_tmp_634, cvt_14_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp);
  assign or_961_nl = (cfg_out_precision_1_sva_st_154!=2'b00);
  assign mux_636_nl = MUX_s_1_2_2(main_stage_v_1, (mux_635_nl), or_961_nl);
  assign nor_1773_nl = ~((cfg_proc_precision_1_sva_st_65[1]) | (~ mux_tmp_641));
  assign mux_642_nl = MUX_s_1_2_2((nor_1773_nl), mux_tmp_641, cfg_proc_precision_1_sva_st_65[0]);
  assign mux_643_nl = MUX_s_1_2_2(main_stage_v_2, (mux_642_nl), or_425_cse);
  assign mux_644_nl = MUX_s_1_2_2((mux_643_nl), (mux_636_nl), or_5189_cse);
  assign mux_2210_nl = MUX_s_1_2_2(mux_tmp_2206, (~ mux_tmp_2203), cfg_proc_precision_1_sva_st_64[1]);
  assign mux_2211_nl = MUX_s_1_2_2((mux_2210_nl), mux_tmp_2206, cfg_proc_precision_1_sva_st_64[0]);
  assign mux_2212_nl = MUX_s_1_2_2((~ mux_tmp_2203), (mux_2211_nl), or_183_cse_1);
  assign and_2487_nl = (cfg_out_precision_1_sva_st_154[1]) & main_stage_v_1;
  assign mux_2213_nl = MUX_s_1_2_2((~ mux_tmp_2203), (mux_2212_nl), and_2487_nl);
  assign mux_2214_nl = MUX_s_1_2_2((mux_2213_nl), (~ mux_tmp_2203), or_4559_cse);
  assign and_216_nl = main_stage_v_1 & cvt_15_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp
      & mux_474_cse;
  assign and_2201_nl = IntShiftRightSat_49U_6U_17U_lor_16_lpi_1_dfm & mux_417_cse;
  assign mux_670_nl = MUX_s_1_2_2((and_2201_nl), mux_417_cse, IsNaN_5U_10U_nor_14_itm_2);
  assign and_218_nl = main_stage_v_2 & (mux_670_nl);
  assign mux_671_nl = MUX_s_1_2_2((and_218_nl), (and_216_nl), or_5189_cse);
  assign nor_1745_nl = ~(((cfg_out_precision_1_sva_st_154[1]) & cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp)
      | (cfg_out_precision_1_sva_st_154[0]) | (~ mux_tmp_634));
  assign mux_676_nl = MUX_s_1_2_2((nor_1745_nl), mux_tmp_634, cvt_15_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp);
  assign mux_677_nl = MUX_s_1_2_2(main_stage_v_1, (mux_676_nl), or_513_cse);
  assign nor_1746_nl = ~((cfg_proc_precision_1_sva_st_65[1]) | (~ mux_tmp_681));
  assign mux_682_nl = MUX_s_1_2_2((nor_1746_nl), mux_tmp_681, cfg_proc_precision_1_sva_st_65[0]);
  assign mux_683_nl = MUX_s_1_2_2(main_stage_v_2, (mux_682_nl), or_451_cse);
  assign mux_684_nl = MUX_s_1_2_2((mux_683_nl), (mux_677_nl), or_5189_cse);
  assign mux_689_nl = MUX_s_1_2_2(nor_1772_cse, mux_tmp_634, cvt_15_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_3_tmp);
  assign mux_690_nl = MUX_s_1_2_2(main_stage_v_1, (mux_689_nl), or_419_cse);
  assign nor_1737_nl = ~((cfg_proc_precision_1_sva_st_65[1]) | (~ mux_tmp_695));
  assign mux_696_nl = MUX_s_1_2_2((nor_1737_nl), mux_tmp_695, cfg_proc_precision_1_sva_st_65[0]);
  assign mux_697_nl = MUX_s_1_2_2(main_stage_v_2, (mux_696_nl), or_423_cse);
  assign mux_698_nl = MUX_s_1_2_2((mux_697_nl), (mux_690_nl), or_5189_cse);
  assign nor_2290_nl = ~((cfg_out_precision_1_sva_st_154[1]) | (~ or_tmp_3840));
  assign mux_2215_nl = MUX_s_1_2_2((nor_2290_nl), or_tmp_3840, or_4559_cse);
  assign mux_2216_nl = MUX_s_1_2_2((mux_2215_nl), or_tmp_3840, nor_2150_cse);
  assign mux_2217_nl = MUX_s_1_2_2(or_tmp_3840, (mux_2216_nl), or_183_cse_1);
  assign mux_2218_nl = MUX_s_1_2_2((mux_2217_nl), or_tmp_3840, nor_8_cse);
  assign and_219_nl = main_stage_v_1 & cvt_16_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_4_tmp
      & mux_344_cse;
  assign and_2196_nl = IntShiftRightSat_49U_6U_17U_lor_lpi_1_dfm & mux_417_cse;
  assign mux_714_nl = MUX_s_1_2_2((and_2196_nl), mux_417_cse, IsNaN_5U_10U_nor_itm_2);
  assign and_221_nl = main_stage_v_2 & (mux_714_nl);
  assign mux_715_nl = MUX_s_1_2_2((and_221_nl), (and_219_nl), or_5189_cse);
  assign nor_1708_nl = ~(((cfg_out_precision_1_sva_st_154[1]) & cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_tmp)
      | (cfg_out_precision_1_sva_st_154[0]) | (~ mux_tmp_720));
  assign mux_721_nl = MUX_s_1_2_2((nor_1708_nl), mux_tmp_720, cvt_16_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_4_tmp);
  assign mux_722_nl = MUX_s_1_2_2(main_stage_v_1, (mux_721_nl), or_513_cse);
  assign nor_1709_nl = ~((cfg_proc_precision_1_sva_st_65[1]) | (~ mux_tmp_727));
  assign mux_728_nl = MUX_s_1_2_2((nor_1709_nl), mux_tmp_727, cfg_proc_precision_1_sva_st_65[0]);
  assign mux_729_nl = MUX_s_1_2_2(main_stage_v_2, (mux_728_nl), or_451_cse);
  assign mux_730_nl = MUX_s_1_2_2((mux_729_nl), (mux_722_nl), or_5189_cse);
  assign nor_1697_nl = ~((cfg_out_precision_1_sva_st_154!=2'b00) | (~ mux_tmp_720));
  assign mux_736_nl = MUX_s_1_2_2((nor_1697_nl), mux_tmp_720, cvt_16_IntShiftRightSat_49U_6U_17U_IntShiftRightSat_49U_6U_17U_oelse_IntShiftRightSat_49U_6U_17U_if_unequal_4_tmp);
  assign mux_737_nl = MUX_s_1_2_2(main_stage_v_1, (mux_736_nl), or_419_cse);
  assign nor_1698_nl = ~((cfg_proc_precision_1_sva_st_65[1]) | (~ mux_tmp_743));
  assign mux_744_nl = MUX_s_1_2_2((nor_1698_nl), mux_tmp_743, cfg_proc_precision_1_sva_st_65[0]);
  assign mux_745_nl = MUX_s_1_2_2(main_stage_v_2, (mux_744_nl), or_423_cse);
  assign mux_746_nl = MUX_s_1_2_2((mux_745_nl), (mux_737_nl), or_5189_cse);
  assign nor_2287_nl = ~((cfg_out_precision_1_sva_st_154[1]) | (~ or_tmp_3849));
  assign mux_2219_nl = MUX_s_1_2_2((nor_2287_nl), or_tmp_3849, or_4559_cse);
  assign mux_2221_nl = MUX_s_1_2_2((mux_2219_nl), or_tmp_3849, nor_2150_cse);
  assign mux_2222_nl = MUX_s_1_2_2(or_tmp_3849, (mux_2221_nl), or_183_cse_1);
  assign mux_2223_nl = MUX_s_1_2_2((mux_2222_nl), or_tmp_3849, nor_8_cse);
  assign mux_792_nl = MUX_s_1_2_2((~ or_tmp_306), and_tmp_8, or_5189_cse);
  assign and_136_nl = main_stage_v_2 & or_tmp_389;
  assign mux_793_nl = MUX_s_1_2_2((and_136_nl), and_tmp_8, or_5189_cse);
  assign mux_794_nl = MUX_s_1_2_2((mux_793_nl), (mux_792_nl), nor_151_cse);
  assign nl_cvt_10_IntSaturation_17U_8U_if_acc_2_nl = conv_s2u_10_11({(~ IntShiftRightSat_49U_6U_17U_o_16_10_sva_2)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_2[14:6]))}) + 11'b1;
  assign cvt_10_IntSaturation_17U_8U_if_acc_2_nl = nl_cvt_10_IntSaturation_17U_8U_if_acc_2_nl[10:0];
  assign nl_cvt_2_IntSaturation_17U_8U_if_acc_1_nl = conv_s2u_10_11({(~ IntShiftRightSat_49U_6U_17U_o_16_2_sva_2)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_2[14:6]))}) + 11'b1;
  assign cvt_2_IntSaturation_17U_8U_if_acc_1_nl = nl_cvt_2_IntSaturation_17U_8U_if_acc_1_nl[10:0];
  assign nl_cvt_4_IntSaturation_17U_8U_if_acc_2_nl = conv_s2u_10_11({(~ IntShiftRightSat_49U_6U_17U_o_16_4_sva_2)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_2[14:6]))}) + 11'b1;
  assign cvt_4_IntSaturation_17U_8U_if_acc_2_nl = nl_cvt_4_IntSaturation_17U_8U_if_acc_2_nl[10:0];
  assign nl_cvt_6_IntSaturation_17U_8U_if_acc_2_nl = conv_s2u_10_11({(~ IntShiftRightSat_49U_6U_17U_o_16_6_sva_2)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_2[14:6]))}) + 11'b1;
  assign cvt_6_IntSaturation_17U_8U_if_acc_2_nl = nl_cvt_6_IntSaturation_17U_8U_if_acc_2_nl[10:0];
  assign nl_cvt_7_IntSaturation_17U_8U_if_acc_2_nl = conv_s2u_10_11({(~ IntShiftRightSat_49U_6U_17U_o_16_7_sva_2)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_2[14:6]))}) + 11'b1;
  assign cvt_7_IntSaturation_17U_8U_if_acc_2_nl = nl_cvt_7_IntSaturation_17U_8U_if_acc_2_nl[10:0];
  assign nl_cvt_16_IntSaturation_17U_8U_if_acc_4_nl = conv_s2u_10_11({(~ IntShiftRightSat_49U_6U_17U_o_16_sva_2)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_sva_2[14:6]))}) + 11'b1;
  assign cvt_16_IntSaturation_17U_8U_if_acc_4_nl = nl_cvt_16_IntSaturation_17U_8U_if_acc_4_nl[10:0];
  assign nl_cvt_8_IntSaturation_17U_8U_if_acc_3_nl = conv_s2u_10_11({(~ IntShiftRightSat_49U_6U_17U_o_16_8_sva_2)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_2[14:6]))}) + 11'b1;
  assign cvt_8_IntSaturation_17U_8U_if_acc_3_nl = nl_cvt_8_IntSaturation_17U_8U_if_acc_3_nl[10:0];
  assign nl_cvt_15_IntSaturation_17U_8U_if_acc_3_nl = conv_s2u_10_11({(~ IntShiftRightSat_49U_6U_17U_o_16_15_sva_2)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_2[14:6]))}) + 11'b1;
  assign cvt_15_IntSaturation_17U_8U_if_acc_3_nl = nl_cvt_15_IntSaturation_17U_8U_if_acc_3_nl[10:0];
  assign nl_cvt_13_IntSaturation_17U_8U_if_acc_2_nl = conv_s2u_10_11({(~ IntShiftRightSat_49U_6U_17U_o_16_13_sva_2)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_2[14:6]))}) + 11'b1;
  assign cvt_13_IntSaturation_17U_8U_if_acc_2_nl = nl_cvt_13_IntSaturation_17U_8U_if_acc_2_nl[10:0];
  assign nl_cvt_11_IntSaturation_17U_8U_if_acc_2_nl = conv_s2u_10_11({(~ IntShiftRightSat_49U_6U_17U_o_16_11_sva_2)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_2[14:6]))}) + 11'b1;
  assign cvt_11_IntSaturation_17U_8U_if_acc_2_nl = nl_cvt_11_IntSaturation_17U_8U_if_acc_2_nl[10:0];
  assign nl_cvt_12_IntSaturation_17U_8U_if_acc_3_nl = conv_s2u_10_11({(~ IntShiftRightSat_49U_6U_17U_o_16_12_sva_2)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_2[14:6]))}) + 11'b1;
  assign cvt_12_IntSaturation_17U_8U_if_acc_3_nl = nl_cvt_12_IntSaturation_17U_8U_if_acc_3_nl[10:0];
  assign nor_1667_nl = ~((~(nor_1056_cse | (chn_idata_data_sva_2_47_31_1[0]))) |
      (cfg_out_precision_1_sva_st_113!=2'b01) | (~ main_stage_v_2) | cfg_mode_eql_1_sva_5);
  assign mux_805_nl = MUX_s_1_2_2((nor_1667_nl), nor_1666_cse, cvt_unequal_tmp_20);
  assign nor_1670_nl = ~((~ (chn_idata_data_sva_2_47_31_1[0])) | (~ main_stage_v_2)
      | cfg_mode_eql_1_sva_5);
  assign mux_806_nl = MUX_s_1_2_2((nor_1670_nl), nor_1669_cse, cvt_unequal_tmp_20);
  assign mux_807_nl = MUX_s_1_2_2((mux_806_nl), (mux_805_nl), nor_50_cse);
  assign nand_208_nl = ~((cvt_1_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_svs_2
      | (chn_idata_data_sva_3_47_31_1[0])) & or_1159_cse);
  assign mux_808_nl = MUX_s_1_2_2((nand_208_nl), or_1159_cse, cvt_unequal_tmp_21);
  assign or_4532_nl = (~(cvt_1_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_svs_2
      | (chn_idata_data_sva_3_47_31_1[0]))) | or_1159_cse;
  assign mux_809_nl = MUX_s_1_2_2((or_4532_nl), nor_1672_cse, cvt_unequal_tmp_21);
  assign mux_810_nl = MUX_s_1_2_2((mux_809_nl), (mux_808_nl), or_1157_cse);
  assign nor_1671_nl = ~((~ main_stage_v_3) | cfg_mode_eql_1_sva_6 | (mux_810_nl));
  assign mux_811_nl = MUX_s_1_2_2((nor_1671_nl), (mux_807_nl), or_5189_cse);
  assign nor_1665_nl = ~((~ cvt_1_FpFloatToInt_16U_5U_10U_if_acc_itm_11_1) | (cfg_proc_precision_1_sva_st_65!=2'b10)
      | (cfg_out_precision_1_sva_st_113!=2'b01));
  assign mux_812_nl = MUX_s_1_2_2((nor_1665_nl), nor_1664_cse, or_309_cse);
  assign and_227_nl = main_stage_v_2 & (cfg_mode_eql_1_sva_5 | (~(cvt_unequal_tmp_20
      | (mux_812_nl))));
  assign nand_2_nl = ~(cvt_1_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_svs_2
      & (~ mux_813_cse));
  assign mux_814_nl = MUX_s_1_2_2((nand_2_nl), cfg_mode_eql_1_sva_6, cvt_unequal_tmp_21);
  assign and_228_nl = main_stage_v_3 & (mux_814_nl);
  assign mux_815_nl = MUX_s_1_2_2((and_228_nl), (and_227_nl), or_5189_cse);
  assign nor_1658_nl = ~((~ cvt_2_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1) | (cfg_proc_precision_1_sva_st_65!=2'b10)
      | (cfg_out_precision_1_sva_st_113!=2'b01));
  assign mux_819_nl = MUX_s_1_2_2((nor_1658_nl), nor_1664_cse, or_309_cse);
  assign and_229_nl = main_stage_v_2 & (cfg_mode_eql_1_sva_5 | (~(cvt_unequal_tmp_20
      | (mux_819_nl))));
  assign nand_3_nl = ~(cvt_2_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2
      & (~ mux_813_cse));
  assign mux_821_nl = MUX_s_1_2_2((nand_3_nl), cfg_mode_eql_1_sva_6, cvt_unequal_tmp_21);
  assign and_230_nl = main_stage_v_3 & (mux_821_nl);
  assign mux_822_nl = MUX_s_1_2_2((and_230_nl), (and_229_nl), or_5189_cse);
  assign or_1201_nl = cvt_1_FpMantRNE_17U_11U_else_and_svs | (cfg_out_precision_1_sva_st_113!=2'b10)
      | (~ FpIntToFloat_17U_5U_10U_else_unequal_tmp);
  assign nand_4_nl = ~(or_1202_cse & (~((~(cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_1_itm_4
      | (~ cvt_1_FpMantRNE_17U_11U_else_and_tmp))) | (cfg_out_precision_1_sva_st_113!=2'b10))));
  assign mux_823_nl = MUX_s_1_2_2((nand_4_nl), (or_1201_nl), cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_svs_st_2);
  assign and_2191_nl = IsNaN_5U_10U_IsNaN_5U_10U_nand_1_itm_2 & cvt_unequal_tmp_20;
  assign mux_825_nl = MUX_s_1_2_2((mux_823_nl), or_1198_cse, and_2191_nl);
  assign mux_826_nl = MUX_s_1_2_2((mux_825_nl), or_1196_cse, nor_50_cse);
  assign nor_1653_nl = ~((~ main_stage_v_2) | cfg_mode_eql_1_sva_5 | (mux_826_nl));
  assign or_1209_nl = (cfg_out_precision_1_sva_st_136!=2'b10) | FpIntToFloat_17U_5U_10U_is_inf_1_lpi_1_dfm_6
      | (cfg_out_precision_1_sva_6[0]) | nand_207_cse;
  assign mux_828_nl = MUX_s_1_2_2(mux_827_cse, (or_1209_nl), cvt_unequal_tmp_21);
  assign nor_1655_nl = ~((~ main_stage_v_3) | cfg_mode_eql_1_sva_6 | (mux_828_nl));
  assign mux_829_nl = MUX_s_1_2_2((nor_1655_nl), (nor_1653_nl), or_5189_cse);
  assign and_2357_nl = cvt_unequal_tmp_20 & (nor_2219_cse | (cfg_out_precision_1_sva_st_113!=2'b10));
  assign mux_2224_nl = MUX_s_1_2_2((and_2357_nl), or_4709_cse, nor_50_cse);
  assign nor_1652_nl = ~((~ cvt_3_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1) | (cfg_proc_precision_1_sva_st_65!=2'b10)
      | (cfg_out_precision_1_sva_st_113!=2'b01));
  assign mux_830_nl = MUX_s_1_2_2((nor_1652_nl), nor_1664_cse, or_309_cse);
  assign and_233_nl = main_stage_v_2 & (cfg_mode_eql_1_sva_5 | (~(cvt_unequal_tmp_20
      | (mux_830_nl))));
  assign nand_5_nl = ~(cvt_3_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2
      & (~ mux_813_cse));
  assign mux_832_nl = MUX_s_1_2_2((nand_5_nl), cfg_mode_eql_1_sva_6, cvt_unequal_tmp_21);
  assign and_234_nl = main_stage_v_3 & (mux_832_nl);
  assign mux_833_nl = MUX_s_1_2_2((and_234_nl), (and_233_nl), or_5189_cse);
  assign nl_cvt_3_FpMantRNE_17U_11U_else_acc_1_nl = (cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[15:6])
      + conv_u2u_1_10(FpMantRNE_17U_11U_else_carry_3_sva);
  assign cvt_3_FpMantRNE_17U_11U_else_acc_1_nl = nl_cvt_3_FpMantRNE_17U_11U_else_acc_1_nl[9:0];
  assign FpIntToFloat_17U_5U_10U_if_not_182_nl = ~ cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2;
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_and_7_nl = MUX_v_10_2_2(10'b0000000000,
      (cvt_3_FpMantRNE_17U_11U_else_acc_1_nl), (FpIntToFloat_17U_5U_10U_if_not_182_nl));
  assign nor_1649_nl = ~((~ cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1) | (cfg_proc_precision_1_sva_st_65!=2'b10)
      | (cfg_out_precision_1_sva_st_113!=2'b01));
  assign mux_834_nl = MUX_s_1_2_2((nor_1649_nl), nor_1664_cse, or_309_cse);
  assign and_235_nl = main_stage_v_2 & (cfg_mode_eql_1_sva_5 | (~(cvt_unequal_tmp_20
      | (mux_834_nl))));
  assign nand_6_nl = ~(cvt_4_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2
      & (~ mux_813_cse));
  assign mux_836_nl = MUX_s_1_2_2((nand_6_nl), cfg_mode_eql_1_sva_6, cvt_unequal_tmp_21);
  assign and_236_nl = main_stage_v_3 & (mux_836_nl);
  assign mux_837_nl = MUX_s_1_2_2((and_236_nl), (and_235_nl), or_5189_cse);
  assign FpFloatToInt_16U_5U_10U_and_37_nl = (~ (chn_idata_data_sva_2_143_127_1[0]))
      & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_3_m1c & and_dcpl_408;
  assign FpFloatToInt_16U_5U_10U_and_38_nl = (chn_idata_data_sva_2_143_127_1[0])
      & FpFloatToInt_16U_5U_10U_FpFloatToInt_16U_5U_10U_nor_3_m1c & and_dcpl_408;
  assign FpFloatToInt_16U_5U_10U_and_7_nl = cvt_4_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1
      & (~ IsNaN_5U_10U_land_4_lpi_1_dfm_4) & and_dcpl_408;
  assign FpFloatToInt_16U_5U_10U_o_int_and_28_nl = IsNaN_5U_10U_land_4_lpi_1_dfm_4
      & and_dcpl_408;
  assign nor_1646_nl = ~((~ cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1) | (cfg_proc_precision_1_sva_st_65!=2'b10)
      | (cfg_out_precision_1_sva_st_113!=2'b01));
  assign mux_838_nl = MUX_s_1_2_2((nor_1646_nl), nor_1664_cse, or_309_cse);
  assign and_237_nl = main_stage_v_2 & (cfg_mode_eql_1_sva_5 | (~(cvt_unequal_tmp_20
      | (mux_838_nl))));
  assign nand_7_nl = ~(cvt_15_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2
      & (~ mux_813_cse));
  assign mux_840_nl = MUX_s_1_2_2((nand_7_nl), cfg_mode_eql_1_sva_6, cvt_unequal_tmp_21);
  assign and_238_nl = main_stage_v_3 & (mux_840_nl);
  assign mux_841_nl = MUX_s_1_2_2((and_238_nl), (and_237_nl), or_5189_cse);
  assign nor_1636_nl = ~((~ (chn_idata_data_sva_2_175_159_1[0])) | (cfg_out_precision_1_sva_st_113!=2'b01)
      | (~ main_stage_v_2) | cfg_mode_eql_1_sva_5);
  assign nor_1637_nl = ~((~(cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1 | (chn_idata_data_sva_2_175_159_1[0])))
      | (cfg_out_precision_1_sva_st_113!=2'b01) | (~ main_stage_v_2) | cfg_mode_eql_1_sva_5);
  assign mux_842_nl = MUX_s_1_2_2((nor_1637_nl), (nor_1636_nl), or_300_cse);
  assign mux_843_nl = MUX_s_1_2_2((mux_842_nl), nor_1666_cse, cvt_unequal_tmp_20);
  assign nor_1640_nl = ~((~ (chn_idata_data_sva_2_175_159_1[0])) | (~ main_stage_v_2)
      | cfg_mode_eql_1_sva_5);
  assign mux_844_nl = MUX_s_1_2_2((nor_1640_nl), nor_1669_cse, cvt_unequal_tmp_20);
  assign mux_845_nl = MUX_s_1_2_2((mux_844_nl), (mux_843_nl), nor_50_cse);
  assign nand_206_nl = ~((cvt_5_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2
      | (chn_idata_data_sva_3_175_159_1[0])) & or_1159_cse);
  assign mux_846_nl = MUX_s_1_2_2((nand_206_nl), or_1159_cse, cvt_unequal_tmp_21);
  assign or_4530_nl = (~(cvt_5_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2
      | (chn_idata_data_sva_3_175_159_1[0]))) | or_1159_cse;
  assign mux_847_nl = MUX_s_1_2_2((or_4530_nl), nor_1672_cse, cvt_unequal_tmp_21);
  assign mux_848_nl = MUX_s_1_2_2((mux_847_nl), (mux_846_nl), or_1157_cse);
  assign nor_1641_nl = ~((~ main_stage_v_3) | cfg_mode_eql_1_sva_6 | (mux_848_nl));
  assign mux_849_nl = MUX_s_1_2_2((nor_1641_nl), (mux_845_nl), or_5189_cse);
  assign nor_1634_nl = ~((~ cvt_5_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1) | (cfg_proc_precision_1_sva_st_65!=2'b10)
      | (cfg_out_precision_1_sva_st_113!=2'b01));
  assign mux_850_nl = MUX_s_1_2_2((nor_1634_nl), nor_1664_cse, or_300_cse);
  assign and_240_nl = main_stage_v_2 & (cfg_mode_eql_1_sva_5 | (~(cvt_unequal_tmp_20
      | (mux_850_nl))));
  assign nand_9_nl = ~(cvt_5_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2
      & (~ mux_813_cse));
  assign mux_852_nl = MUX_s_1_2_2((nand_9_nl), cfg_mode_eql_1_sva_6, cvt_unequal_tmp_21);
  assign and_241_nl = main_stage_v_3 & (mux_852_nl);
  assign mux_853_nl = MUX_s_1_2_2((and_241_nl), (and_240_nl), or_5189_cse);
  assign nor_1625_nl = ~(cvt_16_FpFloatToInt_16U_5U_10U_if_acc_4_itm_11_1 | chn_idata_data_sva_2_511_1
      | (~ main_stage_v_2) | cvt_unequal_tmp_20 | cfg_mode_eql_1_sva_5);
  assign mux_854_nl = MUX_s_1_2_2((nor_1625_nl), nor_1624_cse, or_309_cse);
  assign mux_855_nl = MUX_s_1_2_2(nor_1626_cse, (mux_854_nl), nor_2285_cse);
  assign mux_856_nl = MUX_s_1_2_2(nor_1624_cse, (mux_855_nl), nor_50_cse);
  assign nor_1628_nl = ~(nor_1629_cse | (~ main_stage_v_3) | cvt_unequal_tmp_21 |
      cfg_mode_eql_1_sva_6);
  assign mux_857_nl = MUX_s_1_2_2(nor_1630_cse, (nor_1628_nl), nor_1672_cse);
  assign or_1280_nl = cvt_16_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_4_svs_2
      | IntSaturation_17U_16U_IntSaturation_17U_16U_or_1_itm_3;
  assign mux_858_nl = MUX_s_1_2_2(nor_1630_cse, (mux_857_nl), or_1280_nl);
  assign mux_859_nl = MUX_s_1_2_2((mux_858_nl), (mux_856_nl), or_5189_cse);
  assign nor_1623_nl = ~((~ cvt_14_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1) | (cfg_proc_precision_1_sva_st_65!=2'b10)
      | (cfg_out_precision_1_sva_st_113!=2'b01));
  assign mux_860_nl = MUX_s_1_2_2((nor_1623_nl), nor_1664_cse, or_309_cse);
  assign and_242_nl = main_stage_v_2 & (cfg_mode_eql_1_sva_5 | (~(cvt_unequal_tmp_20
      | (mux_860_nl))));
  assign nand_10_nl = ~(cvt_14_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2
      & (~ mux_813_cse));
  assign mux_862_nl = MUX_s_1_2_2((nand_10_nl), cfg_mode_eql_1_sva_6, cvt_unequal_tmp_21);
  assign and_243_nl = main_stage_v_3 & (mux_862_nl);
  assign mux_863_nl = MUX_s_1_2_2((and_243_nl), (and_242_nl), or_5189_cse);
  assign nor_1620_nl = ~((~ cvt_6_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1) | (cfg_proc_precision_1_sva_st_65!=2'b10)
      | (cfg_out_precision_1_sva_st_113!=2'b01));
  assign mux_864_nl = MUX_s_1_2_2((nor_1620_nl), nor_1664_cse, or_309_cse);
  assign and_244_nl = main_stage_v_2 & (cfg_mode_eql_1_sva_5 | (~(cvt_unequal_tmp_20
      | (mux_864_nl))));
  assign nand_11_nl = ~(cvt_6_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2
      & (~ mux_813_cse));
  assign mux_866_nl = MUX_s_1_2_2((nand_11_nl), cfg_mode_eql_1_sva_6, cvt_unequal_tmp_21);
  assign and_245_nl = main_stage_v_3 & (mux_866_nl);
  assign mux_867_nl = MUX_s_1_2_2((and_245_nl), (and_244_nl), or_5189_cse);
  assign nor_1610_nl = ~((~ (chn_idata_data_sva_2_495_479_1[0])) | (cfg_out_precision_1_sva_st_113!=2'b01)
      | (~ main_stage_v_2) | cfg_mode_eql_1_sva_5);
  assign nor_1611_nl = ~((~(cvt_15_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1 | (chn_idata_data_sva_2_495_479_1[0])))
      | (cfg_out_precision_1_sva_st_113!=2'b01) | (~ main_stage_v_2) | cfg_mode_eql_1_sva_5);
  assign mux_868_nl = MUX_s_1_2_2((nor_1611_nl), (nor_1610_nl), or_309_cse);
  assign mux_869_nl = MUX_s_1_2_2((mux_868_nl), nor_1666_cse, cvt_unequal_tmp_20);
  assign nor_1614_nl = ~((~ (chn_idata_data_sva_2_495_479_1[0])) | (~ main_stage_v_2)
      | cfg_mode_eql_1_sva_5);
  assign mux_870_nl = MUX_s_1_2_2((nor_1614_nl), nor_1669_cse, cvt_unequal_tmp_20);
  assign mux_871_nl = MUX_s_1_2_2((mux_870_nl), (mux_869_nl), nor_50_cse);
  assign nand_205_nl = ~((cvt_15_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2
      | (chn_idata_data_sva_3_495_479_1[0])) & or_1159_cse);
  assign mux_872_nl = MUX_s_1_2_2((nand_205_nl), or_1159_cse, cvt_unequal_tmp_21);
  assign or_4528_nl = (~(cvt_15_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2
      | (chn_idata_data_sva_3_495_479_1[0]))) | or_1159_cse;
  assign mux_873_nl = MUX_s_1_2_2((or_4528_nl), nor_1672_cse, cvt_unequal_tmp_21);
  assign mux_874_nl = MUX_s_1_2_2((mux_873_nl), (mux_872_nl), or_1157_cse);
  assign nor_1615_nl = ~((~ main_stage_v_3) | cfg_mode_eql_1_sva_6 | (mux_874_nl));
  assign mux_875_nl = MUX_s_1_2_2((nor_1615_nl), (mux_871_nl), or_5189_cse);
  assign nor_1608_nl = ~((~ cvt_13_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1) | (cfg_proc_precision_1_sva_st_65!=2'b10)
      | (cfg_out_precision_1_sva_st_113!=2'b01));
  assign mux_876_nl = MUX_s_1_2_2((nor_1608_nl), nor_1664_cse, or_309_cse);
  assign and_247_nl = main_stage_v_2 & (cfg_mode_eql_1_sva_5 | (~(cvt_unequal_tmp_20
      | (mux_876_nl))));
  assign nand_13_nl = ~(cvt_13_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2
      & (~ mux_813_cse));
  assign mux_878_nl = MUX_s_1_2_2((nand_13_nl), cfg_mode_eql_1_sva_6, cvt_unequal_tmp_21);
  assign and_248_nl = main_stage_v_3 & (mux_878_nl);
  assign mux_879_nl = MUX_s_1_2_2((and_248_nl), (and_247_nl), or_5189_cse);
  assign nor_1598_nl = ~((~ (chn_idata_data_sva_2_239_223_1[0])) | (cfg_out_precision_1_sva_st_113!=2'b01)
      | (~ main_stage_v_2) | cfg_mode_eql_1_sva_5);
  assign nor_1599_nl = ~((~(cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1 | (chn_idata_data_sva_2_239_223_1[0])))
      | (cfg_out_precision_1_sva_st_113!=2'b01) | (~ main_stage_v_2) | cfg_mode_eql_1_sva_5);
  assign mux_880_nl = MUX_s_1_2_2((nor_1599_nl), (nor_1598_nl), or_309_cse);
  assign mux_881_nl = MUX_s_1_2_2((mux_880_nl), nor_1666_cse, cvt_unequal_tmp_20);
  assign nor_1602_nl = ~((~ (chn_idata_data_sva_2_239_223_1[0])) | (~ main_stage_v_2)
      | cfg_mode_eql_1_sva_5);
  assign mux_882_nl = MUX_s_1_2_2((nor_1602_nl), nor_1669_cse, cvt_unequal_tmp_20);
  assign mux_883_nl = MUX_s_1_2_2((mux_882_nl), (mux_881_nl), nor_50_cse);
  assign nand_204_nl = ~((cvt_7_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2
      | (chn_idata_data_sva_3_239_223_1[0])) & or_1159_cse);
  assign mux_884_nl = MUX_s_1_2_2((nand_204_nl), or_1159_cse, cvt_unequal_tmp_21);
  assign or_4526_nl = (~(cvt_7_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2
      | (chn_idata_data_sva_3_239_223_1[0]))) | or_1159_cse;
  assign mux_885_nl = MUX_s_1_2_2((or_4526_nl), nor_1672_cse, cvt_unequal_tmp_21);
  assign mux_886_nl = MUX_s_1_2_2((mux_885_nl), (mux_884_nl), or_1157_cse);
  assign nor_1603_nl = ~((~ main_stage_v_3) | cfg_mode_eql_1_sva_6 | (mux_886_nl));
  assign mux_887_nl = MUX_s_1_2_2((nor_1603_nl), (mux_883_nl), or_5189_cse);
  assign nor_1596_nl = ~((~ cvt_7_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1) | (cfg_proc_precision_1_sva_st_65!=2'b10)
      | (cfg_out_precision_1_sva_st_113!=2'b01));
  assign mux_888_nl = MUX_s_1_2_2((nor_1596_nl), nor_1664_cse, or_309_cse);
  assign and_250_nl = main_stage_v_2 & (cfg_mode_eql_1_sva_5 | (~(cvt_unequal_tmp_20
      | (mux_888_nl))));
  assign nand_15_nl = ~(cvt_7_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2
      & (~ mux_813_cse));
  assign mux_890_nl = MUX_s_1_2_2((nand_15_nl), cfg_mode_eql_1_sva_6, cvt_unequal_tmp_21);
  assign and_251_nl = main_stage_v_3 & (mux_890_nl);
  assign mux_891_nl = MUX_s_1_2_2((and_251_nl), (and_250_nl), or_5189_cse);
  assign nand_16_nl = ~(nor_63_cse & nor_1048_cse);
  assign nand_17_nl = ~((~(cvt_6_FpMantRNE_17U_11U_else_and_2_svs | (~ FpIntToFloat_17U_5U_10U_else_unequal_tmp_5)
      | (cfg_out_precision_1_sva_st_149!=2'b10))) & nor_1048_cse);
  assign or_1374_nl = (~(cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4
      | (~ cvt_6_FpMantRNE_17U_11U_else_and_2_tmp))) | (~((~((~((libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_21!=5'b00000)))
      | (cfg_out_precision_1_sva_st_149!=2'b10))) & nor_1048_cse));
  assign mux_892_nl = MUX_s_1_2_2((or_1374_nl), (nand_17_nl), FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_3);
  assign and_2190_nl = cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2
      & cvt_unequal_tmp_20;
  assign mux_894_nl = MUX_s_1_2_2((mux_892_nl), (nand_16_nl), and_2190_nl);
  assign mux_895_nl = MUX_s_1_2_2((mux_894_nl), or_1196_cse, nor_50_cse);
  assign or_1375_nl = (~ main_stage_v_2) | cfg_mode_eql_1_sva_5 | (mux_895_nl);
  assign or_1379_nl = (cfg_out_precision_1_sva_st_156!=2'b10) | FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_7
      | nor_183_cse | nor_213_cse | (cfg_out_precision_1_sva_6!=2'b10) | or_tmp_1375;
  assign or_1383_nl = (~ main_stage_v_3) | cfg_mode_eql_1_sva_6;
  assign mux_897_nl = MUX_s_1_2_2((or_1383_nl), or_tmp_1375, or_1157_cse);
  assign mux_898_nl = MUX_s_1_2_2((mux_897_nl), (or_1379_nl), cvt_unequal_tmp_21);
  assign mux_899_nl = MUX_s_1_2_2((mux_898_nl), (or_1375_nl), or_5189_cse);
  assign nor_1584_nl = ~(cvt_unequal_tmp_20 | (cfg_out_precision_1_sva_st_113!=2'b01));
  assign or_1393_nl = (~((~ cvt_15_FpMantRNE_17U_11U_else_and_3_svs) | cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2))
      | (cfg_out_precision_1_sva_st_113!=2'b10) | (~ mux_tmp_416);
  assign mux_902_nl = MUX_s_1_2_2(or_tmp_1393, (or_1393_nl), FpIntToFloat_17U_5U_10U_else_unequal_tmp_14);
  assign or_1399_nl = (~((libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_30!=5'b00000)
      | cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2)) |
      (cfg_out_precision_1_sva_st_113!=2'b10) | (~ mux_tmp_416);
  assign or_1396_nl = (~ cvt_15_FpMantRNE_17U_11U_else_and_3_tmp) | cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4;
  assign mux_903_nl = MUX_s_1_2_2(or_tmp_1393, (or_1399_nl), or_1396_nl);
  assign mux_904_nl = MUX_s_1_2_2((mux_903_nl), (mux_902_nl), FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_3);
  assign nor_1585_nl = ~((cfg_out_precision_1_sva_st_149!=2'b10) | (mux_904_nl));
  assign mux_906_nl = MUX_s_1_2_2((nor_1585_nl), (nor_1584_nl), nor_50_cse);
  assign and_2189_nl = nor_1666_cse & (mux_906_nl);
  assign or_1402_nl = cvt_unequal_tmp_21 | (cfg_out_precision_1_sva_6!=2'b01);
  assign or_1409_nl = (cfg_out_precision_1_sva_st_156!=2'b10) | FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_8
      | nor_183_cse | nor_213_cse | nor_1589_cse | (cfg_out_precision_1_sva_6!=2'b10);
  assign mux_908_nl = MUX_s_1_2_2((or_1409_nl), (or_1402_nl), nor_1672_cse);
  assign nor_1588_nl = ~((~ main_stage_v_3) | cfg_mode_eql_1_sva_6 | (mux_908_nl));
  assign mux_909_nl = MUX_s_1_2_2((nor_1588_nl), (and_2189_nl), or_5189_cse);
  assign mux_2237_nl = MUX_s_1_2_2(and_2422_cse, mux_2230_cse, nor_50_cse);
  assign or_4793_nl = cvt_unequal_tmp_20 | (~ or_4788_cse);
  assign mux_2239_nl = MUX_s_1_2_2(and_2422_cse, (or_4793_nl), cfg_out_precision_1_sva_st_113[1]);
  assign nor_1583_nl = ~((~ cvt_12_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1) | (cfg_proc_precision_1_sva_st_65!=2'b10)
      | (cfg_out_precision_1_sva_st_113!=2'b01));
  assign mux_910_nl = MUX_s_1_2_2((nor_1583_nl), nor_1664_cse, or_309_cse);
  assign and_252_nl = main_stage_v_2 & (cfg_mode_eql_1_sva_5 | (~(cvt_unequal_tmp_20
      | (mux_910_nl))));
  assign nand_21_nl = ~(cvt_12_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2
      & (~ mux_813_cse));
  assign mux_912_nl = MUX_s_1_2_2((nand_21_nl), cfg_mode_eql_1_sva_6, cvt_unequal_tmp_21);
  assign and_253_nl = main_stage_v_3 & (mux_912_nl);
  assign mux_913_nl = MUX_s_1_2_2((and_253_nl), (and_252_nl), or_5189_cse);
  assign nor_1574_nl = ~((~ (chn_idata_data_sva_2_271_255_1[0])) | (cfg_out_precision_1_sva_st_113!=2'b01)
      | (~ main_stage_v_2) | cfg_mode_eql_1_sva_5);
  assign nor_1575_nl = ~((~(cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1 | (chn_idata_data_sva_2_271_255_1[0])))
      | (cfg_out_precision_1_sva_st_113!=2'b01) | (~ main_stage_v_2) | cfg_mode_eql_1_sva_5);
  assign mux_914_nl = MUX_s_1_2_2((nor_1575_nl), (nor_1574_nl), or_309_cse);
  assign mux_915_nl = MUX_s_1_2_2((mux_914_nl), nor_1666_cse, cvt_unequal_tmp_20);
  assign nor_1577_nl = ~((cfg_out_precision_1_sva_st_113!=2'b00) | (~ main_stage_v_2)
      | cfg_mode_eql_1_sva_5);
  assign nor_1578_nl = ~((~ (chn_idata_data_sva_2_271_255_1[0])) | (~ main_stage_v_2)
      | cfg_mode_eql_1_sva_5);
  assign mux_916_nl = MUX_s_1_2_2((nor_1578_nl), (nor_1577_nl), cvt_unequal_tmp_20);
  assign mux_917_nl = MUX_s_1_2_2((mux_916_nl), (mux_915_nl), nor_50_cse);
  assign or_1431_nl = (cfg_out_precision_1_sva_6!=2'b00);
  assign mux_918_nl = MUX_s_1_2_2(nor_1672_cse, or_1159_cse, or_1431_nl);
  assign mux_919_nl = MUX_s_1_2_2(or_1159_cse, (~ or_1159_cse), nor_1629_cse);
  assign nand_22_nl = ~((cvt_8_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2
      | (chn_idata_data_sva_3_271_255_1[0])) & (mux_919_nl));
  assign mux_920_nl = MUX_s_1_2_2((nand_22_nl), (mux_918_nl), cvt_unequal_tmp_21);
  assign nor_1579_nl = ~((~ main_stage_v_3) | cfg_mode_eql_1_sva_6 | (mux_920_nl));
  assign mux_921_nl = MUX_s_1_2_2((nor_1579_nl), (mux_917_nl), or_5189_cse);
  assign nor_1572_nl = ~((~ cvt_8_FpFloatToInt_16U_5U_10U_if_acc_3_itm_11_1) | (cfg_proc_precision_1_sva_st_65!=2'b10)
      | (cfg_out_precision_1_sva_st_113!=2'b01));
  assign mux_922_nl = MUX_s_1_2_2((nor_1572_nl), nor_1664_cse, or_309_cse);
  assign and_255_nl = main_stage_v_2 & (cfg_mode_eql_1_sva_5 | (~(cvt_unequal_tmp_20
      | (mux_922_nl))));
  assign nand_23_nl = ~(cvt_8_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_3_svs_2
      & (~ mux_813_cse));
  assign mux_924_nl = MUX_s_1_2_2((nand_23_nl), cfg_mode_eql_1_sva_6, cvt_unequal_tmp_21);
  assign and_256_nl = main_stage_v_3 & (mux_924_nl);
  assign mux_925_nl = MUX_s_1_2_2((and_256_nl), (and_255_nl), or_5189_cse);
  assign nor_1569_nl = ~((~ cvt_11_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1) | (cfg_proc_precision_1_sva_st_65!=2'b10)
      | (cfg_out_precision_1_sva_st_113!=2'b01));
  assign mux_926_nl = MUX_s_1_2_2((nor_1569_nl), nor_1664_cse, or_309_cse);
  assign and_257_nl = main_stage_v_2 & (cfg_mode_eql_1_sva_5 | (~(cvt_unequal_tmp_20
      | (mux_926_nl))));
  assign nand_24_nl = ~(cvt_11_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2
      & (~ mux_813_cse));
  assign mux_928_nl = MUX_s_1_2_2((nand_24_nl), cfg_mode_eql_1_sva_6, cvt_unequal_tmp_21);
  assign and_258_nl = main_stage_v_3 & (mux_928_nl);
  assign mux_929_nl = MUX_s_1_2_2((and_258_nl), (and_257_nl), or_5189_cse);
  assign nor_1566_nl = ~((~ cvt_9_FpFloatToInt_16U_5U_10U_if_acc_1_itm_11_1) | (cfg_proc_precision_1_sva_st_65!=2'b10)
      | (cfg_out_precision_1_sva_st_113!=2'b01));
  assign mux_930_nl = MUX_s_1_2_2((nor_1566_nl), nor_1664_cse, or_309_cse);
  assign and_259_nl = main_stage_v_2 & (cfg_mode_eql_1_sva_5 | (~(cvt_unequal_tmp_20
      | (mux_930_nl))));
  assign nand_25_nl = ~(cvt_9_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_1_svs_2
      & (~ mux_813_cse));
  assign mux_932_nl = MUX_s_1_2_2((nand_25_nl), cfg_mode_eql_1_sva_6, cvt_unequal_tmp_21);
  assign and_260_nl = main_stage_v_3 & (mux_932_nl);
  assign mux_933_nl = MUX_s_1_2_2((and_260_nl), (and_259_nl), or_5189_cse);
  assign nor_1563_nl = ~((~ cvt_10_FpFloatToInt_16U_5U_10U_if_acc_2_itm_11_1) | (cfg_proc_precision_1_sva_st_65!=2'b10)
      | (cfg_out_precision_1_sva_st_113!=2'b01));
  assign mux_934_nl = MUX_s_1_2_2((nor_1563_nl), nor_1664_cse, or_309_cse);
  assign and_261_nl = main_stage_v_2 & (cfg_mode_eql_1_sva_5 | (~(cvt_unequal_tmp_20
      | (mux_934_nl))));
  assign nand_26_nl = ~(cvt_10_FpFloatToInt_16U_5U_10U_if_slc_FpFloatToInt_16U_5U_10U_if_acc_11_2_svs_2
      & (~ mux_813_cse));
  assign mux_936_nl = MUX_s_1_2_2((nand_26_nl), cfg_mode_eql_1_sva_6, cvt_unequal_tmp_21);
  assign and_262_nl = main_stage_v_3 & (mux_936_nl);
  assign mux_937_nl = MUX_s_1_2_2((and_262_nl), (and_261_nl), or_5189_cse);
  assign nl_cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_sva_2
      , IntShiftRightSat_49U_6U_17U_o_15_1_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_sva_2})
      + 18'b111111111111111111;
  assign cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl = nl_cvt_16_IntShiftRightSat_49U_6U_17U_oif_1_acc_4_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_24_nl = MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_lpi_1_dfm,
      IntShiftRightSat_49U_6U_17U_lor_lpi_1_dfm_mx1w0, and_tmp_225);
  assign nl_cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_15_sva_2
      , IntShiftRightSat_49U_6U_17U_o_15_1_15_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_15_sva_2})
      + 18'b111111111111111111;
  assign cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl = nl_cvt_15_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_26_nl = MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_16_lpi_1_dfm_mx1w0,
      IntShiftRightSat_49U_6U_17U_lor_16_lpi_1_dfm, or_3817_cse);
  assign nl_cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_14_sva_2
      , IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_14_sva_3})
      + 18'b111111111111111111;
  assign cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl = nl_cvt_14_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_22_nl = MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_15_lpi_1_dfm_mx1w0,
      IntShiftRightSat_49U_6U_17U_lor_15_lpi_1_dfm, or_3817_cse);
  assign nl_cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_13_sva_2
      , IntShiftRightSat_49U_6U_17U_o_15_1_13_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_13_sva_2})
      + 18'b111111111111111111;
  assign cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl = nl_cvt_13_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_28_nl = MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_14_lpi_1_dfm_mx1w0,
      IntShiftRightSat_49U_6U_17U_lor_14_lpi_1_dfm, or_3817_cse);
  assign nl_cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_12_sva_2
      , IntShiftRightSat_49U_6U_17U_o_15_1_12_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_12_sva_2})
      + 18'b111111111111111111;
  assign cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl = nl_cvt_12_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_18_nl = MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_13_lpi_1_dfm,
      IntShiftRightSat_49U_6U_17U_lor_13_lpi_1_dfm_mx1w0, mux_1142_cse);
  assign nl_cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_11_sva_2
      , IntShiftRightSat_49U_6U_17U_o_15_1_11_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_11_sva_2})
      + 18'b111111111111111111;
  assign cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl = nl_cvt_11_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_20_nl = MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_12_lpi_1_dfm_mx1w0,
      IntShiftRightSat_49U_6U_17U_lor_12_lpi_1_dfm, or_3817_cse);
  assign nl_cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_10_sva_2
      , IntShiftRightSat_49U_6U_17U_o_15_1_10_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_10_sva_2})
      + 18'b111111111111111111;
  assign cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl = nl_cvt_10_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_16_nl = MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_11_lpi_1_dfm_mx1w0,
      IntShiftRightSat_49U_6U_17U_lor_11_lpi_1_dfm, or_3817_cse);
  assign nl_cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_9_sva_3
      , IntShiftRightSat_49U_6U_17U_o_15_1_9_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_9_sva_3})
      + 18'b111111111111111111;
  assign cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl = nl_cvt_9_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_30_nl = MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_10_lpi_1_dfm,
      IntShiftRightSat_49U_6U_17U_lor_10_lpi_1_dfm_mx1w0, mux_tmp_455);
  assign nl_cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_8_sva_2
      , IntShiftRightSat_49U_6U_17U_o_15_1_8_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_8_sva_2})
      + 18'b111111111111111111;
  assign cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl = nl_cvt_8_IntShiftRightSat_49U_6U_17U_oif_1_acc_3_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_10_nl = MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_9_lpi_1_dfm_mx1w0,
      IntShiftRightSat_49U_6U_17U_lor_9_lpi_1_dfm, or_3774_cse);
  assign nl_cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_7_sva_2
      , IntShiftRightSat_49U_6U_17U_o_15_1_7_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_7_sva_2})
      + 18'b111111111111111111;
  assign cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl = nl_cvt_7_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_12_nl = MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_8_lpi_1_dfm_mx1w0,
      IntShiftRightSat_49U_6U_17U_lor_8_lpi_1_dfm, or_3774_cse);
  assign nl_cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_6_sva_2
      , IntShiftRightSat_49U_6U_17U_o_15_1_6_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_6_sva_2})
      + 18'b111111111111111111;
  assign cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl = nl_cvt_6_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_8_nl = MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_7_lpi_1_dfm_mx1w0,
      IntShiftRightSat_49U_6U_17U_lor_7_lpi_1_dfm, or_3774_cse);
  assign nl_cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_5_sva_3
      , IntShiftRightSat_49U_6U_17U_o_15_1_5_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_5_sva_3})
      + 18'b111111111111111111;
  assign cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl = nl_cvt_5_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_14_nl = MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_6_lpi_1_dfm_mx1w0,
      IntShiftRightSat_49U_6U_17U_lor_6_lpi_1_dfm, or_dcpl_163);
  assign nl_cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_4_sva_2
      , IntShiftRightSat_49U_6U_17U_o_15_1_4_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_4_sva_2})
      + 18'b111111111111111111;
  assign cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl = nl_cvt_4_IntShiftRightSat_49U_6U_17U_oif_1_acc_2_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_4_nl = MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_5_lpi_1_dfm_mx1w0,
      IntShiftRightSat_49U_6U_17U_lor_5_lpi_1_dfm, or_dcpl_353);
  assign nl_cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_3_sva_3
      , IntShiftRightSat_49U_6U_17U_o_15_1_3_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_3_sva_3})
      + 18'b111111111111111111;
  assign cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl = nl_cvt_3_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_6_nl = MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_4_lpi_1_dfm,
      IntShiftRightSat_49U_6U_17U_lor_4_lpi_1_dfm_mx1w0, and_tmp_50);
  assign nl_cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_2_sva_2
      , IntShiftRightSat_49U_6U_17U_o_15_1_2_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_2_sva_2})
      + 18'b111111111111111111;
  assign cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl = nl_cvt_2_IntShiftRightSat_49U_6U_17U_oif_1_acc_1_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_2_nl = MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_3_lpi_1_dfm_mx1w0,
      IntShiftRightSat_49U_6U_17U_lor_3_lpi_1_dfm, or_dcpl_151);
  assign nl_cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl = conv_s2s_17_18({IntShiftRightSat_49U_6U_17U_o_16_1_sva_3
      , IntShiftRightSat_49U_6U_17U_o_15_1_1_sva_2 , IntShiftRightSat_49U_6U_17U_o_0_1_sva_2})
      + 18'b111111111111111111;
  assign cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl = nl_cvt_1_IntShiftRightSat_49U_6U_17U_oif_1_acc_nl[17:0];
  assign IntShiftRightSat_49U_6U_17U_oelse_mux_32_nl = MUX_s_1_2_2(IntShiftRightSat_49U_6U_17U_lor_2_lpi_1_dfm,
      IntShiftRightSat_49U_6U_17U_lor_2_lpi_1_dfm_mx1w0, or_4862_cse);
  assign or_1483_nl = (~ main_stage_v_2) | (~ cvt_unequal_tmp_20) | cfg_mode_eql_1_sva_5;
  assign or_1484_nl = cvt_1_IntSaturation_17U_8U_if_acc_itm_10_1 | (~ main_stage_v_2)
      | (~ cvt_unequal_tmp_20) | cfg_mode_eql_1_sva_5;
  assign mux_939_nl = MUX_s_1_2_2((or_1484_nl), (or_1483_nl), cfg_out_precision_1_sva_st_113[1]);
  assign nor_1557_nl = ~((cfg_out_precision_1_sva_st_113[0]) | (mux_939_nl));
  assign mux_940_nl = MUX_s_1_2_2((nor_1557_nl), nor_1556_cse, nor_50_cse);
  assign nor_1558_nl = ~((~ main_stage_v_3) | (~ cvt_unequal_tmp_21) | cfg_mode_eql_1_sva_6
      | (cfg_out_precision_1_sva_6[0]) | (~((~((cfg_out_precision_1_sva_st_136!=2'b00)
      | cvt_1_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_svs_st_2))
      | (cfg_out_precision_1_sva_6[1]))));
  assign mux_943_nl = MUX_s_1_2_2((nor_1558_nl), (mux_940_nl), or_5189_cse);
  assign nl_cvt_14_IntSaturation_17U_8U_if_acc_3_nl = conv_s2u_10_11({(~ IntShiftRightSat_49U_6U_17U_o_16_14_sva_2)
      , (~ (IntShiftRightSat_49U_6U_17U_o_15_1_14_sva_2[14:6]))}) + 11'b1;
  assign cvt_14_IntSaturation_17U_8U_if_acc_3_nl = nl_cvt_14_IntSaturation_17U_8U_if_acc_3_nl[10:0];
  assign mux_949_nl = MUX_s_1_2_2(and_2186_cse, mux_tmp_117, main_stage_v_1);
  assign mux_950_nl = MUX_s_1_2_2((mux_949_nl), mux_tmp_321, main_stage_v_2);
  assign nor_1555_nl = ~((cfg_proc_precision_1_sva_st_90[1]) | (~ and_tmp_166));
  assign mux_951_nl = MUX_s_1_2_2((nor_1555_nl), and_tmp_166, cfg_proc_precision_1_sva_st_90[0]);
  assign mux_952_nl = MUX_s_1_2_2(and_tmp_16, mux_tmp_321, main_stage_v_2);
  assign mux_953_nl = MUX_s_1_2_2((mux_952_nl), (mux_951_nl), main_stage_v_3);
  assign mux_954_nl = MUX_s_1_2_2((mux_953_nl), (mux_950_nl), or_5189_cse);
  assign nor_1547_nl = ~((~ main_stage_v_2) | (~ cvt_unequal_tmp_20) | cfg_mode_eql_1_sva_5
      | (cfg_out_precision_1_sva_st_113[0]) | (~((cfg_out_precision_1_sva_st_113[1])
      | (~((cfg_out_precision_1_sva_st_149!=2'b00) | cvt_3_IntSaturation_17U_8U_if_acc_1_itm_10_1
      | nor_2219_cse)))));
  assign nor_1548_nl = ~((~ main_stage_v_3) | (~ cvt_unequal_tmp_21) | cfg_mode_eql_1_sva_6
      | (cfg_out_precision_1_sva_6[0]) | (~((cfg_out_precision_1_sva_6[1]) | (~((cfg_out_precision_1_sva_st_144!=2'b00)
      | cvt_3_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2
      | nor_213_cse)))));
  assign mux_959_nl = MUX_s_1_2_2((nor_1548_nl), (nor_1547_nl), or_5189_cse);
  assign mux_964_nl = MUX_s_1_2_2(mux_tmp_963, mux_tmp_961, or_5189_cse);
  assign nor_1537_nl = ~((~ main_stage_v_2) | (~ cvt_unequal_tmp_20) | cfg_mode_eql_1_sva_5
      | (cfg_out_precision_1_sva_st_113[0]) | (~((cfg_out_precision_1_sva_st_113[1])
      | (~((cfg_out_precision_1_sva_st_149!=2'b00) | cvt_5_IntSaturation_17U_8U_if_acc_1_itm_10_1
      | nor_2219_cse)))));
  assign nor_1538_nl = ~((~ main_stage_v_3) | (~ cvt_unequal_tmp_21) | cfg_mode_eql_1_sva_6
      | (cfg_out_precision_1_sva_6[0]) | (~((cfg_out_precision_1_sva_6[1]) | (~((cfg_out_precision_1_sva_st_144!=2'b00)
      | cvt_5_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2
      | nor_213_cse)))));
  assign mux_982_nl = MUX_s_1_2_2((nor_1538_nl), (nor_1537_nl), or_5189_cse);
  assign mux_995_nl = MUX_s_1_2_2(mux_tmp_994, mux_tmp_992, or_5189_cse);
  assign nor_1526_nl = ~((~ main_stage_v_2) | (~ cvt_unequal_tmp_20) | cfg_mode_eql_1_sva_5
      | (cfg_out_precision_1_sva_st_113[0]) | (~((cfg_out_precision_1_sva_st_113[1])
      | (~((cfg_out_precision_1_sva_st_149!=2'b00) | cvt_9_IntSaturation_17U_8U_if_acc_1_itm_10_1
      | nor_2219_cse)))));
  assign nor_1527_nl = ~((~ main_stage_v_3) | (~ cvt_unequal_tmp_21) | cfg_mode_eql_1_sva_6
      | (cfg_out_precision_1_sva_6[0]) | (~((cfg_out_precision_1_sva_6[1]) | (~((cfg_out_precision_1_sva_st_144!=2'b00)
      | cvt_9_IntSaturation_17U_8U_if_slc_IntSaturation_17U_8U_if_acc_10_1_svs_st_2
      | nor_213_cse)))));
  assign mux_1000_nl = MUX_s_1_2_2((nor_1527_nl), (nor_1526_nl), or_5189_cse);
  assign or_3841_nl = and_dcpl_942 | cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_svs_st_2;
  assign FpMantRNE_17U_11U_else_mux_1_nl = MUX_s_1_2_2(cvt_1_FpMantRNE_17U_11U_else_and_tmp,
      cvt_1_FpMantRNE_17U_11U_else_and_svs, or_3841_nl);
  assign FpIntToFloat_17U_5U_10U_else_mux_1_nl = MUX_s_1_2_2(or_1202_cse, FpIntToFloat_17U_5U_10U_else_unequal_tmp,
      cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_svs_st_2);
  assign nor_1519_nl = ~((~ main_stage_v_2) | (cfg_out_precision_1_sva_st_113!=2'b10)
      | (~ cvt_unequal_tmp_20) | cfg_mode_eql_1_sva_5 | nor_50_cse);
  assign nor_1521_nl = ~(nor_1672_cse | (~ main_stage_v_3) | (~ cvt_unequal_tmp_21)
      | cfg_mode_eql_1_sva_6 | (cfg_out_precision_1_sva_6!=2'b10) | (cfg_out_precision_1_sva_st_136!=2'b10));
  assign mux_1004_nl = MUX_s_1_2_2((nor_1521_nl), (nor_1519_nl), or_5189_cse);
  assign and_2811_nl = (~((FpIntToFloat_17U_5U_10U_else_int_mant_1_sva[16:5]==12'b111111111111)))
      & or_1202_cse;
  assign mux_2250_nl = MUX_s_1_2_2((and_2811_nl), or_1202_cse, cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_1_itm_4);
  assign nor_2461_nl = ~(((~ cvt_1_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_1_itm_4)
      & (FpIntToFloat_17U_5U_10U_else_int_mant_1_sva[16:5]==12'b111111111111)) |
      (cfg_out_precision_1_sva_st_113!=2'b10) | cvt_1_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_svs_st_2
      | IsNaN_5U_10U_IsNaN_5U_10U_nand_1_itm_2 | (~((libraries_leading_sign_17_0_6b58f91630d78ab00051ea7ca02e26cb4a6f_16!=5'b00000))));
  assign mux_2251_nl = MUX_s_1_2_2((nor_2461_nl), nor_2099_cse, nor_50_cse);
  assign nor_1510_nl = ~((~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt
      | (~ main_stage_v_3) | (cfg_out_precision_1_sva_st_136!=2'b00) | (~ or_1159_cse));
  assign nor_1511_nl = ~((~ main_stage_v_3) | (cfg_out_precision_1_sva_st_136!=2'b00)
      | (~ or_1159_cse));
  assign mux_1010_nl = MUX_s_1_2_2((nor_1511_nl), and_2237_cse, or_5189_cse);
  assign mux_1011_nl = MUX_s_1_2_2((mux_1010_nl), (nor_1510_nl), or_425_cse);
  assign or_3850_nl = and_dcpl_946 | cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign FpMantRNE_17U_11U_else_mux_3_nl = MUX_s_1_2_2(cvt_2_FpMantRNE_17U_11U_else_and_1_tmp,
      cvt_2_FpMantRNE_17U_11U_else_and_1_svs, or_3850_nl);
  assign FpIntToFloat_17U_5U_10U_else_mux_4_nl = MUX_s_1_2_2(or_1596_cse, FpIntToFloat_17U_5U_10U_else_unequal_tmp_1,
      cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2);
  assign FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_nor_1_nl
      = ~(((~((~ cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4) & (FpMantRNE_17U_11U_else_mux_3_nl)))
      & (FpIntToFloat_17U_5U_10U_else_mux_4_nl)) | cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2);
  assign nor_1508_nl = ~(main_stage_v_2 | (~ mux_tmp_944));
  assign mux_1012_nl = MUX_s_1_2_2((nor_1508_nl), mux_tmp_945, or_1587_cse);
  assign mux_1016_nl = MUX_s_1_2_2(mux_tmp_1015, (mux_1012_nl), or_5189_cse);
  assign mux_1017_nl = MUX_s_1_2_2(mux_tmp_1015, mux_tmp_945, or_5189_cse);
  assign mux_1018_nl = MUX_s_1_2_2((mux_1017_nl), (mux_1016_nl), nor_63_cse);
  assign and_2809_nl = (~((FpIntToFloat_17U_5U_10U_else_int_mant_2_sva[16:5]==12'b111111111111)))
      & or_1596_cse;
  assign mux_2252_nl = MUX_s_1_2_2((and_2809_nl), or_1596_cse, cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4);
  assign nor_2457_nl = ~((cfg_out_precision_1_sva_st_149!=2'b10) | cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2
      | cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 | nor_2219_cse
      | (~(or_1596_cse & (~(((~ cvt_2_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4)
      & (FpIntToFloat_17U_5U_10U_else_int_mant_2_sva[16:5]==12'b111111111111)) |
      (cfg_out_precision_1_sva_st_113!=2'b10))))));
  assign mux_2253_nl = MUX_s_1_2_2((nor_2457_nl), nor_2099_cse, nor_50_cse);
  assign or_3860_nl = and_dcpl_950 | cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign FpMantRNE_17U_11U_else_mux_5_nl = MUX_s_1_2_2(cvt_3_FpMantRNE_17U_11U_else_and_1_tmp,
      cvt_3_FpMantRNE_17U_11U_else_and_1_svs, or_3860_nl);
  assign FpIntToFloat_17U_5U_10U_else_mux_7_nl = MUX_s_1_2_2(or_1625_cse, FpIntToFloat_17U_5U_10U_else_unequal_tmp_2,
      cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2);
  assign or_3879_nl = and_dcpl_958 | cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign FpMantRNE_17U_11U_else_mux_9_nl = MUX_s_1_2_2(cvt_5_FpMantRNE_17U_11U_else_and_1_tmp,
      cvt_5_FpMantRNE_17U_11U_else_and_1_svs, or_3879_nl);
  assign FpIntToFloat_17U_5U_10U_else_mux_13_nl = MUX_s_1_2_2(or_1693_cse, FpIntToFloat_17U_5U_10U_else_unequal_tmp_4,
      cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2);
  assign and_2807_nl = (~((cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[16:5]==12'b111111111111)))
      & or_1625_cse;
  assign mux_2254_nl = MUX_s_1_2_2((and_2807_nl), or_1625_cse, cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4);
  assign nor_2453_nl = ~((cfg_out_precision_1_sva_st_149!=2'b10) | cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2
      | cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 | nor_2219_cse
      | (~(or_1625_cse & (~(((~ cvt_3_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4)
      & (cvt_3_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[16:5]==12'b111111111111))
      | (cfg_out_precision_1_sva_st_113!=2'b10))))));
  assign mux_2255_nl = MUX_s_1_2_2((nor_2453_nl), nor_2099_cse, nor_50_cse);
  assign mux_1034_nl = MUX_s_1_2_2(nor_1489_cse, and_1078_cse, or_5189_cse);
  assign mux_1035_nl = MUX_s_1_2_2((mux_1034_nl), nor_1488_cse, or_461_cse);
  assign mux_1044_nl = MUX_s_1_2_2(mux_tmp_1043, (~ or_tmp_1650), cfg_proc_precision_1_sva_st_101[1]);
  assign mux_1045_nl = MUX_s_1_2_2((mux_1044_nl), mux_tmp_1043, cfg_proc_precision_1_sva_st_101[0]);
  assign mux_1054_nl = MUX_s_1_2_2(mux_1053_cse, (mux_1045_nl), main_stage_v_2);
  assign and_2805_nl = (~((cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:5]==12'b111111111111)))
      & or_1659_cse_1;
  assign mux_2256_nl = MUX_s_1_2_2((and_2805_nl), or_1659_cse_1, cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4);
  assign nor_2449_nl = ~((cfg_out_precision_1_sva_st_149!=2'b10) | FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_3
      | cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 | nor_2219_cse
      | nor_151_cse | (~(or_1659_cse_1 & (~(((~ cvt_4_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4)
      & (cvt_4_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:5]==12'b111111111111))
      | (cfg_out_precision_1_sva_st_113!=2'b10))))));
  assign mux_2257_nl = MUX_s_1_2_2((nor_2449_nl), nor_2099_cse, nor_50_cse);
  assign and_2803_nl = (~((cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[16:5]==12'b111111111111)))
      & or_1693_cse;
  assign mux_2258_nl = MUX_s_1_2_2((and_2803_nl), or_1693_cse, cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4);
  assign nor_2445_nl = ~((cfg_out_precision_1_sva_st_149!=2'b10) | cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2
      | cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2 | nor_2219_cse
      | (~(or_1693_cse & (~(((~ cvt_5_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4)
      & (cvt_5_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_1_tmp[16:5]==12'b111111111111))
      | (cfg_out_precision_1_sva_st_113!=2'b10))))));
  assign mux_2259_nl = MUX_s_1_2_2((nor_2445_nl), nor_2099_cse, nor_50_cse);
  assign nor_1465_nl = ~((~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt
      | (~ main_stage_v_3) | (cfg_out_precision_1_sva_st_144!=2'b00) | (~ and_tmp_165));
  assign nor_1466_nl = ~((~ main_stage_v_3) | (cfg_out_precision_1_sva_st_144!=2'b00)
      | (~ and_tmp_165));
  assign mux_1069_nl = MUX_s_1_2_2((nor_1466_nl), and_2230_cse, or_5189_cse);
  assign mux_1070_nl = MUX_s_1_2_2((mux_1069_nl), (nor_1465_nl), or_461_cse);
  assign mux_1075_nl = MUX_s_1_2_2(mux_tmp_1074, mux_1071_cse, or_5189_cse);
  assign mux_1076_nl = MUX_s_1_2_2(mux_tmp_1074, mux_tmp_961, or_5189_cse);
  assign mux_1077_nl = MUX_s_1_2_2((mux_1076_nl), (mux_1075_nl), nor_63_cse);
  assign and_2801_nl = (~((cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:5]==12'b111111111111)))
      & or_1720_cse_1;
  assign mux_2260_nl = MUX_s_1_2_2((and_2801_nl), or_1720_cse_1, cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4);
  assign nor_2441_nl = ~((cfg_out_precision_1_sva_st_149!=2'b10) | FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_3
      | cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 | nor_2219_cse
      | nor_151_cse | (~(or_1720_cse_1 & (~(((~ cvt_6_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4)
      & (cvt_6_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:5]==12'b111111111111))
      | (cfg_out_precision_1_sva_st_113!=2'b10))))));
  assign mux_2261_nl = MUX_s_1_2_2((nor_2441_nl), nor_2099_cse, nor_50_cse);
  assign mux_1089_nl = MUX_s_1_2_2(mux_tmp_1088, mux_1071_cse, or_5189_cse);
  assign mux_1090_nl = MUX_s_1_2_2(mux_tmp_1088, mux_tmp_961, or_5189_cse);
  assign mux_1091_nl = MUX_s_1_2_2((mux_1090_nl), (mux_1089_nl), nor_63_cse);
  assign and_2799_nl = (~((cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:5]==12'b111111111111)))
      & or_1752_cse_1;
  assign mux_2262_nl = MUX_s_1_2_2((and_2799_nl), or_1752_cse_1, cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4);
  assign nor_2437_nl = ~((cfg_out_precision_1_sva_st_149!=2'b10) | FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_3
      | cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2 | nor_2219_cse
      | nor_151_cse | (~(or_1752_cse_1 & (~(((~ cvt_7_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4)
      & (cvt_7_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:5]==12'b111111111111))
      | (cfg_out_precision_1_sva_st_113!=2'b10))))));
  assign mux_2263_nl = MUX_s_1_2_2((nor_2437_nl), nor_2099_cse, nor_50_cse);
  assign mux_1106_nl = MUX_s_1_2_2(mux_tmp_1105, (~ or_tmp_1780), cfg_proc_precision_1_sva_st_101[1]);
  assign mux_1107_nl = MUX_s_1_2_2((mux_1106_nl), mux_tmp_1105, cfg_proc_precision_1_sva_st_101[0]);
  assign mux_1112_nl = MUX_s_1_2_2(mux_tmp_1111, (~ or_tmp_1780), cfg_proc_precision_1_sva_st_64[1]);
  assign mux_1113_nl = MUX_s_1_2_2((mux_1112_nl), mux_tmp_1111, cfg_proc_precision_1_sva_st_64[0]);
  assign mux_1114_nl = MUX_s_1_2_2(and_tmp_175, and_2186_cse, or_5189_cse);
  assign mux_1115_nl = MUX_s_1_2_2((mux_1114_nl), (mux_1113_nl), main_stage_v_1);
  assign mux_1116_nl = MUX_s_1_2_2((mux_1115_nl), (mux_1107_nl), main_stage_v_2);
  assign and_2797_nl = (~((cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[16:5]==12'b111111111111)))
      & or_1789_cse_1;
  assign mux_2264_nl = MUX_s_1_2_2((and_2797_nl), or_1789_cse_1, cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4);
  assign nor_2433_nl = ~((cfg_out_precision_1_sva_st_149!=2'b10) | FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_3
      | cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2 | nor_2219_cse
      | nor_151_cse | (~(or_1789_cse_1 & (~(((~ cvt_8_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4)
      & (cvt_8_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[16:5]==12'b111111111111))
      | (cfg_out_precision_1_sva_st_113!=2'b10))))));
  assign mux_2265_nl = MUX_s_1_2_2((nor_2433_nl), nor_2099_cse, nor_50_cse);
  assign or_3920_nl = and_dcpl_974 | cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2;
  assign FpMantRNE_17U_11U_else_mux_17_nl = MUX_s_1_2_2(cvt_9_FpMantRNE_17U_11U_else_and_1_tmp,
      cvt_9_FpMantRNE_17U_11U_else_and_1_svs, or_3920_nl);
  assign FpIntToFloat_17U_5U_10U_else_mux_25_nl = MUX_s_1_2_2(or_1829_cse, FpIntToFloat_17U_5U_10U_else_unequal_tmp_8,
      cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2);
  assign nor_1433_nl = ~((~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | (~ cvt_unequal_tmp_20) | cfg_mode_eql_1_sva_5 | (cfg_out_precision_1_sva_st_113!=2'b10)
      | (~ mux_1126_cse));
  assign mux_1127_nl = MUX_s_1_2_2(nor_1500_cse, (nor_1433_nl), or_5189_cse);
  assign and_2795_nl = (~((FpIntToFloat_17U_5U_10U_else_int_mant_9_sva[16:5]==12'b111111111111)))
      & or_1829_cse;
  assign mux_2266_nl = MUX_s_1_2_2((and_2795_nl), or_1829_cse, cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4);
  assign nor_2429_nl = ~(nor_2219_cse | (cfg_out_precision_1_sva_st_149!=2'b10) |
      cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 | cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_2
      | (~(or_1829_cse & (~(((~ cvt_9_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_2_itm_4)
      & (FpIntToFloat_17U_5U_10U_else_int_mant_9_sva[16:5]==12'b111111111111)) |
      (cfg_out_precision_1_sva_st_113!=2'b10))))));
  assign mux_2267_nl = MUX_s_1_2_2((nor_2429_nl), nor_2099_cse, nor_50_cse);
  assign mux_1133_nl = MUX_s_1_2_2(nor_1489_cse, and_tmp_94, or_5189_cse);
  assign mux_1134_nl = MUX_s_1_2_2((mux_1133_nl), nor_1488_cse, or_461_cse);
  assign and_2793_nl = (~((cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:5]==12'b111111111111)))
      & or_1851_cse_1;
  assign mux_2268_nl = MUX_s_1_2_2((and_2793_nl), or_1851_cse_1, cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4);
  assign nor_2425_nl = ~(nor_2219_cse | (cfg_out_precision_1_sva_st_149!=2'b10) |
      FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_3 | cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2
      | (~(or_400_cse_1 & or_1851_cse_1 & (~(((~ cvt_10_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4)
      & (cvt_10_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:5]==12'b111111111111))
      | (cfg_out_precision_1_sva_st_113!=2'b10))))));
  assign mux_2269_nl = MUX_s_1_2_2((nor_2425_nl), nor_2099_cse, nor_50_cse);
  assign mux_1153_nl = MUX_s_1_2_2(mux_tmp_1152, (~ or_tmp_1650), cfg_proc_precision_1_sva_st_89[1]);
  assign mux_1154_nl = MUX_s_1_2_2((mux_1153_nl), mux_tmp_1152, cfg_proc_precision_1_sva_st_89[0]);
  assign mux_1163_nl = MUX_s_1_2_2(mux_1053_cse, (mux_1154_nl), main_stage_v_2);
  assign and_2791_nl = (~((cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:5]==12'b111111111111)))
      & or_1892_cse_1;
  assign mux_2270_nl = MUX_s_1_2_2((and_2791_nl), or_1892_cse_1, cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4);
  assign and_2789_nl = or_400_cse_1 & (~(nor_2219_cse | (cfg_out_precision_1_sva_st_149!=2'b10)
      | FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_3 | cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2
      | (~(or_1892_cse_1 & (~(((~ cvt_11_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4)
      & (cvt_11_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:5]==12'b111111111111))
      | (cfg_out_precision_1_sva_st_113!=2'b10)))))));
  assign mux_2271_nl = MUX_s_1_2_2((and_2789_nl), nor_2099_cse, nor_50_cse);
  assign and_3372_nl = mux_1142_cse & (~ (cfg_out_precision_1_sva_st_149[1]));
  assign mux_1172_nl = MUX_s_1_2_2((and_3372_nl), mux_1142_cse, cfg_out_precision_1_sva_st_149[0]);
  assign mux_1173_nl = MUX_s_1_2_2(mux_tmp_944, (mux_1172_nl), main_stage_v_2);
  assign mux_1174_nl = MUX_s_1_2_2((mux_1173_nl), mux_tmp_992, or_1587_cse);
  assign nor_1403_nl = ~((cfg_proc_precision_1_sva_st_108[0]) | (~((cfg_proc_precision_1_sva_st_108[1])
      & mux_tmp_987)));
  assign mux_1175_nl = MUX_s_1_2_2(mux_tmp_987, (nor_1403_nl), cfg_out_precision_1_sva_6[1]);
  assign mux_1176_nl = MUX_s_1_2_2((mux_1175_nl), mux_tmp_987, or_1919_cse);
  assign mux_1177_nl = MUX_s_1_2_2(mux_989_cse, (mux_1176_nl), main_stage_v_3);
  assign or_1918_nl = (~ cvt_unequal_tmp_21) | (cfg_out_precision_1_sva_st_156!=2'b10);
  assign mux_1178_nl = MUX_s_1_2_2((mux_1177_nl), mux_tmp_994, or_1918_nl);
  assign mux_1179_nl = MUX_s_1_2_2((mux_1178_nl), (mux_1174_nl), or_5189_cse);
  assign and_2788_nl = (~((cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[16:5]==12'b111111111111)))
      & or_1925_cse_1;
  assign mux_2272_nl = MUX_s_1_2_2((and_2788_nl), or_1925_cse_1, cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4);
  assign and_3373_nl = or_400_cse_1 & (~(nor_2219_cse | (cfg_out_precision_1_sva_st_149!=2'b10)
      | FpIntToFloat_17U_5U_10U_is_inf_12_lpi_1_dfm_3 | cvt_12_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2
      | (~(or_1925_cse_1 & (~(((~ cvt_12_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4)
      & (cvt_12_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[16:5]==12'b111111111111))
      | (cfg_out_precision_1_sva_st_113!=2'b10)))))));
  assign mux_2273_nl = MUX_s_1_2_2((and_3373_nl), nor_2099_cse, nor_50_cse);
  assign and_2786_nl = (~((cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:5]==12'b111111111111)))
      & or_5038_cse;
  assign mux_2274_nl = MUX_s_1_2_2((and_2786_nl), or_5038_cse, cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4);
  assign nor_2411_nl = ~(((~ cvt_13_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_4_tmp_4)
      & (cvt_13_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_2_tmp[16:5]==12'b111111111111))
      | (~(or_5038_cse & or_400_cse_1 & (~(nor_2219_cse | (cfg_out_precision_1_sva_st_149!=2'b10)
      | FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_3 | cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_svs_2
      | (cfg_out_precision_1_sva_st_113!=2'b10))))));
  assign mux_2275_nl = MUX_s_1_2_2((nor_2411_nl), nor_2099_cse, nor_50_cse);
  assign nand_45_nl = ~(main_stage_v_2 & (~(nor_50_cse | nor_2219_cse | nor_151_cse
      | or_425_cse)));
  assign nand_201_nl = ~(cvt_else_equal_tmp_46 & main_stage_v_3 & mux_tmp_1197);
  assign mux_1202_nl = MUX_s_1_2_2(or_tmp_1981, (nand_201_nl), cfg_proc_precision_1_sva_st_108[1]);
  assign mux_1203_nl = MUX_s_1_2_2((mux_1202_nl), or_tmp_1981, cfg_proc_precision_1_sva_st_108[0]);
  assign mux_1204_nl = MUX_s_1_2_2((mux_1203_nl), (nand_45_nl), or_5189_cse);
  assign nand_46_nl = ~(main_stage_v_2 & (~(nor_50_cse | nor_2219_cse | nor_151_cse
      | or_300_cse)));
  assign nand_199_nl = ~(cvt_else_equal_tmp_45 & main_stage_v_3 & mux_tmp_1197);
  assign mux_1211_nl = MUX_s_1_2_2(or_tmp_1992, (nand_199_nl), cfg_proc_precision_1_sva_st_108[1]);
  assign mux_1212_nl = MUX_s_1_2_2((mux_1211_nl), or_tmp_1992, cfg_proc_precision_1_sva_st_108[0]);
  assign mux_1213_nl = MUX_s_1_2_2((mux_1212_nl), (nand_46_nl), or_5189_cse);
  assign and_2784_nl = (~((cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[16:5]==12'b111111111111)))
      & or_5053_cse;
  assign mux_2276_nl = MUX_s_1_2_2((and_2784_nl), or_5053_cse, cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4);
  assign nor_2406_nl = ~(((~ cvt_14_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4)
      & (cvt_14_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[16:5]==12'b111111111111))
      | (~(or_5053_cse & or_400_cse_1 & (~(nor_2219_cse | (cfg_out_precision_1_sva_st_149!=2'b10)
      | FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2 | cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2
      | (cfg_out_precision_1_sva_st_113!=2'b10))))));
  assign mux_2277_nl = MUX_s_1_2_2((nor_2406_nl), nor_2099_cse, nor_50_cse);
  assign and_2782_nl = (~((cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[16:5]==12'b111111111111)))
      & or_5069_cse;
  assign mux_2278_nl = MUX_s_1_2_2((and_2782_nl), or_5069_cse, cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4);
  assign nor_2401_nl = ~(((~ cvt_15_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_6_tmp_4)
      & (cvt_15_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_3_tmp[16:5]==12'b111111111111))
      | (~(or_5069_cse & or_400_cse_1 & (~(nor_2219_cse | (cfg_out_precision_1_sva_st_149!=2'b10)
      | FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_3 | cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_svs_2
      | (cfg_out_precision_1_sva_st_113!=2'b10))))));
  assign mux_2279_nl = MUX_s_1_2_2((nor_2401_nl), nor_2099_cse, nor_50_cse);
  assign and_2780_nl = (~((cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_tmp[16:5]==12'b111111111111)))
      & or_5086_cse;
  assign mux_2280_nl = MUX_s_1_2_2((and_2780_nl), or_5086_cse, cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_8_tmp_4);
  assign nor_2396_nl = ~(((~ cvt_16_FpIntToFloat_17U_5U_10U_else_else_1_if_if_acc_8_tmp_4)
      & (cvt_16_FpIntToFloat_17U_5U_10U_else_int_mant_lshift_4_tmp[16:5]==12'b111111111111))
      | (~(or_5086_cse & (~(nor_151_cse | nor_2219_cse | (cfg_out_precision_1_sva_st_149!=2'b10)
      | FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_3 | cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_svs_2
      | (cfg_out_precision_1_sva_st_113!=2'b10))))));
  assign mux_2281_nl = MUX_s_1_2_2((nor_2396_nl), nor_2099_cse, nor_50_cse);
  assign and_223_nl = main_stage_v_2 & mux_417_cse;
  assign nor_1351_nl = ~((cfg_proc_precision_1_sva_st_108[1]) | (~ mux_tmp_1227));
  assign mux_1252_nl = MUX_s_1_2_2((nor_1351_nl), mux_tmp_1227, cfg_proc_precision_1_sva_st_108[0]);
  assign mux_1262_nl = MUX_s_1_2_2((mux_1252_nl), (and_223_nl), or_5189_cse);
  assign nor_1338_nl = ~((~ reg_chn_out_rsci_ld_core_psct_cse) | chn_out_rsci_bawt
      | (~ and_283_cse));
  assign mux_1265_nl = MUX_s_1_2_2(mux_tmp_1264, (nor_1338_nl), cfg_proc_precision_1_sva_st_101[1]);
  assign mux_1266_nl = MUX_s_1_2_2((mux_1265_nl), mux_tmp_1264, cfg_proc_precision_1_sva_st_101[0]);
  assign nor_2251_nl = ~((cfg_proc_precision_1_sva_st_65[1]) | (~ (cfg_out_precision_1_sva_st_113[1])));
  assign or_4857_nl = cvt_unequal_tmp_20 | (cfg_proc_precision_1_sva_st_65[0]);
  assign mux_2248_nl = MUX_s_1_2_2((nor_2251_nl), (cfg_out_precision_1_sva_st_113[1]),
      or_4857_nl);
  assign nor_2252_nl = ~((~ cvt_unequal_tmp_20) | (cfg_proc_precision_1_sva_st_65!=2'b10));
  assign mux_2249_nl = MUX_s_1_2_2((nor_2252_nl), (mux_2248_nl), cfg_out_precision_1_sva_st_113[0]);
  assign mux_1420_nl = MUX_s_1_2_2(or_5189_cse, (~ mux_tmp_1419), cfg_out_precision_1_sva_st_154[1]);
  assign mux_1421_nl = MUX_s_1_2_2((mux_1420_nl), or_5189_cse, or_4559_cse);
  assign mux_1423_nl = MUX_s_1_2_2((mux_1421_nl), or_5189_cse, nor_2150_cse);
  assign mux_1424_nl = MUX_s_1_2_2((mux_1423_nl), or_5189_cse, nor_8_cse);
  assign or_2251_nl = (cfg_out_precision_1_sva_st_154!=2'b10);
  assign mux_1425_nl = MUX_s_1_2_2(not_tmp_1709, (mux_1424_nl), or_2251_nl);
  assign mux_1426_nl = MUX_s_1_2_2(or_5189_cse, (mux_1425_nl), main_stage_v_1);
  assign mux_1427_nl = MUX_s_1_2_2(nand_tmp_48, (~ (mux_1426_nl)), or_4524_cse);
  assign mux_1428_nl = MUX_s_1_2_2(nand_tmp_48, (mux_1427_nl), chn_in_rsci_bawt);
  assign or_2242_nl = (cfg_out_precision_rsci_d!=2'b10);
  assign mux_1429_nl = MUX_s_1_2_2((mux_1428_nl), nand_tmp_48, or_2242_nl);
  assign nor_2113_nl = ~(nor_8_cse | (cfg_out_precision_1_sva_st_154[0]) | (~((cfg_out_precision_1_sva_st_154[1])
      & mux_1466_cse)));
  assign mux_1467_nl = MUX_s_1_2_2(main_stage_v_1, (nor_2113_nl), or_2289_cse);
  assign nor_1303_nl = ~((cfg_proc_precision_1_sva_st_89[1]) | (~ mux_tmp_1469));
  assign mux_1470_nl = MUX_s_1_2_2((nor_1303_nl), mux_tmp_1469, cfg_proc_precision_1_sva_st_89[0]);
  assign nor_1302_nl = ~(nor_50_cse | (cfg_out_precision_1_sva_st_149[0]) | (~((cfg_out_precision_1_sva_st_149[1])
      & (mux_1470_nl))));
  assign mux_1471_nl = MUX_s_1_2_2(main_stage_v_2, (nor_1302_nl), or_1587_cse);
  assign mux_1472_nl = MUX_s_1_2_2((mux_1471_nl), (mux_1467_nl), or_5189_cse);
  assign mux_1531_nl = MUX_s_1_2_2(or_tmp_2432, (~ chn_in_rsci_bawt), cfg_proc_precision_rsci_d[1]);
  assign or_2433_nl = (cfg_out_precision_rsci_d!=2'b01) | (cfg_proc_precision_rsci_d[0]);
  assign mux_1532_nl = MUX_s_1_2_2((mux_1531_nl), or_tmp_2432, or_2433_nl);
  assign mux_1533_nl = MUX_s_1_2_2(mux_tmp_189, (mux_1532_nl), or_5189_cse);
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_1_sva_2 = conv_u2u_4_5({FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_2_sva_mx0w0
      , (~ (chn_in_rsci_d_mxwt[23]))}) + 5'b1101;
  assign nor_1263_nl = ~(cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_itm_8_1
      | cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1 | (~ cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_tmp);
  assign nor_1264_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_st_2
      | cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_2
      | IsNaN_8U_23U_land_1_lpi_1_dfm_3 | cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_2
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_2
      | nand_164_cse);
  assign mux_1534_nl = MUX_s_1_2_2((nor_1264_nl), (nor_1263_nl), or_5189_cse);
  assign nor_1261_nl = ~((cvt_1_FpMantRNE_24U_11U_else_and_tmp & (cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_tmp==5'b11111))
      | (~ cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_itm_8_1) | cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1
      | (~ cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_itm_8_1) | (cfg_proc_precision_rsci_d!=2'b10)
      | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_tmp);
  assign nor_1262_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_st_2
      | (~ cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_st_2)
      | IsNaN_8U_23U_land_1_lpi_1_dfm_3 | (~ cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_svs_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_1_sva_2
      | nand_164_cse);
  assign mux_1535_nl = MUX_s_1_2_2((nor_1262_nl), (nor_1261_nl), or_5189_cse);
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_2_sva_2 = conv_u2u_4_5({FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_3_sva_mx0w0
      , (~ (chn_in_rsci_d_mxwt[55]))}) + 5'b1101;
  assign nor_1259_nl = ~(cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1
      | cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1 | (~ cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_1_tmp);
  assign nor_1260_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_st_2
      | cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2
      | IsNaN_8U_23U_land_2_lpi_1_dfm_3 | cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_2
      | nand_162_cse);
  assign mux_1536_nl = MUX_s_1_2_2((nor_1260_nl), (nor_1259_nl), or_5189_cse);
  assign nor_1257_nl = ~((cvt_2_FpMantRNE_24U_11U_else_and_1_tmp & (cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp==5'b11111))
      | (~ cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1) | cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1
      | (~ cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1) | (cfg_proc_precision_rsci_d!=2'b10)
      | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_1_tmp);
  assign nor_1258_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_st_2
      | (~ cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2)
      | IsNaN_8U_23U_land_2_lpi_1_dfm_3 | (~ cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_2_sva_2
      | nand_162_cse);
  assign mux_1537_nl = MUX_s_1_2_2((nor_1258_nl), (nor_1257_nl), or_5189_cse);
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_3_sva_2 = conv_u2u_4_5({FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_4_sva_mx0w0
      , (~ (chn_in_rsci_d_mxwt[87]))}) + 5'b1101;
  assign nor_1255_nl = ~(cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1
      | cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1 | (~ cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_2_tmp);
  assign nor_1256_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_st_2
      | cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2
      | IsNaN_8U_23U_land_3_lpi_1_dfm_3 | cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_2
      | nand_160_cse);
  assign mux_1538_nl = MUX_s_1_2_2((nor_1256_nl), (nor_1255_nl), or_5189_cse);
  assign nor_1253_nl = ~((cvt_3_FpMantRNE_24U_11U_else_and_1_tmp & (cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp==5'b11111))
      | (~ cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1) | cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1
      | (~ cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1) | (cfg_proc_precision_rsci_d!=2'b10)
      | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_2_tmp);
  assign nor_1254_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_st_2
      | (~ cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2)
      | IsNaN_8U_23U_land_3_lpi_1_dfm_3 | (~ cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_3_sva_2
      | nand_160_cse);
  assign mux_1539_nl = MUX_s_1_2_2((nor_1254_nl), (nor_1253_nl), or_5189_cse);
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_4_sva_2 = conv_u2u_4_5({FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_5_sva_mx0w0
      , (~ (chn_in_rsci_d_mxwt[119]))}) + 5'b1101;
  assign nor_1251_nl = ~(cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1
      | cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_3_tmp);
  assign nor_1252_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_st_2
      | cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2
      | IsNaN_8U_23U_land_4_lpi_1_dfm_3 | cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_2
      | nand_158_cse);
  assign mux_1540_nl = MUX_s_1_2_2((nor_1252_nl), (nor_1251_nl), or_5189_cse);
  assign nor_1249_nl = ~((cvt_4_FpMantRNE_24U_11U_else_and_2_tmp & (cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp==5'b11111))
      | (~ cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1) | cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1
      | (~ cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1) | (cfg_proc_precision_rsci_d!=2'b10)
      | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_3_tmp);
  assign nor_1250_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_st_2
      | (~ cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2)
      | IsNaN_8U_23U_land_4_lpi_1_dfm_3 | (~ cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_4_sva_2
      | nand_158_cse);
  assign mux_1541_nl = MUX_s_1_2_2((nor_1250_nl), (nor_1249_nl), or_5189_cse);
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_5_sva_2 = conv_u2u_4_5({FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_6_sva_mx0w0
      , (~ (chn_in_rsci_d_mxwt[151]))}) + 5'b1101;
  assign nor_1247_nl = ~((~ or_tmp_2466) | cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1
      | cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1 | (~ cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt));
  assign nor_1248_nl = ~((~ or_tmp_2469) | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_st_2
      | cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2
      | cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_2
      | nand_156_cse);
  assign mux_1542_nl = MUX_s_1_2_2((nor_1248_nl), (nor_1247_nl), or_5189_cse);
  assign nor_1245_nl = ~((cvt_5_FpMantRNE_24U_11U_else_and_1_tmp & (cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp==5'b11111))
      | (~(or_tmp_2466 & cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1
      & (~ cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1) & cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1
      & (cfg_proc_precision_rsci_d==2'b10) & chn_in_rsci_bawt)));
  assign nor_1246_nl = ~((~ or_tmp_2469) | (~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_st_2
      | (~ cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2)
      | (~ cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_5_sva_2
      | nand_156_cse);
  assign mux_1543_nl = MUX_s_1_2_2((nor_1246_nl), (nor_1245_nl), or_5189_cse);
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_6_sva_2 = conv_u2u_4_5({FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_7_sva_mx0w0
      , (~ (chn_in_rsci_d_mxwt[183]))}) + 5'b1101;
  assign nor_1243_nl = ~(cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1
      | cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_5_tmp);
  assign nor_1244_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_st_2
      | cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2
      | IsNaN_8U_23U_land_6_lpi_1_dfm_3 | cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_2
      | nand_153_cse);
  assign mux_1544_nl = MUX_s_1_2_2((nor_1244_nl), (nor_1243_nl), or_5189_cse);
  assign nor_1241_nl = ~((cvt_6_FpMantRNE_24U_11U_else_and_2_tmp & (cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp==5'b11111))
      | (~ cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1) | cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1
      | (~ cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1) | (cfg_proc_precision_rsci_d!=2'b10)
      | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_5_tmp);
  assign nor_1242_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_st_2
      | (~ cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2)
      | IsNaN_8U_23U_land_6_lpi_1_dfm_3 | (~ cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_6_sva_2
      | nand_153_cse);
  assign mux_1545_nl = MUX_s_1_2_2((nor_1242_nl), (nor_1241_nl), or_5189_cse);
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_7_sva_2 = conv_u2u_4_5({FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_8_sva_mx0w0
      , (~ (chn_in_rsci_d_mxwt[215]))}) + 5'b1101;
  assign nor_1239_nl = ~(cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1
      | cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_6_tmp);
  assign nor_1240_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_st_2
      | cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2
      | IsNaN_8U_23U_land_7_lpi_1_dfm_3 | cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_2
      | nand_151_cse);
  assign mux_1546_nl = MUX_s_1_2_2((nor_1240_nl), (nor_1239_nl), or_5189_cse);
  assign nor_1237_nl = ~((cvt_7_FpMantRNE_24U_11U_else_and_2_tmp & (cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp==5'b11111))
      | (~ cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1) | cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1
      | (~ cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1) | (cfg_proc_precision_rsci_d!=2'b10)
      | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_6_tmp);
  assign nor_1238_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_st_2
      | (~ cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2)
      | IsNaN_8U_23U_land_7_lpi_1_dfm_3 | (~ cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_7_sva_2
      | nand_151_cse);
  assign mux_1547_nl = MUX_s_1_2_2((nor_1238_nl), (nor_1237_nl), or_5189_cse);
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_8_sva_2 = conv_u2u_4_5({FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_9_sva_mx0w0
      , (~ (chn_in_rsci_d_mxwt[247]))}) + 5'b1101;
  assign nor_1235_nl = ~(cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1
      | cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 | (~ cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_7_tmp);
  assign nor_1236_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_st_2
      | cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2
      | IsNaN_8U_23U_land_8_lpi_1_dfm_3 | cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_2
      | nand_149_cse);
  assign mux_1548_nl = MUX_s_1_2_2((nor_1236_nl), (nor_1235_nl), or_5189_cse);
  assign nor_1233_nl = ~((cvt_8_FpMantRNE_24U_11U_else_and_3_tmp & (cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp==5'b11111))
      | (~ cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1) | cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1
      | (~ cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1) | (cfg_proc_precision_rsci_d!=2'b10)
      | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_7_tmp);
  assign nor_1234_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_st_2
      | (~ cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2)
      | IsNaN_8U_23U_land_8_lpi_1_dfm_3 | (~ cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_8_sva_2
      | nand_149_cse);
  assign mux_1549_nl = MUX_s_1_2_2((nor_1234_nl), (nor_1233_nl), or_5189_cse);
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_9_sva_2 = conv_u2u_4_5({FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_10_sva_mx0w0
      , (~ (chn_in_rsci_d_mxwt[279]))}) + 5'b1101;
  assign nor_1231_nl = ~(cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1
      | cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1 | (~ cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_8_tmp);
  assign nor_1232_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_st_2
      | cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2
      | IsNaN_8U_23U_land_9_lpi_1_dfm_3 | cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_2
      | nand_147_cse);
  assign mux_1550_nl = MUX_s_1_2_2((nor_1232_nl), (nor_1231_nl), or_5189_cse);
  assign nor_1229_nl = ~((cvt_9_FpMantRNE_24U_11U_else_and_1_tmp & (cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_1_tmp==5'b11111))
      | (~ cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1) | cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1
      | (~ cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1) | (cfg_proc_precision_rsci_d!=2'b10)
      | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_8_tmp);
  assign nor_1230_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_st_2
      | (~ cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_st_2)
      | IsNaN_8U_23U_land_9_lpi_1_dfm_3 | (~ cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_1_svs_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_9_sva_2
      | nand_147_cse);
  assign mux_1551_nl = MUX_s_1_2_2((nor_1230_nl), (nor_1229_nl), or_5189_cse);
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_10_sva_2 = conv_u2u_4_5({FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_11_sva_mx0w0
      , (~ (chn_in_rsci_d_mxwt[311]))}) + 5'b1101;
  assign nor_1227_nl = ~(cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1
      | cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_9_tmp);
  assign nor_1228_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_st_2
      | cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2
      | IsNaN_8U_23U_land_10_lpi_1_dfm_3 | cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_2
      | nand_145_cse);
  assign mux_1552_nl = MUX_s_1_2_2((nor_1228_nl), (nor_1227_nl), or_5189_cse);
  assign nor_1225_nl = ~((cvt_10_FpMantRNE_24U_11U_else_and_2_tmp & (cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp==5'b11111))
      | (~ cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1) | cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1
      | (~ cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1) | (cfg_proc_precision_rsci_d!=2'b10)
      | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_9_tmp);
  assign nor_1226_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_st_2
      | (~ cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2)
      | IsNaN_8U_23U_land_10_lpi_1_dfm_3 | (~ cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_10_sva_2
      | nand_145_cse);
  assign mux_1553_nl = MUX_s_1_2_2((nor_1226_nl), (nor_1225_nl), or_5189_cse);
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_11_sva_2 = conv_u2u_4_5({FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_12_sva_mx0w0
      , (~ (chn_in_rsci_d_mxwt[343]))}) + 5'b1101;
  assign nor_1223_nl = ~(cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1
      | cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_10_tmp);
  assign nor_1224_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_st_2
      | cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2
      | IsNaN_8U_23U_land_11_lpi_1_dfm_3 | cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_2
      | nand_143_cse);
  assign mux_1554_nl = MUX_s_1_2_2((nor_1224_nl), (nor_1223_nl), or_5189_cse);
  assign nor_1221_nl = ~((cvt_11_FpMantRNE_24U_11U_else_and_2_tmp & (cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp==5'b11111))
      | (~ cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1) | cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1
      | (~ cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1) | (cfg_proc_precision_rsci_d!=2'b10)
      | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_10_tmp);
  assign nor_1222_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_st_2
      | (~ cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2)
      | IsNaN_8U_23U_land_11_lpi_1_dfm_3 | (~ cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_11_sva_2
      | nand_143_cse);
  assign mux_1555_nl = MUX_s_1_2_2((nor_1222_nl), (nor_1221_nl), or_5189_cse);
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_12_sva_2 = conv_u2u_4_5({FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_13_sva_mx0w0
      , (~ (chn_in_rsci_d_mxwt[375]))}) + 5'b1101;
  assign nor_1219_nl = ~(cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1
      | cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 | (~ cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_11_tmp);
  assign nor_1220_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_st_2
      | cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2
      | IsNaN_8U_23U_land_12_lpi_1_dfm_3 | cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_2
      | nand_141_cse);
  assign mux_1556_nl = MUX_s_1_2_2((nor_1220_nl), (nor_1219_nl), or_5189_cse);
  assign nor_1217_nl = ~((cvt_12_FpMantRNE_24U_11U_else_and_3_tmp & (cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp==5'b11111))
      | (~ cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1) | cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1
      | (~ cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1) | (cfg_proc_precision_rsci_d!=2'b10)
      | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_11_tmp);
  assign nor_1218_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_st_2
      | (~ cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2)
      | IsNaN_8U_23U_land_12_lpi_1_dfm_3 | (~ cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_12_sva_2
      | nand_141_cse);
  assign mux_1557_nl = MUX_s_1_2_2((nor_1218_nl), (nor_1217_nl), or_5189_cse);
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_13_sva_2 = conv_u2u_4_5({FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_14_sva_mx0w0
      , (~ (chn_in_rsci_d_mxwt[407]))}) + 5'b1101;
  assign nor_1215_nl = ~(cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1
      | cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_12_tmp);
  assign nor_1216_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_st_2
      | cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2
      | IsNaN_8U_23U_land_13_lpi_1_dfm_3 | cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_2
      | nand_139_cse);
  assign mux_1558_nl = MUX_s_1_2_2((nor_1216_nl), (nor_1215_nl), or_5189_cse);
  assign nor_1213_nl = ~((cvt_13_FpMantRNE_24U_11U_else_and_2_tmp & (cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_2_tmp==5'b11111))
      | (~ cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1) | cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1
      | (~ cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1) | (cfg_proc_precision_rsci_d!=2'b10)
      | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_12_tmp);
  assign nor_1214_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_st_2
      | (~ cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_st_2)
      | IsNaN_8U_23U_land_13_lpi_1_dfm_3 | (~ cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_2_svs_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_13_sva_2
      | nand_139_cse);
  assign mux_1559_nl = MUX_s_1_2_2((nor_1214_nl), (nor_1213_nl), or_5189_cse);
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_14_sva_2 = conv_u2u_4_5({FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_15_sva_mx0w0
      , (~ (chn_in_rsci_d_mxwt[439]))}) + 5'b1101;
  assign nor_1211_nl = ~(cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1
      | cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 | (~ cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_13_tmp);
  assign nor_1212_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_st_2
      | cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2
      | IsNaN_8U_23U_land_14_lpi_1_dfm_3 | cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_2
      | nand_137_cse);
  assign mux_1560_nl = MUX_s_1_2_2((nor_1212_nl), (nor_1211_nl), or_5189_cse);
  assign nor_1209_nl = ~((cvt_14_FpMantRNE_24U_11U_else_and_3_tmp & (cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp==5'b11111))
      | (~ cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1) | cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1
      | (~ cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1) | (cfg_proc_precision_rsci_d!=2'b10)
      | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_13_tmp);
  assign nor_1210_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_st_2
      | (~ cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2)
      | IsNaN_8U_23U_land_14_lpi_1_dfm_3 | (~ cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_14_sva_2
      | nand_137_cse);
  assign mux_1561_nl = MUX_s_1_2_2((nor_1210_nl), (nor_1209_nl), or_5189_cse);
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_15_sva_2 = conv_u2u_4_5({FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_16_sva_mx0w0
      , (~ (chn_in_rsci_d_mxwt[471]))}) + 5'b1101;
  assign nor_1207_nl = ~(cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1
      | cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 | (~ cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_14_tmp);
  assign nor_1208_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_st_2
      | cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2
      | IsNaN_8U_23U_land_15_lpi_1_dfm_3 | cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_2
      | nand_135_cse);
  assign mux_1562_nl = MUX_s_1_2_2((nor_1208_nl), (nor_1207_nl), or_5189_cse);
  assign nor_1205_nl = ~((cvt_15_FpMantRNE_24U_11U_else_and_3_tmp & (cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_3_tmp==5'b11111))
      | (~ cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1) | cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1
      | (~ cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1) | (cfg_proc_precision_rsci_d!=2'b10)
      | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_14_tmp);
  assign nor_1206_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_st_2
      | (~ cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_st_2)
      | IsNaN_8U_23U_land_15_lpi_1_dfm_3 | (~ cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_3_svs_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_15_sva_2
      | nand_135_cse);
  assign mux_1563_nl = MUX_s_1_2_2((nor_1206_nl), (nor_1205_nl), or_5189_cse);
  assign nl_FpMantDecShiftRight_23U_8U_10U_guard_mask_acc_1_psp_sva_2 = conv_u2u_4_5({FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_i_shift_acc_psp_1_sva_mx0w0
      , (~ (chn_in_rsci_d_mxwt[503]))}) + 5'b1101;
  assign nor_1203_nl = ~(cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_itm_8_1
      | cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_itm_7_1 | (~ cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_itm_8_1)
      | (cfg_proc_precision_rsci_d!=2'b10) | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_15_tmp);
  assign nor_1204_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_2
      | cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_st_2
      | IsNaN_8U_23U_land_lpi_1_dfm_3 | cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_2
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_2
      | nand_133_cse);
  assign mux_1564_nl = MUX_s_1_2_2((nor_1204_nl), (nor_1203_nl), or_5189_cse);
  assign nor_1201_nl = ~((cvt_16_FpMantRNE_24U_11U_else_and_4_tmp & (cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_else_if_acc_4_tmp==5'b11111))
      | (~ cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_itm_8_1) | cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_itm_7_1
      | (~ cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_itm_8_1) | (cfg_proc_precision_rsci_d!=2'b10)
      | (~ chn_in_rsci_bawt) | IsNaN_8U_23U_IsNaN_8U_23U_nor_15_tmp);
  assign nor_1202_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64!=2'b10)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_st_2
      | (~ cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_st_2)
      | IsNaN_8U_23U_land_lpi_1_dfm_3 | (~ cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_8_4_svs_2)
      | FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_slc_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_7_mdf_sva_2
      | nand_133_cse);
  assign mux_1565_nl = MUX_s_1_2_2((nor_1202_nl), (nor_1201_nl), or_5189_cse);
  assign mux_1567_nl = MUX_s_1_2_2(or_tmp_2569, mux_tmp_1566, cvt_16_FpMantRNE_24U_11U_else_and_4_tmp);
  assign mux_1568_nl = MUX_s_1_2_2(or_tmp_2569, mux_tmp_1566, cvt_16_FpMantRNE_24U_11U_else_and_4_svs);
  assign nor_597_nl = ~((~ cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_4_itm_8_1)
      | cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_4_itm_7_1 | (~ cvt_16_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_4_itm_8_1));
  assign mux_1569_nl = MUX_s_1_2_2((mux_1568_nl), (mux_1567_nl), nor_597_nl);
  assign mux_1571_nl = MUX_s_1_2_2(or_tmp_2571, mux_tmp_1570, cvt_15_FpMantRNE_24U_11U_else_and_3_tmp);
  assign mux_1572_nl = MUX_s_1_2_2(or_tmp_2571, mux_tmp_1570, cvt_15_FpMantRNE_24U_11U_else_and_3_svs);
  assign nor_598_nl = ~((~ cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1)
      | cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 | (~ cvt_15_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1));
  assign mux_1573_nl = MUX_s_1_2_2((mux_1572_nl), (mux_1571_nl), nor_598_nl);
  assign mux_1575_nl = MUX_s_1_2_2(or_tmp_2573, mux_tmp_1574, cvt_14_FpMantRNE_24U_11U_else_and_3_tmp);
  assign mux_1576_nl = MUX_s_1_2_2(or_tmp_2573, mux_tmp_1574, cvt_14_FpMantRNE_24U_11U_else_and_3_svs);
  assign nor_599_nl = ~((~ cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1)
      | cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 | (~ cvt_14_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1));
  assign mux_1577_nl = MUX_s_1_2_2((mux_1576_nl), (mux_1575_nl), nor_599_nl);
  assign mux_1579_nl = MUX_s_1_2_2(or_tmp_2575, mux_tmp_1578, cvt_13_FpMantRNE_24U_11U_else_and_2_tmp);
  assign mux_1580_nl = MUX_s_1_2_2(or_tmp_2575, mux_tmp_1578, cvt_13_FpMantRNE_24U_11U_else_and_2_svs);
  assign nor_600_nl = ~((~ cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1)
      | cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_13_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1));
  assign mux_1581_nl = MUX_s_1_2_2((mux_1580_nl), (mux_1579_nl), nor_600_nl);
  assign mux_1583_nl = MUX_s_1_2_2(or_tmp_2577, mux_tmp_1582, cvt_12_FpMantRNE_24U_11U_else_and_3_tmp);
  assign mux_1584_nl = MUX_s_1_2_2(or_tmp_2577, mux_tmp_1582, cvt_12_FpMantRNE_24U_11U_else_and_3_svs);
  assign nor_601_nl = ~((~ cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1)
      | cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 | (~ cvt_12_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1));
  assign mux_1585_nl = MUX_s_1_2_2((mux_1584_nl), (mux_1583_nl), nor_601_nl);
  assign mux_1587_nl = MUX_s_1_2_2(or_tmp_2579, mux_tmp_1586, cvt_11_FpMantRNE_24U_11U_else_and_2_tmp);
  assign mux_1588_nl = MUX_s_1_2_2(or_tmp_2579, mux_tmp_1586, cvt_11_FpMantRNE_24U_11U_else_and_2_svs);
  assign nor_602_nl = ~((~ cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1)
      | cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_11_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1));
  assign mux_1589_nl = MUX_s_1_2_2((mux_1588_nl), (mux_1587_nl), nor_602_nl);
  assign and_2243_nl = cvt_10_FpMantRNE_24U_11U_else_and_2_tmp & (cfg_proc_precision_rsci_d==2'b10)
      & chn_in_rsci_bawt;
  assign and_2162_nl = cvt_10_FpMantRNE_24U_11U_else_and_2_svs & (cfg_proc_precision_rsci_d==2'b10)
      & chn_in_rsci_bawt;
  assign nor_603_nl = ~((~ cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1)
      | cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_10_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1));
  assign mux_1590_nl = MUX_s_1_2_2((and_2162_nl), (and_2243_nl), nor_603_nl);
  assign nor_1200_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64[0])
      | (~((cfg_proc_precision_1_sva_st_64[1]) & cvt_10_FpMantRNE_24U_11U_else_and_2_svs_2)));
  assign mux_1591_nl = MUX_s_1_2_2((nor_1200_nl), (mux_1590_nl), or_5189_cse);
  assign mux_1593_nl = MUX_s_1_2_2(or_tmp_2588, mux_tmp_1592, cvt_9_FpMantRNE_24U_11U_else_and_1_tmp);
  assign mux_1594_nl = MUX_s_1_2_2(or_tmp_2588, mux_tmp_1592, cvt_9_FpMantRNE_24U_11U_else_and_1_svs);
  assign nor_605_nl = ~((~ cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1)
      | cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1 | (~ cvt_9_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1));
  assign mux_1595_nl = MUX_s_1_2_2((mux_1594_nl), (mux_1593_nl), nor_605_nl);
  assign mux_1597_nl = MUX_s_1_2_2(or_tmp_2590, mux_tmp_1596, cvt_8_FpMantRNE_24U_11U_else_and_3_tmp);
  assign mux_1598_nl = MUX_s_1_2_2(or_tmp_2590, mux_tmp_1596, cvt_8_FpMantRNE_24U_11U_else_and_3_svs);
  assign nor_606_nl = ~((~ cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_3_itm_8_1)
      | cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_3_itm_7_1 | (~ cvt_8_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_3_itm_8_1));
  assign mux_1599_nl = MUX_s_1_2_2((mux_1598_nl), (mux_1597_nl), nor_606_nl);
  assign mux_1601_nl = MUX_s_1_2_2(or_tmp_2595, mux_tmp_1600, cvt_7_FpMantRNE_24U_11U_else_and_2_tmp);
  assign mux_1602_nl = MUX_s_1_2_2(or_tmp_2595, mux_tmp_1600, cvt_7_FpMantRNE_24U_11U_else_and_2_svs);
  assign nor_607_nl = ~((~ cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1)
      | cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_7_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1));
  assign mux_1603_nl = MUX_s_1_2_2((mux_1602_nl), (mux_1601_nl), nor_607_nl);
  assign and_nl = cvt_6_FpMantRNE_24U_11U_else_and_2_tmp & (cfg_proc_precision_rsci_d==2'b10)
      & chn_in_rsci_bawt;
  assign and_2161_nl = cvt_6_FpMantRNE_24U_11U_else_and_2_svs & (cfg_proc_precision_rsci_d==2'b10)
      & chn_in_rsci_bawt;
  assign nor_608_nl = ~((~ cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1)
      | cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_6_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1));
  assign mux_1604_nl = MUX_s_1_2_2((and_2161_nl), (and_nl), nor_608_nl);
  assign nor_1198_nl = ~((~ main_stage_v_1) | (cfg_proc_precision_1_sva_st_64[0])
      | (~((cfg_proc_precision_1_sva_st_64[1]) & cvt_6_FpMantRNE_24U_11U_else_and_2_svs_2)));
  assign mux_1605_nl = MUX_s_1_2_2((nor_1198_nl), (mux_1604_nl), or_5189_cse);
  assign mux_1607_nl = MUX_s_1_2_2(or_tmp_2604, mux_tmp_1606, cvt_5_FpMantRNE_24U_11U_else_and_1_tmp);
  assign mux_1608_nl = MUX_s_1_2_2(or_tmp_2604, mux_tmp_1606, cvt_5_FpMantRNE_24U_11U_else_and_1_svs);
  assign nor_610_nl = ~((~ cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1)
      | cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1 | (~ cvt_5_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1));
  assign mux_1609_nl = MUX_s_1_2_2((mux_1608_nl), (mux_1607_nl), nor_610_nl);
  assign mux_1611_nl = MUX_s_1_2_2(or_tmp_2606, mux_tmp_1610, cvt_4_FpMantRNE_24U_11U_else_and_2_tmp);
  assign mux_1612_nl = MUX_s_1_2_2(or_tmp_2606, mux_tmp_1610, cvt_4_FpMantRNE_24U_11U_else_and_2_svs);
  assign nor_611_nl = ~((~ cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_2_itm_8_1)
      | cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_2_itm_7_1 | (~ cvt_4_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_2_itm_8_1));
  assign mux_1613_nl = MUX_s_1_2_2((mux_1612_nl), (mux_1611_nl), nor_611_nl);
  assign mux_1615_nl = MUX_s_1_2_2(or_tmp_2608, mux_tmp_1614, cvt_3_FpMantRNE_24U_11U_else_and_1_tmp);
  assign mux_1616_nl = MUX_s_1_2_2(or_tmp_2608, mux_tmp_1614, cvt_3_FpMantRNE_24U_11U_else_and_1_svs);
  assign nor_612_nl = ~((~ cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1)
      | cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1 | (~ cvt_3_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1));
  assign mux_1617_nl = MUX_s_1_2_2((mux_1616_nl), (mux_1615_nl), nor_612_nl);
  assign mux_1619_nl = MUX_s_1_2_2(or_tmp_2610, mux_tmp_1618, cvt_2_FpMantRNE_24U_11U_else_and_1_tmp);
  assign mux_1620_nl = MUX_s_1_2_2(or_tmp_2610, mux_tmp_1618, cvt_2_FpMantRNE_24U_11U_else_and_1_svs);
  assign nor_613_nl = ~((~ cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_1_itm_8_1)
      | cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_1_itm_7_1 | (~ cvt_2_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_1_itm_8_1));
  assign mux_1621_nl = MUX_s_1_2_2((mux_1620_nl), (mux_1619_nl), nor_613_nl);
  assign mux_1623_nl = MUX_s_1_2_2(or_tmp_2612, mux_tmp_1622, cvt_1_FpMantRNE_24U_11U_else_and_tmp);
  assign mux_1624_nl = MUX_s_1_2_2(or_tmp_2612, mux_tmp_1622, cvt_1_FpMantRNE_24U_11U_else_and_svs);
  assign nor_614_nl = ~((~ cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_acc_itm_8_1) | cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_if_acc_itm_7_1
      | (~ cvt_1_FpWidthDec_8U_23U_5U_10U_1U_1U_else_else_acc_itm_8_1));
  assign mux_1625_nl = MUX_s_1_2_2((mux_1624_nl), (mux_1623_nl), nor_614_nl);
  assign and_2160_nl = cfg_mode_eql_1_sva_5 & main_stage_v_2;
  assign mux_1627_nl = MUX_s_1_2_2((and_2160_nl), and_2239_cse, or_5189_cse);
  assign IsNaN_5U_10U_nor_nl = ~((FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_1_lpi_1_dfm_5_mx0!=10'b0000000000));
  assign mux_1632_nl = MUX_s_1_2_2(mux_tmp_719, nor_1185_cse, cfg_proc_precision_1_sva_st_64[1]);
  assign mux_1633_nl = MUX_s_1_2_2((mux_1632_nl), mux_tmp_719, cfg_proc_precision_1_sva_st_64[0]);
  assign mux_1638_nl = MUX_s_1_2_2(mux_767_cse, nor_1186_cse, cfg_proc_precision_1_sva_st_65[1]);
  assign mux_1639_nl = MUX_s_1_2_2((mux_1638_nl), mux_767_cse, cfg_proc_precision_1_sva_st_65[0]);
  assign mux_1640_nl = MUX_s_1_2_2((mux_1639_nl), (mux_1633_nl), or_5189_cse);
  assign IsNaN_5U_10U_IsNaN_5U_10U_nand_nl = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_7_4_mx0w0
      & (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_1_lpi_1_dfm_7_3_0_mx0w0==4'b1111));
  assign mux_1643_nl = MUX_s_1_2_2(mux_1460_cse, nor_1185_cse, cfg_proc_precision_1_sva_st_64[1]);
  assign mux_1644_nl = MUX_s_1_2_2((mux_1643_nl), mux_1460_cse, cfg_proc_precision_1_sva_st_64[0]);
  assign mux_1647_nl = MUX_s_1_2_2(mux_1463_cse, nor_1186_cse, cfg_proc_precision_1_sva_st_65[1]);
  assign mux_1648_nl = MUX_s_1_2_2((mux_1647_nl), mux_1463_cse, cfg_proc_precision_1_sva_st_65[0]);
  assign mux_1649_nl = MUX_s_1_2_2((mux_1648_nl), (mux_1644_nl), or_5189_cse);
  assign IsNaN_5U_10U_nor_1_nl = ~((FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_2_lpi_1_dfm_5_mx0!=10'b0000000000));
  assign mux_1658_nl = MUX_s_1_2_2(mux_660_cse, nor_1186_cse, cfg_proc_precision_1_sva_st_65[1]);
  assign mux_1659_nl = MUX_s_1_2_2((mux_1658_nl), mux_660_cse, cfg_proc_precision_1_sva_st_65[0]);
  assign mux_1660_nl = MUX_s_1_2_2((mux_1659_nl), mux_1654_cse, or_5189_cse);
  assign IsNaN_5U_10U_IsNaN_5U_10U_nand_1_nl = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_7_4_mx0w0
      & (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_2_lpi_1_dfm_7_3_0_mx0w0==4'b1111));
  assign mux_1661_nl = MUX_s_1_2_2(nor_1309_cse, nor_1185_cse, nor_8_cse);
  assign mux_1662_nl = MUX_s_1_2_2(nor_1310_cse, nor_1186_cse, nor_50_cse);
  assign mux_1663_nl = MUX_s_1_2_2((mux_1662_nl), (mux_1661_nl), or_5189_cse);
  assign IsNaN_5U_10U_nor_14_nl = ~((FpWidthDec_8U_23U_5U_10U_1U_1U_o_mant_15_lpi_1_dfm_5_mx0!=10'b0000000000));
  assign mux_1672_nl = MUX_s_1_2_2(mux_786_cse_1, nor_1186_cse, cfg_proc_precision_1_sva_st_65[1]);
  assign mux_1673_nl = MUX_s_1_2_2((mux_1672_nl), mux_786_cse_1, cfg_proc_precision_1_sva_st_65[0]);
  assign mux_1674_nl = MUX_s_1_2_2((mux_1673_nl), mux_1654_cse, or_5189_cse);
  assign IsNaN_5U_10U_IsNaN_5U_10U_nand_14_nl = ~(FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_7_4_mx0w0
      & (FpWidthDec_8U_23U_5U_10U_1U_1U_o_expo_15_lpi_1_dfm_7_3_0_mx0w0==4'b1111));
  assign mux_1683_nl = MUX_s_1_2_2(mux_201_cse, nor_1186_cse, cfg_proc_precision_1_sva_st_65[1]);
  assign mux_1684_nl = MUX_s_1_2_2((mux_1683_nl), mux_201_cse, cfg_proc_precision_1_sva_st_65[0]);
  assign mux_1685_nl = MUX_s_1_2_2((mux_1684_nl), mux_1654_cse, or_5189_cse);
  assign or_724_nl = main_stage_v_2 | (~ mux_tmp_129);
  assign mux_449_nl = MUX_s_1_2_2((or_724_nl), or_5379_cse, or_5189_cse);
  assign or_733_nl = main_stage_v_2 | (~ and_tmp_18);
  assign mux_454_nl = MUX_s_1_2_2((or_733_nl), or_5379_cse, or_5189_cse);
  assign or_1118_nl = main_stage_v_2 | (~ mux_tmp_151);
  assign mux_770_nl = MUX_s_1_2_2((or_1118_nl), or_5379_cse, or_5189_cse);
  assign or_1134_nl = main_stage_v_2 | (~ and_tmp_33);
  assign mux_789_nl = MUX_s_1_2_2((or_1134_nl), or_5379_cse, or_5189_cse);
  assign or_1145_nl = (cfg_proc_precision_1_sva_st_101[0]) | (~((cfg_proc_precision_1_sva_st_101[1])
      & mux_tmp_455));
  assign mux_798_nl = MUX_s_1_2_2((~ and_1386_cse), (or_1145_nl), main_stage_v_2);
  assign mux_799_nl = MUX_s_1_2_2((mux_798_nl), or_5379_cse, or_5189_cse);
  assign mux_92_nl = MUX_s_1_2_2(and_dcpl_3, or_186_cse, or_183_cse_1);
  assign mux_801_nl = MUX_s_1_2_2((~ and_2186_cse), (mux_92_nl), main_stage_v_1);
  assign mux_207_nl = MUX_s_1_2_2(or_tmp_389, (~ or_4862_cse), cfg_proc_precision_1_sva_st_101[1]);
  assign mux_208_nl = MUX_s_1_2_2((mux_207_nl), or_tmp_389, cfg_proc_precision_1_sva_st_101[0]);
  assign mux_802_nl = MUX_s_1_2_2((~ and_tmp_11), (mux_208_nl), main_stage_v_2);
  assign mux_803_nl = MUX_s_1_2_2((mux_802_nl), (mux_801_nl), or_5189_cse);
  assign or_2688_nl = (~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp | (~ mux_344_cse);
  assign or_2691_nl = nor_2219_cse | (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | cvt_2_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 |
      nor_50_cse;
  assign mux_1687_nl = MUX_s_1_2_2((or_2691_nl), (or_2688_nl), or_5189_cse);
  assign or_2696_nl = (~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp | (~ mux_344_cse);
  assign or_2699_nl = nor_2219_cse | (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | cvt_3_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 |
      nor_50_cse;
  assign mux_1689_nl = MUX_s_1_2_2((or_2699_nl), (or_2696_nl), or_5189_cse);
  assign or_2705_nl = (~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_4_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp | (~ mux_474_cse);
  assign or_2709_nl = nor_151_cse | nor_2219_cse | (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | FpIntToFloat_17U_5U_10U_is_inf_4_lpi_1_dfm_3 | nor_50_cse;
  assign mux_1692_nl = MUX_s_1_2_2((or_2709_nl), (or_2705_nl), or_5189_cse);
  assign or_2714_nl = (~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp | (~ mux_344_cse);
  assign or_2717_nl = nor_2219_cse | (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | cvt_5_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 |
      nor_50_cse;
  assign mux_1694_nl = MUX_s_1_2_2((or_2717_nl), (or_2714_nl), or_5189_cse);
  assign or_2723_nl = (~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_6_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp | (~ mux_344_cse);
  assign or_2727_nl = nor_151_cse | nor_2219_cse | (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | FpIntToFloat_17U_5U_10U_is_inf_6_lpi_1_dfm_3 | nor_50_cse;
  assign mux_1697_nl = MUX_s_1_2_2((or_2727_nl), (or_2723_nl), or_5189_cse);
  assign or_2733_nl = (~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_7_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp | (~ mux_344_cse);
  assign or_2737_nl = nor_151_cse | nor_2219_cse | (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | FpIntToFloat_17U_5U_10U_is_inf_7_lpi_1_dfm_3 | nor_50_cse;
  assign mux_1700_nl = MUX_s_1_2_2((or_2737_nl), (or_2733_nl), or_5189_cse);
  assign or_2744_nl = (~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_8_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp | (~ mux_344_cse);
  assign or_2749_nl = nor_151_cse | nor_2219_cse | (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | FpIntToFloat_17U_5U_10U_is_inf_8_lpi_1_dfm_3 | nor_50_cse;
  assign mux_1704_nl = MUX_s_1_2_2((or_2749_nl), (or_2744_nl), or_5189_cse);
  assign or_2754_nl = (~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_tmp | (~ mux_344_cse);
  assign or_2758_nl = (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | cvt_9_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_1_svs_st_2 |
      (~ mux_1126_cse);
  assign mux_1707_nl = MUX_s_1_2_2((or_2758_nl), (or_2754_nl), or_5189_cse);
  assign or_2764_nl = (~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_10_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp | (~
      mux_474_cse);
  assign or_2768_nl = nor_151_cse | (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | FpIntToFloat_17U_5U_10U_is_inf_10_lpi_1_dfm_3 | (~ mux_1126_cse);
  assign mux_1711_nl = MUX_s_1_2_2((or_2768_nl), (or_2764_nl), or_5189_cse);
  assign or_2774_nl = (~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_11_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp | (~
      mux_474_cse);
  assign or_2778_nl = nor_151_cse | (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | FpIntToFloat_17U_5U_10U_is_inf_11_lpi_1_dfm_3 | (~ mux_1126_cse);
  assign mux_1715_nl = MUX_s_1_2_2((or_2778_nl), (or_2774_nl), or_5189_cse);
  assign or_2784_nl = (~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_13_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_2_tmp | (~
      mux_474_cse);
  assign or_2789_nl = (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | FpIntToFloat_17U_5U_10U_is_inf_13_lpi_1_dfm_3 | (~ mux_382_cse);
  assign mux_1720_nl = MUX_s_1_2_2((or_2789_nl), (or_2784_nl), or_5189_cse);
  assign or_2796_nl = (~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_14_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp | (~
      mux_474_cse);
  assign or_2802_nl = (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | FpIntToFloat_17U_5U_10U_is_inf_14_lpi_1_dfm_2 | (~ mux_417_cse);
  assign mux_1727_nl = MUX_s_1_2_2((or_2802_nl), (or_2796_nl), or_5189_cse);
  assign or_2809_nl = (~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_15_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_3_tmp | (~
      mux_474_cse);
  assign or_2815_nl = (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | FpIntToFloat_17U_5U_10U_is_inf_15_lpi_1_dfm_3 | (~ mux_417_cse);
  assign mux_1734_nl = MUX_s_1_2_2((or_2815_nl), (or_2809_nl), or_5189_cse);
  assign or_2823_nl = (~ main_stage_v_1) | (cfg_out_precision_1_sva_st_154!=2'b10)
      | cvt_16_FpIntToFloat_17U_5U_10U_FpIntToFloat_17U_5U_10U_if_nor_4_tmp | (~
      mux_344_cse);
  assign or_2830_nl = (~ main_stage_v_2) | (cfg_out_precision_1_sva_st_149!=2'b10)
      | FpIntToFloat_17U_5U_10U_is_inf_lpi_1_dfm_3 | (~ mux_417_cse);
  assign mux_1743_nl = MUX_s_1_2_2((or_2830_nl), (or_2823_nl), or_5189_cse);
  assign mux_1412_nl = MUX_s_1_2_2(mux_tmp_1409, (~ mux_1437_cse), cfg_out_precision_1_sva_st_154[1]);
  assign mux_1413_nl = MUX_s_1_2_2((mux_1412_nl), mux_tmp_1409, or_4559_cse);
  assign mux_1414_nl = MUX_s_1_2_2((mux_1413_nl), mux_tmp_1409, nor_2150_cse);
  assign mux_1415_nl = MUX_s_1_2_2((mux_1414_nl), mux_tmp_1409, nor_8_cse);
  assign mux_121_nl = MUX_s_1_2_2(or_tmp_218, or_tmp_213, or_5189_cse);
  assign or_236_nl = (cfg_out_precision_1_sva_st_154!=2'b10) | (~ mux_tmp_129);
  assign mux_131_nl = MUX_s_1_2_2((or_236_nl), or_tmp_213, or_5189_cse);
  assign or_263_nl = (cfg_out_precision_1_sva_st_154[0]) | (~((cfg_out_precision_1_sva_st_154[1])
      & and_tmp_16));
  assign mux_143_nl = MUX_s_1_2_2((or_263_nl), or_tmp_213, or_5189_cse);
  assign or_270_nl = (cfg_out_precision_1_sva_st_154!=2'b10) | (~ and_tmp_33);
  assign mux_150_nl = MUX_s_1_2_2((or_270_nl), or_tmp_213, or_5189_cse);
  assign or_275_nl = (cfg_out_precision_1_sva_st_154!=2'b10) | (~ mux_tmp_151);
  assign mux_153_nl = MUX_s_1_2_2((or_275_nl), or_tmp_213, or_5189_cse);
  function [0:0] MUX1HOT_s_1_1_2;
    input [0:0] input_0;
    input [0:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    MUX1HOT_s_1_1_2 = result;
  end
  endfunction
  function [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction
  function [0:0] MUX1HOT_s_1_5_2;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [4:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction
  function [14:0] MUX1HOT_v_15_3_2;
    input [14:0] input_2;
    input [14:0] input_1;
    input [14:0] input_0;
    input [2:0] sel;
    reg [14:0] result;
  begin
    result = input_0 & {15{sel[0]}};
    result = result | ( input_1 & {15{sel[1]}});
    result = result | ( input_2 & {15{sel[2]}});
    MUX1HOT_v_15_3_2 = result;
  end
  endfunction
  function [14:0] MUX1HOT_v_15_6_2;
    input [14:0] input_5;
    input [14:0] input_4;
    input [14:0] input_3;
    input [14:0] input_2;
    input [14:0] input_1;
    input [14:0] input_0;
    input [5:0] sel;
    reg [14:0] result;
  begin
    result = input_0 & {15{sel[0]}};
    result = result | ( input_1 & {15{sel[1]}});
    result = result | ( input_2 & {15{sel[2]}});
    result = result | ( input_3 & {15{sel[3]}});
    result = result | ( input_4 & {15{sel[4]}});
    result = result | ( input_5 & {15{sel[5]}});
    MUX1HOT_v_15_6_2 = result;
  end
  endfunction
  function [14:0] MUX1HOT_v_15_7_2;
    input [14:0] input_6;
    input [14:0] input_5;
    input [14:0] input_4;
    input [14:0] input_3;
    input [14:0] input_2;
    input [14:0] input_1;
    input [14:0] input_0;
    input [6:0] sel;
    reg [14:0] result;
  begin
    result = input_0 & {15{sel[0]}};
    result = result | ( input_1 & {15{sel[1]}});
    result = result | ( input_2 & {15{sel[2]}});
    result = result | ( input_3 & {15{sel[3]}});
    result = result | ( input_4 & {15{sel[4]}});
    result = result | ( input_5 & {15{sel[5]}});
    result = result | ( input_6 & {15{sel[6]}});
    MUX1HOT_v_15_7_2 = result;
  end
  endfunction
  function [15:0] MUX1HOT_v_16_3_2;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [2:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | ( input_1 & {16{sel[1]}});
    result = result | ( input_2 & {16{sel[2]}});
    MUX1HOT_v_16_3_2 = result;
  end
  endfunction
  function [3:0] MUX1HOT_v_4_4_2;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [3:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    result = result | ( input_3 & {4{sel[3]}});
    MUX1HOT_v_4_4_2 = result;
  end
  endfunction
  function [3:0] MUX1HOT_v_4_6_2;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [5:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    result = result | ( input_3 & {4{sel[3]}});
    result = result | ( input_4 & {4{sel[4]}});
    result = result | ( input_5 & {4{sel[5]}});
    MUX1HOT_v_4_6_2 = result;
  end
  endfunction
  function [4:0] MUX1HOT_v_5_3_2;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [2:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | ( input_1 & {5{sel[1]}});
    result = result | ( input_2 & {5{sel[2]}});
    MUX1HOT_v_5_3_2 = result;
  end
  endfunction
  function [6:0] MUX1HOT_v_7_3_2;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [2:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | ( input_1 & {7{sel[1]}});
    result = result | ( input_2 & {7{sel[2]}});
    MUX1HOT_v_7_3_2 = result;
  end
  endfunction
  function [8:0] MUX1HOT_v_9_4_2;
    input [8:0] input_3;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [3:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | ( input_1 & {9{sel[1]}});
    result = result | ( input_2 & {9{sel[2]}});
    result = result | ( input_3 & {9{sel[3]}});
    MUX1HOT_v_9_4_2 = result;
  end
  endfunction
  function [8:0] MUX1HOT_v_9_5_2;
    input [8:0] input_4;
    input [8:0] input_3;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [4:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | ( input_1 & {9{sel[1]}});
    result = result | ( input_2 & {9{sel[2]}});
    result = result | ( input_3 & {9{sel[3]}});
    result = result | ( input_4 & {9{sel[4]}});
    MUX1HOT_v_9_5_2 = result;
  end
  endfunction
  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction
  function [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction
  function [14:0] MUX_v_15_2_2;
    input [14:0] input_0;
    input [14:0] input_1;
    input [0:0] sel;
    reg [14:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_15_2_2 = result;
  end
  endfunction
  function [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction
  function [23:0] MUX_v_24_2_2;
    input [23:0] input_0;
    input [23:0] input_1;
    input [0:0] sel;
    reg [23:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_24_2_2 = result;
  end
  endfunction
  function [48:0] MUX_v_49_2_2;
    input [48:0] input_0;
    input [48:0] input_1;
    input [0:0] sel;
    reg [48:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_49_2_2 = result;
  end
  endfunction
  function [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction
  function [0:0] readslicef_11_1_10;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_11_1_10 = tmp[0:0];
  end
  endfunction
  function [0:0] readslicef_12_1_11;
    input [11:0] vector;
    reg [11:0] tmp;
  begin
    tmp = vector >> 11;
    readslicef_12_1_11 = tmp[0:0];
  end
  endfunction
  function [0:0] readslicef_3_1_2;
    input [2:0] vector;
    reg [2:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_3_1_2 = tmp[0:0];
  end
  endfunction
  function [0:0] readslicef_5_1_4;
    input [4:0] vector;
    reg [4:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_5_1_4 = tmp[0:0];
  end
  endfunction
  function [0:0] readslicef_8_1_7;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_8_1_7 = tmp[0:0];
  end
  endfunction
  function [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction
  function [3:0] signext_4_1;
    input [0:0] vector;
  begin
    signext_4_1= {{3{vector[0]}}, vector};
  end
  endfunction
  function [17:0] conv_s2s_17_18 ;
    input [16:0] vector ;
  begin
    conv_s2s_17_18 = {vector[16], vector};
  end
  endfunction
  function [48:0] conv_s2s_17_49 ;
    input [16:0] vector ;
  begin
    conv_s2s_17_49 = {{32{vector[16]}}, vector};
  end
  endfunction
  function [48:0] conv_s2s_18_49 ;
    input [17:0] vector ;
  begin
    conv_s2s_18_49 = {{31{vector[17]}}, vector};
  end
  endfunction
  function [32:0] conv_s2s_32_33 ;
    input [31:0] vector ;
  begin
    conv_s2s_32_33 = {vector[31], vector};
  end
  endfunction
  function [44:0] conv_s2s_44_45 ;
    input [43:0] vector ;
  begin
    conv_s2s_44_45 = {vector[43], vector};
  end
  endfunction
  function [49:0] conv_s2s_49_50 ;
    input [48:0] vector ;
  begin
    conv_s2s_49_50 = {vector[48], vector};
  end
  endfunction
  function [2:0] conv_s2u_2_3 ;
    input [1:0] vector ;
  begin
    conv_s2u_2_3 = {vector[1], vector};
  end
  endfunction
  function [10:0] conv_s2u_10_11 ;
    input [9:0] vector ;
  begin
    conv_s2u_10_11 = {vector[9], vector};
  end
  endfunction
  function [48:0] conv_s2u_49_49 ;
    input [48:0] vector ;
  begin
    conv_s2u_49_49 = vector;
  end
  endfunction
  function [44:0] conv_u2s_1_45 ;
    input [0:0] vector ;
  begin
    conv_u2s_1_45 = {{44{1'b0}}, vector};
  end
  endfunction
  function [49:0] conv_u2s_1_50 ;
    input [0:0] vector ;
  begin
    conv_u2s_1_50 = {{49{1'b0}}, vector};
  end
  endfunction
  function [8:0] conv_u2s_8_9 ;
    input [7:0] vector ;
  begin
    conv_u2s_8_9 = {1'b0, vector};
  end
  endfunction
  function [9:0] conv_u2u_1_10 ;
    input [0:0] vector ;
  begin
    conv_u2u_1_10 = {{9{1'b0}}, vector};
  end
  endfunction
  function [10:0] conv_u2u_1_11 ;
    input [0:0] vector ;
  begin
    conv_u2u_1_11 = {{10{1'b0}}, vector};
  end
  endfunction
  function [4:0] conv_u2u_4_5 ;
    input [3:0] vector ;
  begin
    conv_u2u_4_5 = {1'b0, vector};
  end
  endfunction
  function [7:0] conv_u2u_7_8 ;
    input [6:0] vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction
  function [16:0] conv_u2u_16_17 ;
    input [15:0] vector ;
  begin
    conv_u2u_16_17 = {1'b0, vector};
  end
  endfunction
endmodule
// ------------------------------------------------------------------
// Design Unit: NV_NVDLA_SDP_CORE_c
// ------------------------------------------------------------------
module NV_NVDLA_SDP_CORE_c (
  nvdla_core_clk, nvdla_core_rstn, chn_in_rsc_z, chn_in_rsc_vz, chn_in_rsc_lz, cfg_offset_rsc_z,
      cfg_scale_rsc_z, cfg_truncate_rsc_z, cfg_proc_precision_rsc_z, cfg_out_precision_rsc_z,
      cfg_mode_eql_rsc_z, chn_out_rsc_z, chn_out_rsc_vz, chn_out_rsc_lz
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [511:0] chn_in_rsc_z;
  input chn_in_rsc_vz;
  output chn_in_rsc_lz;
  input [31:0] cfg_offset_rsc_z;
  input [15:0] cfg_scale_rsc_z;
  input [5:0] cfg_truncate_rsc_z;
  input [1:0] cfg_proc_precision_rsc_z;
  input [1:0] cfg_out_precision_rsc_z;
  input cfg_mode_eql_rsc_z;
  output [271:0] chn_out_rsc_z;
  input chn_out_rsc_vz;
  output chn_out_rsc_lz;
// Interconnect Declarations
  wire chn_in_rsci_oswt;
  wire chn_in_rsci_oswt_unreg;
  wire chn_out_rsci_oswt;
  wire chn_out_rsci_oswt_unreg;
// Interconnect Declarations for Component Instantiations
  SDP_C_chn_in_rsci_unreg chn_in_rsci_unreg_inst (
      .in_0(chn_in_rsci_oswt_unreg),
      .outsig(chn_in_rsci_oswt)
    );
  SDP_C_chn_out_rsci_unreg chn_out_rsci_unreg_inst (
      .in_0(chn_out_rsci_oswt_unreg),
      .outsig(chn_out_rsci_oswt)
    );
  NV_NVDLA_SDP_CORE_c_core NV_NVDLA_SDP_CORE_c_core_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_in_rsc_z(chn_in_rsc_z),
      .chn_in_rsc_vz(chn_in_rsc_vz),
      .chn_in_rsc_lz(chn_in_rsc_lz),
      .cfg_offset_rsc_z(cfg_offset_rsc_z),
      .cfg_scale_rsc_z(cfg_scale_rsc_z),
      .cfg_truncate_rsc_z(cfg_truncate_rsc_z),
      .cfg_proc_precision_rsc_z(cfg_proc_precision_rsc_z),
      .cfg_out_precision_rsc_z(cfg_out_precision_rsc_z),
      .cfg_mode_eql_rsc_z(cfg_mode_eql_rsc_z),
      .chn_out_rsc_z(chn_out_rsc_z),
      .chn_out_rsc_vz(chn_out_rsc_vz),
      .chn_out_rsc_lz(chn_out_rsc_lz),
      .chn_in_rsci_oswt(chn_in_rsci_oswt),
      .chn_in_rsci_oswt_unreg(chn_in_rsci_oswt_unreg),
      .chn_out_rsci_oswt(chn_out_rsci_oswt),
      .chn_out_rsci_oswt_unreg(chn_out_rsci_oswt_unreg)
    );
endmodule
