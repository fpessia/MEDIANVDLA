// ================================================================
// NVDLA Open Source Project
// 
// Copyright(c) 2016 - 2017 NVIDIA Corporation.  Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with 
// this distribution for more information.
// ================================================================

// File Name: HLS_fp17_add.v
`timescale 10ps/1ps
module FP17_ADD_mgc_in_wire_wait_v1 (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  output [width-1:0] d;
  output             lz;
  input              vz;
  input  [width-1:0] z;

  wire               vd;
  wire   [width-1:0] d;
  wire               lz;

  assign d = z;
  assign lz = ld;
  assign vd = vz;

endmodule


//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/FP17_ADD_mgc_out_stdreg_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module FP17_ADD_mgc_out_stdreg_wait_v1 (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  input  [width-1:0] d;
  output             lz;
  input              vz;
  output [width-1:0] z;

  wire               vd;
  wire               lz;
  wire   [width-1:0] z;

  assign z = d;
  assign lz = ld;
  assign vd = vz;

endmodule



//------> ../td_ccore_solutions/leading_sign_23_0_b9d2f049d7a95593b985a5e76dea79445444_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.0/264918 Production Release
//  HLS Date:       Mon Aug  8 13:35:54 PDT 2016
// 
//  Generated by:   ezhang@hk-sim-11-144
//  Generated date: Sun Dec 11 16:48:02 2016
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    FP17_ADD_leading_sign_23_0
// ------------------------------------------------------------------


module FP17_ADD_leading_sign_23_0 (
  mantissa, rtn
);
  input [22:0] mantissa;
  output [4:0] rtn;


  // Interconnect Declarations
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_2;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_2;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_2;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1;
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_9;
  wire c_h_1_10;

  wire[0:0] IntLeadZero_23U_leading_sign_23_0_rtn_and_85_nl;
  wire[0:0] IntLeadZero_23U_leading_sign_23_0_rtn_and_83_nl;
  wire[0:0] IntLeadZero_23U_leading_sign_23_0_rtn_and_90_nl;
  wire[0:0] IntLeadZero_23U_leading_sign_23_0_rtn_IntLeadZero_23U_leading_sign_23_0_rtn_or_2_nl;

  // Interconnect Declarations for Component Instantiations 
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_2 = ~((mantissa[20:19]!=2'b00));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1 = ~((mantissa[22:21]!=2'b00));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1 = ~((mantissa[18:17]!=2'b00));
  assign c_h_1_2 = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1 & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_2;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3 = (mantissa[16:15]==2'b00)
      & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_2 = ~((mantissa[12:11]!=2'b00));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1 = ~((mantissa[14:13]!=2'b00));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1 = ~((mantissa[10:9]!=2'b00));
  assign c_h_1_5 = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1 & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4 = (mantissa[8:7]==2'b00)
      & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1 & c_h_1_5;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_2 = ~((mantissa[4:3]!=2'b00));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1 = ~((mantissa[6:5]!=2'b00));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1 = ~((mantissa[2:1]!=2'b00));
  assign c_h_1_9 = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1 & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_2;
  assign c_h_1_10 = c_h_1_6 & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_and_85_nl = c_h_1_6 & (~ IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4);
  assign IntLeadZero_23U_leading_sign_23_0_rtn_and_83_nl = c_h_1_2 & (c_h_1_5 | (~
      IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3)) & (c_h_1_9 | (~ c_h_1_10));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_and_90_nl = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1
      & (IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1 | (~ IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_2))
      & (~((~(IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1 & (IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1
      | (~ IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_2)))) & c_h_1_6))
      & (~((~(IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1 & (IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1
      | (~ IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_2)))) & c_h_1_10));
  assign IntLeadZero_23U_leading_sign_23_0_rtn_IntLeadZero_23U_leading_sign_23_0_rtn_or_2_nl
      = ((~((mantissa[22]) | (~((mantissa[21:20]!=2'b01))))) & (~(((mantissa[18])
      | (~((mantissa[17:16]!=2'b01)))) & c_h_1_2)) & (~((~((~((mantissa[14]) | (~((mantissa[13:12]!=2'b01)))))
      & (~(((mantissa[10]) | (~((mantissa[9:8]!=2'b01)))) & c_h_1_5)))) & c_h_1_6))
      & (~((~((~((mantissa[6]) | (~((mantissa[5:4]!=2'b01))))) & (~((~((mantissa[2:1]==2'b01)))
      & c_h_1_9)))) & c_h_1_10))) | ((~ (mantissa[0])) & IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1
      & c_h_1_9 & c_h_1_10);
  assign rtn = {c_h_1_10 , (IntLeadZero_23U_leading_sign_23_0_rtn_and_85_nl) , (IntLeadZero_23U_leading_sign_23_0_rtn_and_83_nl)
      , (IntLeadZero_23U_leading_sign_23_0_rtn_and_90_nl) , (IntLeadZero_23U_leading_sign_23_0_rtn_IntLeadZero_23U_leading_sign_23_0_rtn_or_2_nl)};
endmodule




//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/mgc_shift_bl_beh_v4.v 
module FP17_ADD_mgc_shift_bl_v4(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate if ( signd_a )
   begin: SIGNED
     assign z = fshl_s(a,s,a[width_a-1]);
   end
   else
   begin: UNSIGNED
     assign z = fshl_s(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift left - signed shift argument
   function [width_z-1:0] fshl_s;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      reg [width_a:0] sbit_arg1;
      begin
        // Ignoring the possibility that arg2[width_s-1] could be X
        // because of customer complaints regarding X'es in simulation results
        if ( arg2[width_s-1] == 1'b0 )
        begin
          sbit_arg1[width_a:0] = {(width_a+1){1'b0}};
          fshl_s = fshl_u(arg1, arg2, sbit);
        end
        else
        begin
          sbit_arg1[width_a] = sbit;
          sbit_arg1[width_a-1:0] = arg1;
          fshl_s = fshr_u(sbit_arg1[width_a:1], ~arg2, sbit);
        end
      end
   endfunction

endmodule

//------> /home/tools/calypto/catapult-10.0-264918/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v4.v 
module FP17_ADD_mgc_shift_l_v4(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SIGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSIGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.0/264918 Production Release
//  HLS Date:       Mon Aug  8 13:35:54 PDT 2016
// 
//  Generated by:   ezhang@hk-sim-10-184
//  Generated date: Fri Jun 16 21:49:51 2017
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    FP17_ADD_chn_o_rsci_unreg
// ------------------------------------------------------------------


module FP17_ADD_chn_o_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    FP17_ADD_chn_b_rsci_unreg
// ------------------------------------------------------------------


module FP17_ADD_chn_b_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    FP17_ADD_chn_a_rsci_unreg
// ------------------------------------------------------------------


module FP17_ADD_chn_a_rsci_unreg (
  in_0, outsig
);
  input in_0;
  output outsig;



  // Interconnect Declarations for Component Instantiations 
  assign outsig = in_0;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_add_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module HLS_fp17_add_core_core_fsm (
  nvdla_core_clk, nvdla_core_rstn, core_wen, fsm_output
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for HLS_fp17_add_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : HLS_fp17_add_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b1;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_add_core_staller
// ------------------------------------------------------------------


module HLS_fp17_add_core_staller (
  nvdla_core_clk, nvdla_core_rstn, core_wen, chn_a_rsci_wen_comp, core_wten, chn_b_rsci_wen_comp,
      chn_o_rsci_wen_comp
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output core_wen;
  input chn_a_rsci_wen_comp;
  output core_wten;
  reg core_wten;
  input chn_b_rsci_wen_comp;
  input chn_o_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign core_wen = chn_a_rsci_wen_comp & chn_b_rsci_wen_comp & chn_o_rsci_wen_comp;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      core_wten <= 1'b0;
    end
    else begin
      core_wten <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_add_core_chn_o_rsci_chn_o_wait_dp
// ------------------------------------------------------------------


module HLS_fp17_add_core_chn_o_rsci_chn_o_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_o_rsci_oswt, chn_o_rsci_bawt, chn_o_rsci_wen_comp,
      chn_o_rsci_biwt, chn_o_rsci_bdwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_o_rsci_oswt;
  output chn_o_rsci_bawt;
  output chn_o_rsci_wen_comp;
  input chn_o_rsci_biwt;
  input chn_o_rsci_bdwt;


  // Interconnect Declarations
  reg chn_o_rsci_bcwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_o_rsci_bawt = chn_o_rsci_biwt | chn_o_rsci_bcwt;
  assign chn_o_rsci_wen_comp = (~ chn_o_rsci_oswt) | chn_o_rsci_bawt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_bcwt <= 1'b0;
    end
    else begin
      chn_o_rsci_bcwt <= ~((~(chn_o_rsci_bcwt | chn_o_rsci_biwt)) | chn_o_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_add_core_chn_o_rsci_chn_o_wait_ctrl
// ------------------------------------------------------------------


module HLS_fp17_add_core_chn_o_rsci_chn_o_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_o_rsci_oswt, core_wen, core_wten, chn_o_rsci_iswt0,
      chn_o_rsci_ld_core_psct, chn_o_rsci_biwt, chn_o_rsci_bdwt, chn_o_rsci_ld_core_sct,
      chn_o_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_o_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_o_rsci_iswt0;
  input chn_o_rsci_ld_core_psct;
  output chn_o_rsci_biwt;
  output chn_o_rsci_bdwt;
  output chn_o_rsci_ld_core_sct;
  input chn_o_rsci_vd;


  // Interconnect Declarations
  wire chn_o_rsci_ogwt;
  wire chn_o_rsci_pdswt0;
  reg chn_o_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_o_rsci_pdswt0 = (~ core_wten) & chn_o_rsci_iswt0;
  assign chn_o_rsci_biwt = chn_o_rsci_ogwt & chn_o_rsci_vd;
  assign chn_o_rsci_ogwt = chn_o_rsci_pdswt0 | chn_o_rsci_icwt;
  assign chn_o_rsci_bdwt = chn_o_rsci_oswt & core_wen;
  assign chn_o_rsci_ld_core_sct = chn_o_rsci_ld_core_psct & chn_o_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_icwt <= 1'b0;
    end
    else begin
      chn_o_rsci_icwt <= ~((~(chn_o_rsci_icwt | chn_o_rsci_pdswt0)) | chn_o_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_add_core_chn_b_rsci_chn_b_wait_dp
// ------------------------------------------------------------------


module HLS_fp17_add_core_chn_b_rsci_chn_b_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_b_rsci_oswt, chn_b_rsci_bawt, chn_b_rsci_wen_comp,
      chn_b_rsci_d_mxwt, chn_b_rsci_biwt, chn_b_rsci_bdwt, chn_b_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_b_rsci_oswt;
  output chn_b_rsci_bawt;
  output chn_b_rsci_wen_comp;
  output [16:0] chn_b_rsci_d_mxwt;
  input chn_b_rsci_biwt;
  input chn_b_rsci_bdwt;
  input [16:0] chn_b_rsci_d;


  // Interconnect Declarations
  reg chn_b_rsci_bcwt;
  reg [16:0] chn_b_rsci_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_b_rsci_bawt = chn_b_rsci_biwt | chn_b_rsci_bcwt;
  assign chn_b_rsci_wen_comp = (~ chn_b_rsci_oswt) | chn_b_rsci_bawt;
  assign chn_b_rsci_d_mxwt = MUX_v_17_2_2(chn_b_rsci_d, chn_b_rsci_d_bfwt, chn_b_rsci_bcwt);
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_b_rsci_bcwt <= 1'b0;
      chn_b_rsci_d_bfwt <= 17'b0;
    end
    else begin
      chn_b_rsci_bcwt <= ~((~(chn_b_rsci_bcwt | chn_b_rsci_biwt)) | chn_b_rsci_bdwt);
      chn_b_rsci_d_bfwt <= chn_b_rsci_d_mxwt;
    end
  end

  function [16:0] MUX_v_17_2_2;
    input [16:0] input_0;
    input [16:0] input_1;
    input [0:0] sel;
    reg [16:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_17_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_add_core_chn_b_rsci_chn_b_wait_ctrl
// ------------------------------------------------------------------


module HLS_fp17_add_core_chn_b_rsci_chn_b_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_b_rsci_oswt, core_wen, core_wten, chn_b_rsci_iswt0,
      chn_b_rsci_ld_core_psct, chn_b_rsci_biwt, chn_b_rsci_bdwt, chn_b_rsci_ld_core_sct,
      chn_b_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_b_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_b_rsci_iswt0;
  input chn_b_rsci_ld_core_psct;
  output chn_b_rsci_biwt;
  output chn_b_rsci_bdwt;
  output chn_b_rsci_ld_core_sct;
  input chn_b_rsci_vd;


  // Interconnect Declarations
  wire chn_b_rsci_ogwt;
  wire chn_b_rsci_pdswt0;
  reg chn_b_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_b_rsci_pdswt0 = (~ core_wten) & chn_b_rsci_iswt0;
  assign chn_b_rsci_biwt = chn_b_rsci_ogwt & chn_b_rsci_vd;
  assign chn_b_rsci_ogwt = chn_b_rsci_pdswt0 | chn_b_rsci_icwt;
  assign chn_b_rsci_bdwt = chn_b_rsci_oswt & core_wen;
  assign chn_b_rsci_ld_core_sct = chn_b_rsci_ld_core_psct & chn_b_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_b_rsci_icwt <= 1'b0;
    end
    else begin
      chn_b_rsci_icwt <= ~((~(chn_b_rsci_icwt | chn_b_rsci_pdswt0)) | chn_b_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_add_core_chn_a_rsci_chn_a_wait_dp
// ------------------------------------------------------------------


module HLS_fp17_add_core_chn_a_rsci_chn_a_wait_dp (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsci_oswt, chn_a_rsci_bawt, chn_a_rsci_wen_comp,
      chn_a_rsci_d_mxwt, chn_a_rsci_biwt, chn_a_rsci_bdwt, chn_a_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_a_rsci_oswt;
  output chn_a_rsci_bawt;
  output chn_a_rsci_wen_comp;
  output [16:0] chn_a_rsci_d_mxwt;
  input chn_a_rsci_biwt;
  input chn_a_rsci_bdwt;
  input [16:0] chn_a_rsci_d;


  // Interconnect Declarations
  reg chn_a_rsci_bcwt;
  reg [16:0] chn_a_rsci_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_a_rsci_bawt = chn_a_rsci_biwt | chn_a_rsci_bcwt;
  assign chn_a_rsci_wen_comp = (~ chn_a_rsci_oswt) | chn_a_rsci_bawt;
  assign chn_a_rsci_d_mxwt = MUX_v_17_2_2(chn_a_rsci_d, chn_a_rsci_d_bfwt, chn_a_rsci_bcwt);
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_a_rsci_bcwt <= 1'b0;
      chn_a_rsci_d_bfwt <= 17'b0;
    end
    else begin
      chn_a_rsci_bcwt <= ~((~(chn_a_rsci_bcwt | chn_a_rsci_biwt)) | chn_a_rsci_bdwt);
      chn_a_rsci_d_bfwt <= chn_a_rsci_d_mxwt;
    end
  end

  function [16:0] MUX_v_17_2_2;
    input [16:0] input_0;
    input [16:0] input_1;
    input [0:0] sel;
    reg [16:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_17_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_add_core_chn_a_rsci_chn_a_wait_ctrl
// ------------------------------------------------------------------


module HLS_fp17_add_core_chn_a_rsci_chn_a_wait_ctrl (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsci_oswt, core_wen, chn_a_rsci_iswt0, chn_a_rsci_ld_core_psct,
      core_wten, chn_a_rsci_biwt, chn_a_rsci_bdwt, chn_a_rsci_ld_core_sct, chn_a_rsci_vd
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input chn_a_rsci_oswt;
  input core_wen;
  input chn_a_rsci_iswt0;
  input chn_a_rsci_ld_core_psct;
  input core_wten;
  output chn_a_rsci_biwt;
  output chn_a_rsci_bdwt;
  output chn_a_rsci_ld_core_sct;
  input chn_a_rsci_vd;


  // Interconnect Declarations
  wire chn_a_rsci_ogwt;
  wire chn_a_rsci_pdswt0;
  reg chn_a_rsci_icwt;


  // Interconnect Declarations for Component Instantiations 
  assign chn_a_rsci_pdswt0 = (~ core_wten) & chn_a_rsci_iswt0;
  assign chn_a_rsci_biwt = chn_a_rsci_ogwt & chn_a_rsci_vd;
  assign chn_a_rsci_ogwt = chn_a_rsci_pdswt0 | chn_a_rsci_icwt;
  assign chn_a_rsci_bdwt = chn_a_rsci_oswt & core_wen;
  assign chn_a_rsci_ld_core_sct = chn_a_rsci_ld_core_psct & chn_a_rsci_ogwt;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_a_rsci_icwt <= 1'b0;
    end
    else begin
      chn_a_rsci_icwt <= ~((~(chn_a_rsci_icwt | chn_a_rsci_pdswt0)) | chn_a_rsci_biwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_add_core_chn_o_rsci
// ------------------------------------------------------------------


module HLS_fp17_add_core_chn_o_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_o_rsc_z, chn_o_rsc_vz, chn_o_rsc_lz, chn_o_rsci_oswt,
      core_wen, core_wten, chn_o_rsci_iswt0, chn_o_rsci_bawt, chn_o_rsci_wen_comp,
      chn_o_rsci_ld_core_psct, chn_o_rsci_d
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  output [16:0] chn_o_rsc_z;
  input chn_o_rsc_vz;
  output chn_o_rsc_lz;
  input chn_o_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_o_rsci_iswt0;
  output chn_o_rsci_bawt;
  output chn_o_rsci_wen_comp;
  input chn_o_rsci_ld_core_psct;
  input [16:0] chn_o_rsci_d;


  // Interconnect Declarations
  wire chn_o_rsci_biwt;
  wire chn_o_rsci_bdwt;
  wire chn_o_rsci_ld_core_sct;
  wire chn_o_rsci_vd;


  // Interconnect Declarations for Component Instantiations 
  FP17_ADD_mgc_out_stdreg_wait_v1 #(.rscid(32'sd3),
  .width(32'sd17)) chn_o_rsci (
      .ld(chn_o_rsci_ld_core_sct),
      .vd(chn_o_rsci_vd),
      .d(chn_o_rsci_d),
      .lz(chn_o_rsc_lz),
      .vz(chn_o_rsc_vz),
      .z(chn_o_rsc_z)
    );
  HLS_fp17_add_core_chn_o_rsci_chn_o_wait_ctrl HLS_fp17_add_core_chn_o_rsci_chn_o_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_o_rsci_oswt(chn_o_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_o_rsci_iswt0(chn_o_rsci_iswt0),
      .chn_o_rsci_ld_core_psct(chn_o_rsci_ld_core_psct),
      .chn_o_rsci_biwt(chn_o_rsci_biwt),
      .chn_o_rsci_bdwt(chn_o_rsci_bdwt),
      .chn_o_rsci_ld_core_sct(chn_o_rsci_ld_core_sct),
      .chn_o_rsci_vd(chn_o_rsci_vd)
    );
  HLS_fp17_add_core_chn_o_rsci_chn_o_wait_dp HLS_fp17_add_core_chn_o_rsci_chn_o_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_o_rsci_oswt(chn_o_rsci_oswt),
      .chn_o_rsci_bawt(chn_o_rsci_bawt),
      .chn_o_rsci_wen_comp(chn_o_rsci_wen_comp),
      .chn_o_rsci_biwt(chn_o_rsci_biwt),
      .chn_o_rsci_bdwt(chn_o_rsci_bdwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_add_core_chn_b_rsci
// ------------------------------------------------------------------


module HLS_fp17_add_core_chn_b_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_b_rsc_z, chn_b_rsc_vz, chn_b_rsc_lz, chn_b_rsci_oswt,
      core_wen, core_wten, chn_b_rsci_iswt0, chn_b_rsci_bawt, chn_b_rsci_wen_comp,
      chn_b_rsci_ld_core_psct, chn_b_rsci_d_mxwt
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [16:0] chn_b_rsc_z;
  input chn_b_rsc_vz;
  output chn_b_rsc_lz;
  input chn_b_rsci_oswt;
  input core_wen;
  input core_wten;
  input chn_b_rsci_iswt0;
  output chn_b_rsci_bawt;
  output chn_b_rsci_wen_comp;
  input chn_b_rsci_ld_core_psct;
  output [16:0] chn_b_rsci_d_mxwt;


  // Interconnect Declarations
  wire chn_b_rsci_biwt;
  wire chn_b_rsci_bdwt;
  wire chn_b_rsci_ld_core_sct;
  wire chn_b_rsci_vd;
  wire [16:0] chn_b_rsci_d;


  // Interconnect Declarations for Component Instantiations 
  FP17_ADD_mgc_in_wire_wait_v1 #(.rscid(32'sd2),
  .width(32'sd17)) chn_b_rsci (
      .ld(chn_b_rsci_ld_core_sct),
      .vd(chn_b_rsci_vd),
      .d(chn_b_rsci_d),
      .lz(chn_b_rsc_lz),
      .vz(chn_b_rsc_vz),
      .z(chn_b_rsc_z)
    );
  HLS_fp17_add_core_chn_b_rsci_chn_b_wait_ctrl HLS_fp17_add_core_chn_b_rsci_chn_b_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_b_rsci_oswt(chn_b_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_b_rsci_iswt0(chn_b_rsci_iswt0),
      .chn_b_rsci_ld_core_psct(chn_b_rsci_ld_core_psct),
      .chn_b_rsci_biwt(chn_b_rsci_biwt),
      .chn_b_rsci_bdwt(chn_b_rsci_bdwt),
      .chn_b_rsci_ld_core_sct(chn_b_rsci_ld_core_sct),
      .chn_b_rsci_vd(chn_b_rsci_vd)
    );
  HLS_fp17_add_core_chn_b_rsci_chn_b_wait_dp HLS_fp17_add_core_chn_b_rsci_chn_b_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_b_rsci_oswt(chn_b_rsci_oswt),
      .chn_b_rsci_bawt(chn_b_rsci_bawt),
      .chn_b_rsci_wen_comp(chn_b_rsci_wen_comp),
      .chn_b_rsci_d_mxwt(chn_b_rsci_d_mxwt),
      .chn_b_rsci_biwt(chn_b_rsci_biwt),
      .chn_b_rsci_bdwt(chn_b_rsci_bdwt),
      .chn_b_rsci_d(chn_b_rsci_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_add_core_chn_a_rsci
// ------------------------------------------------------------------


module HLS_fp17_add_core_chn_a_rsci (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsc_z, chn_a_rsc_vz, chn_a_rsc_lz, chn_a_rsci_oswt,
      core_wen, chn_a_rsci_iswt0, chn_a_rsci_bawt, chn_a_rsci_wen_comp, chn_a_rsci_ld_core_psct,
      chn_a_rsci_d_mxwt, core_wten
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [16:0] chn_a_rsc_z;
  input chn_a_rsc_vz;
  output chn_a_rsc_lz;
  input chn_a_rsci_oswt;
  input core_wen;
  input chn_a_rsci_iswt0;
  output chn_a_rsci_bawt;
  output chn_a_rsci_wen_comp;
  input chn_a_rsci_ld_core_psct;
  output [16:0] chn_a_rsci_d_mxwt;
  input core_wten;


  // Interconnect Declarations
  wire chn_a_rsci_biwt;
  wire chn_a_rsci_bdwt;
  wire chn_a_rsci_ld_core_sct;
  wire chn_a_rsci_vd;
  wire [16:0] chn_a_rsci_d;


  // Interconnect Declarations for Component Instantiations 
  FP17_ADD_mgc_in_wire_wait_v1 #(.rscid(32'sd1),
  .width(32'sd17)) chn_a_rsci (
      .ld(chn_a_rsci_ld_core_sct),
      .vd(chn_a_rsci_vd),
      .d(chn_a_rsci_d),
      .lz(chn_a_rsc_lz),
      .vz(chn_a_rsc_vz),
      .z(chn_a_rsc_z)
    );
  HLS_fp17_add_core_chn_a_rsci_chn_a_wait_ctrl HLS_fp17_add_core_chn_a_rsci_chn_a_wait_ctrl_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_a_rsci_oswt(chn_a_rsci_oswt),
      .core_wen(core_wen),
      .chn_a_rsci_iswt0(chn_a_rsci_iswt0),
      .chn_a_rsci_ld_core_psct(chn_a_rsci_ld_core_psct),
      .core_wten(core_wten),
      .chn_a_rsci_biwt(chn_a_rsci_biwt),
      .chn_a_rsci_bdwt(chn_a_rsci_bdwt),
      .chn_a_rsci_ld_core_sct(chn_a_rsci_ld_core_sct),
      .chn_a_rsci_vd(chn_a_rsci_vd)
    );
  HLS_fp17_add_core_chn_a_rsci_chn_a_wait_dp HLS_fp17_add_core_chn_a_rsci_chn_a_wait_dp_inst
      (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_a_rsci_oswt(chn_a_rsci_oswt),
      .chn_a_rsci_bawt(chn_a_rsci_bawt),
      .chn_a_rsci_wen_comp(chn_a_rsci_wen_comp),
      .chn_a_rsci_d_mxwt(chn_a_rsci_d_mxwt),
      .chn_a_rsci_biwt(chn_a_rsci_biwt),
      .chn_a_rsci_bdwt(chn_a_rsci_bdwt),
      .chn_a_rsci_d(chn_a_rsci_d)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_add_core
// ------------------------------------------------------------------


module HLS_fp17_add_core (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsc_z, chn_a_rsc_vz, chn_a_rsc_lz, chn_b_rsc_z,
      chn_b_rsc_vz, chn_b_rsc_lz, chn_o_rsc_z, chn_o_rsc_vz, chn_o_rsc_lz, chn_a_rsci_oswt,
      chn_b_rsci_oswt, chn_o_rsci_oswt, chn_o_rsci_oswt_unreg, chn_a_rsci_oswt_unreg_pff
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [16:0] chn_a_rsc_z;
  input chn_a_rsc_vz;
  output chn_a_rsc_lz;
  input [16:0] chn_b_rsc_z;
  input chn_b_rsc_vz;
  output chn_b_rsc_lz;
  output [16:0] chn_o_rsc_z;
  input chn_o_rsc_vz;
  output chn_o_rsc_lz;
  input chn_a_rsci_oswt;
  input chn_b_rsci_oswt;
  input chn_o_rsci_oswt;
  output chn_o_rsci_oswt_unreg;
  output chn_a_rsci_oswt_unreg_pff;


  // Interconnect Declarations
  wire core_wen;
  wire chn_a_rsci_bawt;
  wire chn_a_rsci_wen_comp;
  wire [16:0] chn_a_rsci_d_mxwt;
  wire core_wten;
  wire chn_b_rsci_bawt;
  wire chn_b_rsci_wen_comp;
  wire [16:0] chn_b_rsci_d_mxwt;
  reg chn_o_rsci_iswt0;
  wire chn_o_rsci_bawt;
  wire chn_o_rsci_wen_comp;
  reg chn_o_rsci_d_16;
  reg [5:0] chn_o_rsci_d_15_10;
  reg [9:0] chn_o_rsci_d_9_0;
  wire [1:0] fsm_output;
  wire IsNaN_6U_10U_IsNaN_6U_10U_nor_tmp;
  wire FpAdd_6U_10U_is_a_greater_oif_equal_tmp;
  wire FpMantRNE_23U_11U_else_and_tmp;
  wire IsNaN_6U_10U_1_IsNaN_6U_10U_1_nor_tmp;
  wire nor_tmp_1;
  wire mux_tmp_2;
  wire or_tmp_10;
  wire mux_tmp_6;
  wire mux_tmp_8;
  wire or_tmp_25;
  wire nor_tmp_8;
  wire or_tmp_43;
  wire not_tmp_34;
  wire and_dcpl_7;
  wire and_dcpl_13;
  wire and_dcpl_14;
  wire and_dcpl_15;
  wire and_dcpl_38;
  wire or_tmp_47;
  wire or_tmp_53;
  reg main_stage_v_1;
  reg main_stage_v_2;
  reg main_stage_v_3;
  reg IsNaN_6U_10U_1_land_lpi_1_dfm_4;
  reg IsNaN_6U_10U_1_land_lpi_1_dfm_5;
  reg IsNaN_6U_10U_1_land_lpi_1_dfm_6;
  reg [23:0] FpAdd_6U_10U_int_mant_p1_sva_3;
  reg FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_3;
  reg [5:0] FpAdd_6U_10U_qr_lpi_1_dfm_3;
  reg [5:0] FpAdd_6U_10U_qr_lpi_1_dfm_4;
  reg [5:0] FpAdd_6U_10U_o_expo_lpi_1_dfm_10;
  reg FpAdd_6U_10U_is_inf_lpi_1_dfm_4;
  reg FpMantRNE_23U_11U_else_carry_sva_2;
  reg FpMantRNE_23U_11U_else_and_svs_2;
  reg IsNaN_6U_10U_land_lpi_1_dfm_6;
  reg FpAdd_6U_10U_IsZero_6U_10U_or_itm_2;
  reg [6:0] FpAdd_6U_10U_a_left_shift_acc_itm_2;
  wire [7:0] nl_FpAdd_6U_10U_a_left_shift_acc_itm_2;
  reg FpAdd_6U_10U_IsZero_6U_10U_1_or_itm_2;
  reg [6:0] FpAdd_6U_10U_b_left_shift_acc_itm_2;
  wire [7:0] nl_FpAdd_6U_10U_b_left_shift_acc_itm_2;
  reg [9:0] FpSignedBitsToFloat_6U_10U_1_slc_FpSignedBitsToFloat_6U_10U_1_ubits_9_0_itm_3;
  reg [9:0] FpSignedBitsToFloat_6U_10U_1_slc_FpSignedBitsToFloat_6U_10U_1_ubits_9_0_itm_4;
  reg FpAdd_6U_10U_mux_13_itm_4;
  reg FpAdd_6U_10U_mux_13_itm_5;
  reg FpAdd_6U_10U_mux_13_itm_6;
  reg [5:0] FpSignedBitsToFloat_6U_10U_1_slc_FpSignedBitsToFloat_6U_10U_1_ubits_15_10_itm_3;
  reg [5:0] FpSignedBitsToFloat_6U_10U_1_slc_FpSignedBitsToFloat_6U_10U_1_ubits_15_10_itm_4;
  reg IsNaN_6U_10U_land_lpi_1_dfm_st_4;
  reg IsNaN_6U_10U_land_lpi_1_dfm_st_5;
  reg [15:0] FpSignedBitsToFloat_6U_10U_bits_sva_1_15_0_1;
  reg [15:0] FpSignedBitsToFloat_6U_10U_bits_1_sva_1_15_0_1;
  wire main_stage_en_1;
  wire FpAdd_6U_10U_is_inf_lpi_1_dfm_2_mx0;
  wire FpAdd_6U_10U_FpAdd_6U_10U_nor_2_m1c;
  wire and_58_m1c;
  reg reg_chn_b_rsci_iswt0_cse;
  reg reg_chn_b_rsci_ld_core_psct_cse;
  wire chn_o_and_1_cse;
  wire nor_24_cse;
  wire FpAdd_6U_10U_or_cse;
  wire nor_3_cse;
  reg reg_chn_o_rsci_ld_core_psct_cse;
  wire or_61_cse;
  wire or_5_cse;
  wire nor_7_cse;
  wire and_41_cse;
  wire FpAdd_6U_10U_o_expo_FpAdd_6U_10U_o_expo_nor_rgt;
  wire FpAdd_6U_10U_and_1_rgt;
  wire FpAdd_6U_10U_and_2_rgt;
  wire and_47_rgt;
  wire and_51_rgt;
  wire FpSignedBitsToFloat_6U_10U_or_1_rgt;
  wire [22:0] FpNormalize_6U_23U_else_lshift_itm;
  wire FpAdd_6U_10U_a_right_shift_qelse_and_tmp;
  wire [5:0] z_out;
  wire FpAdd_6U_10U_if_2_and_tmp;
  wire chn_o_rsci_d_9_0_mx0c1;
  wire main_stage_v_1_mx0c1;
  wire main_stage_v_2_mx0c1;
  wire main_stage_v_3_mx0c1;
  wire FpMantRNE_23U_11U_else_carry_sva_mx0w0;
  wire FpAdd_6U_10U_and_tmp;
  wire [22:0] FpAdd_6U_10U_addend_larger_asn_1_mx0w1;
  wire [22:0] FpAdd_6U_10U_addend_larger_qr_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_addend_smaller_qr_lpi_1_dfm_mx0;
  wire [22:0] FpAdd_6U_10U_a_int_mant_p1_sva;
  wire [21:0] FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0;
  wire [22:0] FpAdd_6U_10U_int_mant_1_lpi_1_dfm_1;
  wire FpNormalize_6U_23U_oelse_not_3;
  wire [4:0] libraries_leading_sign_23_0_b9d2f049d7a95593b985a5e76dea79445444_1;
  wire IsNaN_6U_10U_aelse_and_cse;
  wire FpAdd_6U_10U_and_8_cse;
  wire IsNaN_6U_10U_1_aelse_and_cse;
  wire FpSignedBitsToFloat_6U_10U_1_FpSignedBitsToFloat_6U_10U_1_or_1_cse;
  reg reg_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_st_1_cse;
  wire mux_24_cse;
  wire or_75_cse;
  wire nand_cse;
  wire FpAdd_6U_10U_is_a_greater_acc_1_itm_6_1;
  wire FpAdd_6U_10U_if_3_if_acc_1_itm_5_1;
  wire FpAdd_6U_10U_if_4_if_acc_1_itm_5_1;
  wire FpAdd_6U_10U_is_a_greater_oif_aelse_acc_itm_10_1;

  wire[9:0] FpAdd_6U_10U_FpAdd_6U_10U_or_2_nl;
  wire[9:0] FpMantRNE_23U_11U_else_acc_nl;
  wire[10:0] nl_FpMantRNE_23U_11U_else_acc_nl;
  wire[0:0] FpSignedBitsToFloat_6U_10U_1_and_nl;
  wire[5:0] FpAdd_6U_10U_if_4_if_acc_nl;
  wire[6:0] nl_FpAdd_6U_10U_if_4_if_acc_nl;
  wire[0:0] FpAdd_6U_10U_and_nl;
  wire[0:0] FpAdd_6U_10U_and_3_nl;
  wire[0:0] FpAdd_6U_10U_and_7_nl;
  wire[24:0] acc_1_nl;
  wire[25:0] nl_acc_1_nl;
  wire[22:0] FpAdd_6U_10U_else_2_mux_2_nl;
  wire[22:0] FpAdd_6U_10U_else_2_mux_3_nl;
  wire[0:0] mux_3_nl;
  wire[0:0] nor_35_nl;
  wire[0:0] nor_36_nl;
  wire[5:0] FpNormalize_6U_23U_FpNormalize_6U_23U_and_nl;
  wire[5:0] FpNormalize_6U_23U_else_acc_nl;
  wire[7:0] nl_FpNormalize_6U_23U_else_acc_nl;
  wire[5:0] FpAdd_6U_10U_if_3_if_acc_nl;
  wire[6:0] nl_FpAdd_6U_10U_if_3_if_acc_nl;
  wire[0:0] mux_10_nl;
  wire[0:0] mux_9_nl;
  wire[0:0] and_11_nl;
  wire[0:0] or_18_nl;
  wire[0:0] mux_14_nl;
  wire[0:0] mux_12_nl;
  wire[0:0] mux_11_nl;
  wire[0:0] mux_13_nl;
  wire[0:0] nor_25_nl;
  wire[0:0] and_84_nl;
  wire[0:0] mux_16_nl;
  wire[0:0] or_31_nl;
  wire[0:0] mux_15_nl;
  wire[0:0] nor_23_nl;
  wire[0:0] mux_18_nl;
  wire[0:0] or_35_nl;
  wire[0:0] mux_17_nl;
  wire[0:0] nor_22_nl;
  wire[0:0] and_82_nl;
  wire[0:0] or_1_nl;
  wire[0:0] mux_nl;
  wire[0:0] nor_39_nl;
  wire[5:0] FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl;
  wire[5:0] FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl;
  wire[0:0] FpAdd_6U_10U_is_a_greater_oelse_not_5_nl;
  wire[0:0] mux_33_nl;
  wire[0:0] mux_32_nl;
  wire[0:0] mux_31_nl;
  wire[0:0] and_91_nl;
  wire[0:0] mux_35_nl;
  wire[0:0] mux_34_nl;
  wire[0:0] or_44_nl;
  wire[6:0] FpAdd_6U_10U_is_a_greater_acc_1_nl;
  wire[8:0] nl_FpAdd_6U_10U_is_a_greater_acc_1_nl;
  wire[5:0] FpAdd_6U_10U_if_3_if_acc_1_nl;
  wire[6:0] nl_FpAdd_6U_10U_if_3_if_acc_1_nl;
  wire[5:0] FpAdd_6U_10U_if_4_if_acc_1_nl;
  wire[6:0] nl_FpAdd_6U_10U_if_4_if_acc_1_nl;
  wire[0:0] FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_1_nl;
  wire[6:0] FpNormalize_6U_23U_acc_nl;
  wire[8:0] nl_FpNormalize_6U_23U_acc_nl;
  wire[0:0] or_3_nl;
  wire[0:0] nor_38_nl;
  wire[0:0] nor_33_nl;
  wire[0:0] mux_5_nl;
  wire[0:0] nor_34_nl;
  wire[0:0] mux_7_nl;
  wire[0:0] or_13_nl;
  wire[0:0] mux_4_nl;
  wire[0:0] nor_31_nl;
  wire[0:0] nor_32_nl;
  wire[10:0] FpAdd_6U_10U_is_a_greater_oif_aelse_acc_nl;
  wire[12:0] nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_nl;
  wire[6:0] acc_nl;
  wire[7:0] nl_acc_nl;
  wire[5:0] FpAdd_6U_10U_b_right_shift_qif_mux_2_nl;
  wire[5:0] FpAdd_6U_10U_b_right_shift_qif_mux_3_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [22:0] nl_leading_sign_23_0_rg_mantissa;
  assign nl_leading_sign_23_0_rg_mantissa = FpAdd_6U_10U_int_mant_p1_sva_3[22:0];
  wire [10:0] nl_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a;
  assign nl_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a = {FpAdd_6U_10U_IsZero_6U_10U_1_or_itm_2
      , (FpSignedBitsToFloat_6U_10U_bits_1_sva_1_15_0_1[9:0])};
  wire [10:0] nl_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a;
  assign nl_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a = {FpAdd_6U_10U_IsZero_6U_10U_or_itm_2
      , (FpSignedBitsToFloat_6U_10U_bits_sva_1_15_0_1[9:0])};
  wire [22:0] nl_FpNormalize_6U_23U_else_lshift_rg_a;
  assign nl_FpNormalize_6U_23U_else_lshift_rg_a = FpAdd_6U_10U_int_mant_p1_sva_3[22:0];
  wire [16:0] nl_HLS_fp17_add_core_chn_o_rsci_inst_chn_o_rsci_d;
  assign nl_HLS_fp17_add_core_chn_o_rsci_inst_chn_o_rsci_d = {chn_o_rsci_d_16 , chn_o_rsci_d_15_10
      , chn_o_rsci_d_9_0};
  FP17_ADD_leading_sign_23_0  leading_sign_23_0_rg (
      .mantissa(nl_leading_sign_23_0_rg_mantissa[22:0]),
      .rtn(libraries_leading_sign_23_0_b9d2f049d7a95593b985a5e76dea79445444_1)
    );
  FP17_ADD_mgc_shift_bl_v4 #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) FpAdd_6U_10U_b_int_mant_p1_lshift_rg (
      .a(nl_FpAdd_6U_10U_b_int_mant_p1_lshift_rg_a[10:0]),
      .s(FpAdd_6U_10U_b_left_shift_acc_itm_2),
      .z(FpAdd_6U_10U_addend_larger_asn_1_mx0w1)
    );
  FP17_ADD_mgc_shift_bl_v4 #(.width_a(32'sd11),
  .signd_a(32'sd0),
  .width_s(32'sd7),
  .width_z(32'sd23)) FpAdd_6U_10U_a_int_mant_p1_lshift_rg (
      .a(nl_FpAdd_6U_10U_a_int_mant_p1_lshift_rg_a[10:0]),
      .s(FpAdd_6U_10U_a_left_shift_acc_itm_2),
      .z(FpAdd_6U_10U_a_int_mant_p1_sva)
    );
  FP17_ADD_mgc_shift_l_v4 #(.width_a(32'sd23),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd23)) FpNormalize_6U_23U_else_lshift_rg (
      .a(nl_FpNormalize_6U_23U_else_lshift_rg_a[22:0]),
      .s(libraries_leading_sign_23_0_b9d2f049d7a95593b985a5e76dea79445444_1),
      .z(FpNormalize_6U_23U_else_lshift_itm)
    );
  HLS_fp17_add_core_chn_a_rsci HLS_fp17_add_core_chn_a_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_a_rsc_z(chn_a_rsc_z),
      .chn_a_rsc_vz(chn_a_rsc_vz),
      .chn_a_rsc_lz(chn_a_rsc_lz),
      .chn_a_rsci_oswt(chn_a_rsci_oswt),
      .core_wen(core_wen),
      .chn_a_rsci_iswt0(reg_chn_b_rsci_iswt0_cse),
      .chn_a_rsci_bawt(chn_a_rsci_bawt),
      .chn_a_rsci_wen_comp(chn_a_rsci_wen_comp),
      .chn_a_rsci_ld_core_psct(reg_chn_b_rsci_ld_core_psct_cse),
      .chn_a_rsci_d_mxwt(chn_a_rsci_d_mxwt),
      .core_wten(core_wten)
    );
  HLS_fp17_add_core_chn_b_rsci HLS_fp17_add_core_chn_b_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_b_rsc_z(chn_b_rsc_z),
      .chn_b_rsc_vz(chn_b_rsc_vz),
      .chn_b_rsc_lz(chn_b_rsc_lz),
      .chn_b_rsci_oswt(chn_b_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_b_rsci_iswt0(reg_chn_b_rsci_iswt0_cse),
      .chn_b_rsci_bawt(chn_b_rsci_bawt),
      .chn_b_rsci_wen_comp(chn_b_rsci_wen_comp),
      .chn_b_rsci_ld_core_psct(reg_chn_b_rsci_ld_core_psct_cse),
      .chn_b_rsci_d_mxwt(chn_b_rsci_d_mxwt)
    );
  HLS_fp17_add_core_chn_o_rsci HLS_fp17_add_core_chn_o_rsci_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_o_rsc_z(chn_o_rsc_z),
      .chn_o_rsc_vz(chn_o_rsc_vz),
      .chn_o_rsc_lz(chn_o_rsc_lz),
      .chn_o_rsci_oswt(chn_o_rsci_oswt),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .chn_o_rsci_iswt0(chn_o_rsci_iswt0),
      .chn_o_rsci_bawt(chn_o_rsci_bawt),
      .chn_o_rsci_wen_comp(chn_o_rsci_wen_comp),
      .chn_o_rsci_ld_core_psct(reg_chn_o_rsci_ld_core_psct_cse),
      .chn_o_rsci_d(nl_HLS_fp17_add_core_chn_o_rsci_inst_chn_o_rsci_d[16:0])
    );
  HLS_fp17_add_core_staller HLS_fp17_add_core_staller_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .chn_a_rsci_wen_comp(chn_a_rsci_wen_comp),
      .core_wten(core_wten),
      .chn_b_rsci_wen_comp(chn_b_rsci_wen_comp),
      .chn_o_rsci_wen_comp(chn_o_rsci_wen_comp)
    );
  HLS_fp17_add_core_core_fsm HLS_fp17_add_core_core_fsm_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign chn_o_and_1_cse = core_wen & (~(and_dcpl_7 | (~ main_stage_v_3)));
  assign FpAdd_6U_10U_or_cse = IsNaN_6U_10U_1_land_lpi_1_dfm_6 | IsNaN_6U_10U_land_lpi_1_dfm_6;
  assign IsNaN_6U_10U_aelse_and_cse = core_wen & (~ and_dcpl_7) & mux_24_cse;
  assign FpAdd_6U_10U_and_8_cse = core_wen & (~ and_dcpl_7) & mux_tmp_2;
  assign and_41_cse = or_5_cse & main_stage_v_2;
  assign nor_3_cse = ~(FpAdd_6U_10U_if_3_if_acc_1_itm_5_1 | (~ (FpAdd_6U_10U_int_mant_p1_sva_3[23])));
  assign or_5_cse = (~ reg_chn_o_rsci_ld_core_psct_cse) | chn_o_rsci_bawt;
  assign FpAdd_6U_10U_o_expo_FpAdd_6U_10U_o_expo_nor_rgt = ~((FpAdd_6U_10U_int_mant_p1_sva_3[23])
      | and_dcpl_7);
  assign FpAdd_6U_10U_and_1_rgt = (~ FpAdd_6U_10U_if_3_if_acc_1_itm_5_1) & (FpAdd_6U_10U_int_mant_p1_sva_3[23])
      & (~ and_dcpl_7);
  assign FpAdd_6U_10U_and_2_rgt = FpAdd_6U_10U_if_3_if_acc_1_itm_5_1 & (FpAdd_6U_10U_int_mant_p1_sva_3[23])
      & (~ and_dcpl_7);
  assign nor_24_cse = ~(FpAdd_6U_10U_if_3_if_acc_1_itm_5_1 | (~ (FpAdd_6U_10U_int_mant_p1_sva_3[23]))
      | IsNaN_6U_10U_1_land_lpi_1_dfm_5);
  assign and_47_rgt = (~(IsNaN_6U_10U_land_lpi_1_dfm_st_5 | IsNaN_6U_10U_1_land_lpi_1_dfm_5))
      & or_5_cse;
  assign or_31_nl = nor_7_cse | main_stage_v_2;
  assign nor_23_nl = ~(reg_chn_o_rsci_ld_core_psct_cse | (~ main_stage_v_2));
  assign mux_15_nl = MUX_s_1_2_2((nor_23_nl), main_stage_v_2, chn_o_rsci_bawt);
  assign mux_16_nl = MUX_s_1_2_2((mux_15_nl), (or_31_nl), main_stage_v_3);
  assign IsNaN_6U_10U_1_aelse_and_cse = core_wen & (~ and_dcpl_7) & (mux_16_nl);
  assign nor_7_cse = ~(chn_o_rsci_bawt | (~ reg_chn_o_rsci_ld_core_psct_cse));
  assign or_61_cse = (FpAdd_6U_10U_is_a_greater_oif_equal_tmp & (~ FpAdd_6U_10U_is_a_greater_oif_aelse_acc_itm_10_1))
      | FpAdd_6U_10U_is_a_greater_acc_1_itm_6_1;
  assign and_51_rgt = or_5_cse & (~ FpAdd_6U_10U_is_a_greater_acc_1_itm_6_1) & ((~
      FpAdd_6U_10U_is_a_greater_oif_equal_tmp) | FpAdd_6U_10U_is_a_greater_oif_aelse_acc_itm_10_1);
  assign or_1_nl = nor_7_cse | nor_tmp_1;
  assign nor_39_nl = ~(reg_chn_o_rsci_ld_core_psct_cse | (~ nor_tmp_1));
  assign mux_nl = MUX_s_1_2_2((nor_39_nl), nor_tmp_1, chn_o_rsci_bawt);
  assign mux_24_cse = MUX_s_1_2_2((mux_nl), (or_1_nl), main_stage_v_1);
  assign FpSignedBitsToFloat_6U_10U_1_FpSignedBitsToFloat_6U_10U_1_or_1_cse = (or_5_cse
      & (~ IsNaN_6U_10U_land_lpi_1_dfm_st_4)) | and_dcpl_38;
  assign or_75_cse = chn_o_rsci_bawt | (~ reg_chn_o_rsci_ld_core_psct_cse) | nor_tmp_8;
  assign and_58_m1c = or_5_cse & (~(IsNaN_6U_10U_IsNaN_6U_10U_nor_tmp | IsNaN_6U_10U_1_IsNaN_6U_10U_1_nor_tmp));
  assign FpSignedBitsToFloat_6U_10U_or_1_rgt = (or_5_cse & (~ IsNaN_6U_10U_IsNaN_6U_10U_nor_tmp)
      & IsNaN_6U_10U_1_IsNaN_6U_10U_1_nor_tmp) | ((~ or_61_cse) & and_58_m1c);
  assign FpAdd_6U_10U_is_a_greater_oif_equal_tmp = (chn_a_rsci_d_mxwt[15:10]) ==
      (chn_b_rsci_d_mxwt[15:10]);
  assign IsNaN_6U_10U_IsNaN_6U_10U_nor_tmp = ~((~((chn_a_rsci_d_mxwt[9:0]!=10'b0000000000)))
      | (chn_a_rsci_d_mxwt[15:10]!=6'b111111));
  assign FpMantRNE_23U_11U_else_carry_sva_mx0w0 = (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[11])
      & ((FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[0]) | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[1])
      | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[2]) | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[3])
      | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[4]) | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[5])
      | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[6]) | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[7])
      | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[8]) | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[9])
      | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[10]) | (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[12]));
  assign FpMantRNE_23U_11U_else_and_tmp = FpMantRNE_23U_11U_else_carry_sva_mx0w0
      & (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[21:12]==10'b1111111111) & ((FpAdd_6U_10U_int_mant_1_lpi_1_dfm_1[22])
      | (FpAdd_6U_10U_int_mant_p1_sva_3[23]));
  assign IsNaN_6U_10U_1_IsNaN_6U_10U_1_nor_tmp = ~((~((chn_b_rsci_d_mxwt[9:0]!=10'b0000000000)))
      | (chn_b_rsci_d_mxwt[15:10]!=6'b111111));
  assign nl_FpAdd_6U_10U_is_a_greater_acc_1_nl = ({1'b1 , (chn_b_rsci_d_mxwt[15:10])})
      + conv_u2u_6_7(~ (chn_a_rsci_d_mxwt[15:10])) + 7'b1;
  assign FpAdd_6U_10U_is_a_greater_acc_1_nl = nl_FpAdd_6U_10U_is_a_greater_acc_1_nl[6:0];
  assign FpAdd_6U_10U_is_a_greater_acc_1_itm_6_1 = readslicef_7_1_6((FpAdd_6U_10U_is_a_greater_acc_1_nl));
  assign nl_FpAdd_6U_10U_if_3_if_acc_1_nl = ({1'b1 , (FpAdd_6U_10U_qr_lpi_1_dfm_4[5:1])})
      + 6'b1;
  assign FpAdd_6U_10U_if_3_if_acc_1_nl = nl_FpAdd_6U_10U_if_3_if_acc_1_nl[5:0];
  assign FpAdd_6U_10U_if_3_if_acc_1_itm_5_1 = readslicef_6_1_5((FpAdd_6U_10U_if_3_if_acc_1_nl));
  assign nl_FpAdd_6U_10U_if_4_if_acc_1_nl = ({1'b1 , (FpAdd_6U_10U_o_expo_lpi_1_dfm_10[5:1])})
      + 6'b1;
  assign FpAdd_6U_10U_if_4_if_acc_1_nl = nl_FpAdd_6U_10U_if_4_if_acc_1_nl[5:0];
  assign FpAdd_6U_10U_if_4_if_acc_1_itm_5_1 = readslicef_6_1_5((FpAdd_6U_10U_if_4_if_acc_1_nl));
  assign FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_1_nl = FpAdd_6U_10U_is_inf_lpi_1_dfm_4
      | (~ FpAdd_6U_10U_if_4_if_acc_1_itm_5_1);
  assign FpAdd_6U_10U_is_inf_lpi_1_dfm_2_mx0 = MUX_s_1_2_2(FpAdd_6U_10U_is_inf_lpi_1_dfm_4,
      (FpAdd_6U_10U_if_4_FpAdd_6U_10U_if_4_or_1_nl), FpMantRNE_23U_11U_else_and_svs_2);
  assign FpAdd_6U_10U_and_tmp = FpAdd_6U_10U_if_4_if_acc_1_itm_5_1 & FpMantRNE_23U_11U_else_and_svs_2;
  assign FpAdd_6U_10U_FpAdd_6U_10U_nor_2_m1c = ~(IsNaN_6U_10U_1_land_lpi_1_dfm_6
      | IsNaN_6U_10U_land_lpi_1_dfm_6);
  assign main_stage_en_1 = chn_a_rsci_bawt & chn_b_rsci_bawt & or_5_cse;
  assign FpAdd_6U_10U_addend_larger_qr_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_addend_larger_asn_1_mx0w1,
      FpAdd_6U_10U_a_int_mant_p1_sva, FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_3);
  assign FpAdd_6U_10U_addend_smaller_qr_lpi_1_dfm_mx0 = MUX_v_23_2_2(FpAdd_6U_10U_a_int_mant_p1_sva,
      FpAdd_6U_10U_addend_larger_asn_1_mx0w1, FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_3);
  assign FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0 = MUX_v_22_2_2((FpAdd_6U_10U_int_mant_1_lpi_1_dfm_1[21:0]),
      (FpAdd_6U_10U_int_mant_p1_sva_3[22:1]), FpAdd_6U_10U_int_mant_p1_sva_3[23]);
  assign FpAdd_6U_10U_int_mant_1_lpi_1_dfm_1 = MUX_v_23_2_2(23'b00000000000000000000000,
      FpNormalize_6U_23U_else_lshift_itm, FpNormalize_6U_23U_oelse_not_3);
  assign nl_FpNormalize_6U_23U_acc_nl = ({1'b1 , (~ FpAdd_6U_10U_qr_lpi_1_dfm_4)})
      + conv_u2s_5_7(libraries_leading_sign_23_0_b9d2f049d7a95593b985a5e76dea79445444_1)
      + 7'b1;
  assign FpNormalize_6U_23U_acc_nl = nl_FpNormalize_6U_23U_acc_nl[6:0];
  assign FpNormalize_6U_23U_oelse_not_3 = ((FpAdd_6U_10U_int_mant_p1_sva_3[22:0]!=23'b00000000000000000000000))
      & (readslicef_7_1_6((FpNormalize_6U_23U_acc_nl)));
  assign nor_tmp_1 = chn_a_rsci_bawt & chn_b_rsci_bawt;
  assign or_3_nl = chn_o_rsci_bawt | (~ reg_chn_o_rsci_ld_core_psct_cse) | main_stage_v_2;
  assign nor_38_nl = ~(chn_o_rsci_bawt | (~(reg_chn_o_rsci_ld_core_psct_cse & main_stage_v_2)));
  assign mux_tmp_2 = MUX_s_1_2_2((nor_38_nl), (or_3_nl), main_stage_v_1);
  assign or_tmp_10 = IsNaN_6U_10U_land_lpi_1_dfm_st_5 | IsNaN_6U_10U_1_land_lpi_1_dfm_5;
  assign nor_34_nl = ~((FpAdd_6U_10U_int_mant_p1_sva_3[23]) | (~ or_5_cse));
  assign mux_5_nl = MUX_s_1_2_2((nor_34_nl), or_5_cse, FpAdd_6U_10U_if_3_if_acc_1_itm_5_1);
  assign nor_33_nl = ~(or_tmp_10 | (~ (mux_5_nl)));
  assign mux_tmp_6 = MUX_s_1_2_2((nor_33_nl), or_5_cse, FpMantRNE_23U_11U_else_and_tmp);
  assign nor_31_nl = ~(FpAdd_6U_10U_if_3_if_acc_1_itm_5_1 | (~((FpAdd_6U_10U_int_mant_p1_sva_3[23])
      & or_5_cse)));
  assign mux_4_nl = MUX_s_1_2_2((nor_31_nl), or_5_cse, or_tmp_10);
  assign or_13_nl = FpMantRNE_23U_11U_else_and_tmp | (~ (mux_4_nl));
  assign mux_7_nl = MUX_s_1_2_2(mux_tmp_6, (or_13_nl), main_stage_v_3);
  assign nor_32_nl = ~((~ main_stage_v_3) | (~ reg_chn_o_rsci_ld_core_psct_cse) |
      chn_o_rsci_bawt);
  assign mux_tmp_8 = MUX_s_1_2_2((nor_32_nl), (mux_7_nl), main_stage_v_2);
  assign or_tmp_25 = main_stage_v_2 | (~ or_5_cse);
  assign nor_tmp_8 = or_tmp_10 & main_stage_v_2;
  assign nand_cse = ~(reg_chn_o_rsci_ld_core_psct_cse & nor_tmp_8);
  assign or_tmp_43 = chn_o_rsci_bawt | nand_cse;
  assign not_tmp_34 = ~(chn_o_rsci_bawt | nand_cse);
  assign and_dcpl_7 = reg_chn_o_rsci_ld_core_psct_cse & (~ chn_o_rsci_bawt);
  assign and_dcpl_13 = or_5_cse & main_stage_v_3;
  assign and_dcpl_14 = reg_chn_o_rsci_ld_core_psct_cse & chn_o_rsci_bawt;
  assign and_dcpl_15 = and_dcpl_14 & (~ main_stage_v_3);
  assign and_dcpl_38 = or_5_cse & IsNaN_6U_10U_land_lpi_1_dfm_st_4;
  assign or_tmp_47 = main_stage_en_1 | (fsm_output[0]);
  assign or_tmp_53 = chn_b_rsci_bawt & chn_a_rsci_bawt & or_5_cse & (fsm_output[1]);
  assign chn_o_rsci_d_9_0_mx0c1 = or_5_cse & main_stage_v_3 & (~ IsNaN_6U_10U_land_lpi_1_dfm_6);
  assign main_stage_v_1_mx0c1 = (~(chn_b_rsci_bawt & chn_a_rsci_bawt)) & or_5_cse
      & main_stage_v_1;
  assign main_stage_v_2_mx0c1 = or_5_cse & main_stage_v_2 & (~ main_stage_v_1);
  assign main_stage_v_3_mx0c1 = or_5_cse & (~ main_stage_v_2) & main_stage_v_3;
  assign nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_nl = ({1'b1 , (chn_a_rsci_d_mxwt[9:0])})
      + conv_u2u_10_11(~ (chn_b_rsci_d_mxwt[9:0])) + 11'b1;
  assign FpAdd_6U_10U_is_a_greater_oif_aelse_acc_nl = nl_FpAdd_6U_10U_is_a_greater_oif_aelse_acc_nl[10:0];
  assign FpAdd_6U_10U_is_a_greater_oif_aelse_acc_itm_10_1 = readslicef_11_1_10((FpAdd_6U_10U_is_a_greater_oif_aelse_acc_nl));
  assign chn_a_rsci_oswt_unreg_pff = or_tmp_53;
  assign chn_o_rsci_oswt_unreg = and_dcpl_14;
  assign FpAdd_6U_10U_a_right_shift_qelse_and_tmp = (fsm_output[1]) & (~((~(FpAdd_6U_10U_is_a_greater_oif_aelse_acc_itm_10_1
      | (~ FpAdd_6U_10U_is_a_greater_oif_equal_tmp))) | FpAdd_6U_10U_is_a_greater_acc_1_itm_6_1));
  assign FpAdd_6U_10U_if_2_and_tmp = (fsm_output[1]) & reg_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_st_1_cse;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_b_rsci_iswt0_cse <= 1'b0;
      chn_o_rsci_iswt0 <= 1'b0;
    end
    else if ( core_wen ) begin
      reg_chn_b_rsci_iswt0_cse <= ~((~ main_stage_en_1) & (fsm_output[1]));
      chn_o_rsci_iswt0 <= and_dcpl_13;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_b_rsci_ld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & or_tmp_47 ) begin
      reg_chn_b_rsci_ld_core_psct_cse <= or_tmp_47;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_d_9_0 <= 10'b0;
    end
    else if ( core_wen & ((or_5_cse & main_stage_v_3 & IsNaN_6U_10U_land_lpi_1_dfm_6)
        | chn_o_rsci_d_9_0_mx0c1) ) begin
      chn_o_rsci_d_9_0 <= MUX_v_10_2_2(FpSignedBitsToFloat_6U_10U_1_slc_FpSignedBitsToFloat_6U_10U_1_ubits_9_0_itm_4,
          (FpAdd_6U_10U_FpAdd_6U_10U_or_2_nl), FpSignedBitsToFloat_6U_10U_1_and_nl);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      chn_o_rsci_d_15_10 <= 6'b0;
      chn_o_rsci_d_16 <= 1'b0;
    end
    else if ( chn_o_and_1_cse ) begin
      chn_o_rsci_d_15_10 <= MUX1HOT_v_6_4_2(FpAdd_6U_10U_o_expo_lpi_1_dfm_10, (FpAdd_6U_10U_if_4_if_acc_nl),
          6'b111110, FpSignedBitsToFloat_6U_10U_1_slc_FpSignedBitsToFloat_6U_10U_1_ubits_15_10_itm_4,
          {(FpAdd_6U_10U_and_nl) , (FpAdd_6U_10U_and_3_nl) , (FpAdd_6U_10U_and_7_nl)
          , FpAdd_6U_10U_or_cse});
      chn_o_rsci_d_16 <= FpAdd_6U_10U_mux_13_itm_6;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      reg_chn_o_rsci_ld_core_psct_cse <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_13 | and_dcpl_15) ) begin
      reg_chn_o_rsci_ld_core_psct_cse <= ~ and_dcpl_15;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_1 <= 1'b0;
    end
    else if ( core_wen & (or_tmp_53 | main_stage_v_1_mx0c1) ) begin
      main_stage_v_1 <= ~ main_stage_v_1_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_land_lpi_1_dfm_st_4 <= 1'b0;
      reg_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_st_1_cse <=
          1'b0;
      FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_3 <= 1'b0;
      FpAdd_6U_10U_IsZero_6U_10U_1_or_itm_2 <= 1'b0;
      FpSignedBitsToFloat_6U_10U_bits_1_sva_1_15_0_1 <= 16'b0;
      FpAdd_6U_10U_b_left_shift_acc_itm_2 <= 7'b0;
      FpAdd_6U_10U_IsZero_6U_10U_or_itm_2 <= 1'b0;
      FpSignedBitsToFloat_6U_10U_bits_sva_1_15_0_1 <= 16'b0;
      FpAdd_6U_10U_a_left_shift_acc_itm_2 <= 7'b0;
      IsNaN_6U_10U_1_land_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_aelse_and_cse ) begin
      IsNaN_6U_10U_land_lpi_1_dfm_st_4 <= IsNaN_6U_10U_IsNaN_6U_10U_nor_tmp;
      reg_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_st_1_cse <=
          ~((chn_a_rsci_d_mxwt[16]) ^ (chn_b_rsci_d_mxwt[16]));
      FpAdd_6U_10U_is_a_greater_lor_lpi_1_dfm_3 <= or_61_cse;
      FpAdd_6U_10U_IsZero_6U_10U_1_or_itm_2 <= (chn_b_rsci_d_mxwt[15:0]!=16'b0000000000000000);
      FpSignedBitsToFloat_6U_10U_bits_1_sva_1_15_0_1 <= chn_b_rsci_d_mxwt[15:0];
      FpAdd_6U_10U_b_left_shift_acc_itm_2 <= nl_FpAdd_6U_10U_b_left_shift_acc_itm_2[6:0];
      FpAdd_6U_10U_IsZero_6U_10U_or_itm_2 <= (chn_a_rsci_d_mxwt[15:0]!=16'b0000000000000000);
      FpSignedBitsToFloat_6U_10U_bits_sva_1_15_0_1 <= chn_a_rsci_d_mxwt[15:0];
      FpAdd_6U_10U_a_left_shift_acc_itm_2 <= nl_FpAdd_6U_10U_a_left_shift_acc_itm_2[6:0];
      IsNaN_6U_10U_1_land_lpi_1_dfm_4 <= IsNaN_6U_10U_1_IsNaN_6U_10U_1_nor_tmp;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_2 <= 1'b0;
    end
    else if ( core_wen & ((or_5_cse & main_stage_v_1) | main_stage_v_2_mx0c1) ) begin
      main_stage_v_2 <= ~ main_stage_v_2_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_qr_lpi_1_dfm_4 <= 6'b0;
      IsNaN_6U_10U_land_lpi_1_dfm_st_5 <= 1'b0;
      IsNaN_6U_10U_1_land_lpi_1_dfm_5 <= 1'b0;
      FpAdd_6U_10U_mux_13_itm_5 <= 1'b0;
    end
    else if ( FpAdd_6U_10U_and_8_cse ) begin
      FpAdd_6U_10U_qr_lpi_1_dfm_4 <= FpAdd_6U_10U_qr_lpi_1_dfm_3;
      IsNaN_6U_10U_land_lpi_1_dfm_st_5 <= IsNaN_6U_10U_land_lpi_1_dfm_st_4;
      IsNaN_6U_10U_1_land_lpi_1_dfm_5 <= IsNaN_6U_10U_1_land_lpi_1_dfm_4;
      FpAdd_6U_10U_mux_13_itm_5 <= FpAdd_6U_10U_mux_13_itm_4;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_int_mant_p1_sva_3 <= 24'b0;
    end
    else if ( core_wen & (~((~(or_5_cse & (~ reg_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_st_1_cse)))
        & (~(or_5_cse & reg_FpAdd_6U_10U_is_addition_FpAdd_6U_10U_is_addition_xnor_svs_st_1_cse))))
        & mux_tmp_2 ) begin
      FpAdd_6U_10U_int_mant_p1_sva_3 <= readslicef_25_24_1((acc_1_nl));
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      main_stage_v_3 <= 1'b0;
    end
    else if ( core_wen & (and_41_cse | main_stage_v_3_mx0c1) ) begin
      main_stage_v_3 <= ~ main_stage_v_3_mx0c1;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpMantRNE_23U_11U_else_carry_sva_2 <= 1'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_3_nl) ) begin
      FpMantRNE_23U_11U_else_carry_sva_2 <= FpMantRNE_23U_11U_else_carry_sva_mx0w0;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_o_expo_lpi_1_dfm_10 <= 6'b0;
    end
    else if ( core_wen & (FpAdd_6U_10U_o_expo_FpAdd_6U_10U_o_expo_nor_rgt | FpAdd_6U_10U_and_1_rgt
        | FpAdd_6U_10U_and_2_rgt) & (mux_10_nl) ) begin
      FpAdd_6U_10U_o_expo_lpi_1_dfm_10 <= MUX1HOT_v_6_3_2((FpNormalize_6U_23U_FpNormalize_6U_23U_and_nl),
          FpAdd_6U_10U_qr_lpi_1_dfm_4, (FpAdd_6U_10U_if_3_if_acc_nl), {FpAdd_6U_10U_o_expo_FpAdd_6U_10U_o_expo_nor_rgt
          , FpAdd_6U_10U_and_1_rgt , FpAdd_6U_10U_and_2_rgt});
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpSignedBitsToFloat_6U_10U_1_slc_FpSignedBitsToFloat_6U_10U_1_ubits_9_0_itm_4
          <= 10'b0;
    end
    else if ( core_wen & ((or_tmp_10 & or_5_cse) | and_47_rgt) & (mux_14_nl) ) begin
      FpSignedBitsToFloat_6U_10U_1_slc_FpSignedBitsToFloat_6U_10U_1_ubits_9_0_itm_4
          <= MUX_v_10_2_2(FpSignedBitsToFloat_6U_10U_1_slc_FpSignedBitsToFloat_6U_10U_1_ubits_9_0_itm_3,
          (FpAdd_6U_10U_int_mant_1_lpi_1_dfm_2_21_0_mx0[21:12]), and_47_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      IsNaN_6U_10U_1_land_lpi_1_dfm_6 <= 1'b0;
      FpAdd_6U_10U_mux_13_itm_6 <= 1'b0;
      IsNaN_6U_10U_land_lpi_1_dfm_6 <= 1'b0;
      FpMantRNE_23U_11U_else_and_svs_2 <= 1'b0;
      FpAdd_6U_10U_is_inf_lpi_1_dfm_4 <= 1'b0;
    end
    else if ( IsNaN_6U_10U_1_aelse_and_cse ) begin
      IsNaN_6U_10U_1_land_lpi_1_dfm_6 <= IsNaN_6U_10U_1_land_lpi_1_dfm_5;
      FpAdd_6U_10U_mux_13_itm_6 <= FpAdd_6U_10U_mux_13_itm_5;
      IsNaN_6U_10U_land_lpi_1_dfm_6 <= IsNaN_6U_10U_land_lpi_1_dfm_st_5;
      FpMantRNE_23U_11U_else_and_svs_2 <= FpMantRNE_23U_11U_else_and_tmp;
      FpAdd_6U_10U_is_inf_lpi_1_dfm_4 <= nor_3_cse;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpSignedBitsToFloat_6U_10U_1_slc_FpSignedBitsToFloat_6U_10U_1_ubits_15_10_itm_4
          <= 6'b0;
    end
    else if ( core_wen & (~ and_dcpl_7) & (mux_18_nl) ) begin
      FpSignedBitsToFloat_6U_10U_1_slc_FpSignedBitsToFloat_6U_10U_1_ubits_15_10_itm_4
          <= FpSignedBitsToFloat_6U_10U_1_slc_FpSignedBitsToFloat_6U_10U_1_ubits_15_10_itm_3;
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_qr_lpi_1_dfm_3 <= 6'b0;
    end
    else if ( core_wen & ((or_61_cse & or_5_cse) | and_51_rgt) & mux_24_cse ) begin
      FpAdd_6U_10U_qr_lpi_1_dfm_3 <= MUX_v_6_2_2((chn_a_rsci_d_mxwt[15:10]), (chn_b_rsci_d_mxwt[15:10]),
          and_51_rgt);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpSignedBitsToFloat_6U_10U_1_slc_FpSignedBitsToFloat_6U_10U_1_ubits_9_0_itm_3
          <= 10'b0;
    end
    else if ( core_wen & FpSignedBitsToFloat_6U_10U_1_FpSignedBitsToFloat_6U_10U_1_or_1_cse
        & (mux_33_nl) ) begin
      FpSignedBitsToFloat_6U_10U_1_slc_FpSignedBitsToFloat_6U_10U_1_ubits_9_0_itm_3
          <= MUX_v_10_2_2((FpSignedBitsToFloat_6U_10U_bits_1_sva_1_15_0_1[9:0]),
          (FpSignedBitsToFloat_6U_10U_bits_sva_1_15_0_1[9:0]), and_dcpl_38);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpSignedBitsToFloat_6U_10U_1_slc_FpSignedBitsToFloat_6U_10U_1_ubits_15_10_itm_3
          <= 6'b0;
    end
    else if ( core_wen & FpSignedBitsToFloat_6U_10U_1_FpSignedBitsToFloat_6U_10U_1_or_1_cse
        & (mux_35_nl) ) begin
      FpSignedBitsToFloat_6U_10U_1_slc_FpSignedBitsToFloat_6U_10U_1_ubits_15_10_itm_3
          <= MUX_v_6_2_2((FpSignedBitsToFloat_6U_10U_bits_1_sva_1_15_0_1[15:10]),
          (FpSignedBitsToFloat_6U_10U_bits_sva_1_15_0_1[15:10]), and_dcpl_38);
    end
  end
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn) begin
    if ( ~ nvdla_core_rstn ) begin
      FpAdd_6U_10U_mux_13_itm_4 <= 1'b0;
    end
    else if ( core_wen & ((or_5_cse & IsNaN_6U_10U_IsNaN_6U_10U_nor_tmp) | (or_61_cse
        & and_58_m1c) | FpSignedBitsToFloat_6U_10U_or_1_rgt) & mux_24_cse ) begin
      FpAdd_6U_10U_mux_13_itm_4 <= MUX_s_1_2_2((chn_a_rsci_d_mxwt[16]), (chn_b_rsci_d_mxwt[16]),
          FpSignedBitsToFloat_6U_10U_or_1_rgt);
    end
  end
  assign nl_FpMantRNE_23U_11U_else_acc_nl = FpSignedBitsToFloat_6U_10U_1_slc_FpSignedBitsToFloat_6U_10U_1_ubits_9_0_itm_4
      + conv_u2u_1_10(FpMantRNE_23U_11U_else_carry_sva_2);
  assign FpMantRNE_23U_11U_else_acc_nl = nl_FpMantRNE_23U_11U_else_acc_nl[9:0];
  assign FpAdd_6U_10U_FpAdd_6U_10U_or_2_nl = MUX_v_10_2_2((FpMantRNE_23U_11U_else_acc_nl),
      10'b1111111111, FpAdd_6U_10U_is_inf_lpi_1_dfm_2_mx0);
  assign FpSignedBitsToFloat_6U_10U_1_and_nl = (~ IsNaN_6U_10U_1_land_lpi_1_dfm_6)
      & chn_o_rsci_d_9_0_mx0c1;
  assign nl_FpAdd_6U_10U_if_4_if_acc_nl = FpAdd_6U_10U_o_expo_lpi_1_dfm_10 + 6'b1;
  assign FpAdd_6U_10U_if_4_if_acc_nl = nl_FpAdd_6U_10U_if_4_if_acc_nl[5:0];
  assign FpAdd_6U_10U_and_nl = (~(FpAdd_6U_10U_and_tmp | FpAdd_6U_10U_is_inf_lpi_1_dfm_2_mx0))
      & FpAdd_6U_10U_FpAdd_6U_10U_nor_2_m1c;
  assign FpAdd_6U_10U_and_3_nl = FpAdd_6U_10U_and_tmp & (~ FpAdd_6U_10U_is_inf_lpi_1_dfm_2_mx0)
      & FpAdd_6U_10U_FpAdd_6U_10U_nor_2_m1c;
  assign FpAdd_6U_10U_and_7_nl = FpAdd_6U_10U_is_inf_lpi_1_dfm_2_mx0 & FpAdd_6U_10U_FpAdd_6U_10U_nor_2_m1c;
  assign FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl = ~(MUX_v_6_2_2(6'b000000,
      z_out, or_61_cse));
  assign nl_FpAdd_6U_10U_b_left_shift_acc_itm_2  = ({1'b1 , (FpAdd_6U_10U_b_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl)})
      + 7'b1101;
  assign FpAdd_6U_10U_is_a_greater_oelse_not_5_nl = ~ or_61_cse;
  assign FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl = ~(MUX_v_6_2_2(6'b000000,
      z_out, (FpAdd_6U_10U_is_a_greater_oelse_not_5_nl)));
  assign nl_FpAdd_6U_10U_a_left_shift_acc_itm_2  = ({1'b1 , (FpAdd_6U_10U_a_left_shift_FpAdd_6U_10U_a_right_shift_nand_nl)})
      + 7'b1101;
  assign FpAdd_6U_10U_else_2_mux_2_nl = MUX_v_23_2_2((~ FpAdd_6U_10U_addend_smaller_qr_lpi_1_dfm_mx0),
      FpAdd_6U_10U_addend_larger_qr_lpi_1_dfm_mx0, FpAdd_6U_10U_if_2_and_tmp);
  assign FpAdd_6U_10U_else_2_mux_3_nl = MUX_v_23_2_2(FpAdd_6U_10U_addend_larger_qr_lpi_1_dfm_mx0,
      FpAdd_6U_10U_addend_smaller_qr_lpi_1_dfm_mx0, FpAdd_6U_10U_if_2_and_tmp);
  assign nl_acc_1_nl = ({(~ FpAdd_6U_10U_if_2_and_tmp) , (FpAdd_6U_10U_else_2_mux_2_nl)
      , (~ FpAdd_6U_10U_if_2_and_tmp)}) + conv_u2u_24_25({(FpAdd_6U_10U_else_2_mux_3_nl)
      , 1'b1});
  assign acc_1_nl = nl_acc_1_nl[24:0];
  assign nor_35_nl = ~(nor_3_cse | (~ main_stage_v_2) | IsNaN_6U_10U_land_lpi_1_dfm_st_5
      | IsNaN_6U_10U_1_land_lpi_1_dfm_5);
  assign nor_36_nl = ~((~ main_stage_v_3) | IsNaN_6U_10U_land_lpi_1_dfm_6 | IsNaN_6U_10U_1_land_lpi_1_dfm_6
      | FpAdd_6U_10U_is_inf_lpi_1_dfm_4);
  assign mux_3_nl = MUX_s_1_2_2((nor_36_nl), (nor_35_nl), or_5_cse);
  assign nl_FpNormalize_6U_23U_else_acc_nl = FpAdd_6U_10U_qr_lpi_1_dfm_4 + ({1'b1
      , (~ libraries_leading_sign_23_0_b9d2f049d7a95593b985a5e76dea79445444_1)})
      + 6'b1;
  assign FpNormalize_6U_23U_else_acc_nl = nl_FpNormalize_6U_23U_else_acc_nl[5:0];
  assign FpNormalize_6U_23U_FpNormalize_6U_23U_and_nl = MUX_v_6_2_2(6'b000000, (FpNormalize_6U_23U_else_acc_nl),
      FpNormalize_6U_23U_oelse_not_3);
  assign nl_FpAdd_6U_10U_if_3_if_acc_nl = FpAdd_6U_10U_qr_lpi_1_dfm_4 + 6'b1;
  assign FpAdd_6U_10U_if_3_if_acc_nl = nl_FpAdd_6U_10U_if_3_if_acc_nl[5:0];
  assign and_11_nl = main_stage_v_2 & mux_tmp_6;
  assign or_18_nl = IsNaN_6U_10U_land_lpi_1_dfm_6 | IsNaN_6U_10U_1_land_lpi_1_dfm_6
      | FpAdd_6U_10U_is_inf_lpi_1_dfm_4;
  assign mux_9_nl = MUX_s_1_2_2(mux_tmp_8, (and_11_nl), or_18_nl);
  assign mux_10_nl = MUX_s_1_2_2((mux_9_nl), mux_tmp_8, FpMantRNE_23U_11U_else_and_svs_2);
  assign mux_11_nl = MUX_s_1_2_2(or_tmp_25, (~ or_5_cse), nor_24_cse);
  assign mux_12_nl = MUX_s_1_2_2((mux_11_nl), or_tmp_25, IsNaN_6U_10U_land_lpi_1_dfm_st_5);
  assign nor_25_nl = ~(nor_24_cse | (~ and_41_cse));
  assign mux_13_nl = MUX_s_1_2_2((nor_25_nl), and_41_cse, IsNaN_6U_10U_land_lpi_1_dfm_st_5);
  assign and_84_nl = ((~ FpAdd_6U_10U_is_inf_lpi_1_dfm_4) | IsNaN_6U_10U_1_land_lpi_1_dfm_6
      | IsNaN_6U_10U_land_lpi_1_dfm_6) & main_stage_v_3;
  assign mux_14_nl = MUX_s_1_2_2((mux_13_nl), (mux_12_nl), and_84_nl);
  assign or_35_nl = nor_7_cse | nor_tmp_8;
  assign nor_22_nl = ~(reg_chn_o_rsci_ld_core_psct_cse | (~ nor_tmp_8));
  assign mux_17_nl = MUX_s_1_2_2((nor_22_nl), nor_tmp_8, chn_o_rsci_bawt);
  assign and_82_nl = FpAdd_6U_10U_or_cse & main_stage_v_3;
  assign mux_18_nl = MUX_s_1_2_2((mux_17_nl), (or_35_nl), and_82_nl);
  assign and_91_nl = (~ nor_tmp_8) & reg_chn_o_rsci_ld_core_psct_cse & (~ chn_o_rsci_bawt);
  assign mux_31_nl = MUX_s_1_2_2(or_tmp_43, (and_91_nl), IsNaN_6U_10U_1_land_lpi_1_dfm_4);
  assign mux_32_nl = MUX_s_1_2_2((~ (mux_31_nl)), or_75_cse, IsNaN_6U_10U_land_lpi_1_dfm_st_4);
  assign mux_33_nl = MUX_s_1_2_2((~ or_tmp_43), (mux_32_nl), main_stage_v_1);
  assign or_44_nl = IsNaN_6U_10U_land_lpi_1_dfm_st_4 | IsNaN_6U_10U_1_land_lpi_1_dfm_4;
  assign mux_34_nl = MUX_s_1_2_2(not_tmp_34, or_75_cse, or_44_nl);
  assign mux_35_nl = MUX_s_1_2_2(not_tmp_34, (mux_34_nl), main_stage_v_1);
  assign FpAdd_6U_10U_b_right_shift_qif_mux_2_nl = MUX_v_6_2_2((chn_a_rsci_d_mxwt[15:10]),
      (chn_b_rsci_d_mxwt[15:10]), FpAdd_6U_10U_a_right_shift_qelse_and_tmp);
  assign FpAdd_6U_10U_b_right_shift_qif_mux_3_nl = MUX_v_6_2_2((~ (chn_b_rsci_d_mxwt[15:10])),
      (~ (chn_a_rsci_d_mxwt[15:10])), FpAdd_6U_10U_a_right_shift_qelse_and_tmp);
  assign nl_acc_nl = ({(FpAdd_6U_10U_b_right_shift_qif_mux_2_nl) , 1'b1}) + ({(FpAdd_6U_10U_b_right_shift_qif_mux_3_nl)
      , 1'b1});
  assign acc_nl = nl_acc_nl[6:0];
  assign z_out = readslicef_7_6_1((acc_nl));

  function [5:0] MUX1HOT_v_6_3_2;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [2:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | ( input_1 & {6{sel[1]}});
    result = result | ( input_2 & {6{sel[2]}});
    MUX1HOT_v_6_3_2 = result;
  end
  endfunction


  function [5:0] MUX1HOT_v_6_4_2;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [3:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | ( input_1 & {6{sel[1]}});
    result = result | ( input_2 & {6{sel[2]}});
    result = result | ( input_3 & {6{sel[3]}});
    MUX1HOT_v_6_4_2 = result;
  end
  endfunction


  function [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function [21:0] MUX_v_22_2_2;
    input [21:0] input_0;
    input [21:0] input_1;
    input [0:0] sel;
    reg [21:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_22_2_2 = result;
  end
  endfunction


  function [22:0] MUX_v_23_2_2;
    input [22:0] input_0;
    input [22:0] input_1;
    input [0:0] sel;
    reg [22:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_23_2_2 = result;
  end
  endfunction


  function [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function [0:0] readslicef_11_1_10;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_11_1_10 = tmp[0:0];
  end
  endfunction


  function [23:0] readslicef_25_24_1;
    input [24:0] vector;
    reg [24:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_25_24_1 = tmp[23:0];
  end
  endfunction


  function [0:0] readslicef_6_1_5;
    input [5:0] vector;
    reg [5:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_6_1_5 = tmp[0:0];
  end
  endfunction


  function [0:0] readslicef_7_1_6;
    input [6:0] vector;
    reg [6:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_7_1_6 = tmp[0:0];
  end
  endfunction


  function [5:0] readslicef_7_6_1;
    input [6:0] vector;
    reg [6:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_7_6_1 = tmp[5:0];
  end
  endfunction


  function  [6:0] conv_u2s_5_7 ;
    input [4:0]  vector ;
  begin
    conv_u2s_5_7 = {{2{1'b0}}, vector};
  end
  endfunction


  function  [9:0] conv_u2u_1_10 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_10 = {{9{1'b0}}, vector};
  end
  endfunction


  function  [6:0] conv_u2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_7 = {1'b0, vector};
  end
  endfunction


  function  [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction


  function  [24:0] conv_u2u_24_25 ;
    input [23:0]  vector ;
  begin
    conv_u2u_24_25 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    HLS_fp17_add
// ------------------------------------------------------------------


module HLS_fp17_add (
  nvdla_core_clk, nvdla_core_rstn, chn_a_rsc_z, chn_a_rsc_vz, chn_a_rsc_lz, chn_b_rsc_z,
      chn_b_rsc_vz, chn_b_rsc_lz, chn_o_rsc_z, chn_o_rsc_vz, chn_o_rsc_lz
);
  input nvdla_core_clk;
  input nvdla_core_rstn;
  input [16:0] chn_a_rsc_z;
  input chn_a_rsc_vz;
  output chn_a_rsc_lz;
  input [16:0] chn_b_rsc_z;
  input chn_b_rsc_vz;
  output chn_b_rsc_lz;
  output [16:0] chn_o_rsc_z;
  input chn_o_rsc_vz;
  output chn_o_rsc_lz;


  // Interconnect Declarations
  wire chn_a_rsci_oswt;
  wire chn_b_rsci_oswt;
  wire chn_o_rsci_oswt;
  wire chn_o_rsci_oswt_unreg;
  wire chn_a_rsci_oswt_unreg_iff;


  // Interconnect Declarations for Component Instantiations 
  FP17_ADD_chn_a_rsci_unreg chn_a_rsci_unreg_inst (
      .in_0(chn_a_rsci_oswt_unreg_iff),
      .outsig(chn_a_rsci_oswt)
    );
  FP17_ADD_chn_b_rsci_unreg chn_b_rsci_unreg_inst (
      .in_0(chn_a_rsci_oswt_unreg_iff),
      .outsig(chn_b_rsci_oswt)
    );
  FP17_ADD_chn_o_rsci_unreg chn_o_rsci_unreg_inst (
      .in_0(chn_o_rsci_oswt_unreg),
      .outsig(chn_o_rsci_oswt)
    );
  HLS_fp17_add_core HLS_fp17_add_core_inst (
      .nvdla_core_clk(nvdla_core_clk),
      .nvdla_core_rstn(nvdla_core_rstn),
      .chn_a_rsc_z(chn_a_rsc_z),
      .chn_a_rsc_vz(chn_a_rsc_vz),
      .chn_a_rsc_lz(chn_a_rsc_lz),
      .chn_b_rsc_z(chn_b_rsc_z),
      .chn_b_rsc_vz(chn_b_rsc_vz),
      .chn_b_rsc_lz(chn_b_rsc_lz),
      .chn_o_rsc_z(chn_o_rsc_z),
      .chn_o_rsc_vz(chn_o_rsc_vz),
      .chn_o_rsc_lz(chn_o_rsc_lz),
      .chn_a_rsci_oswt(chn_a_rsci_oswt),
      .chn_b_rsci_oswt(chn_b_rsci_oswt),
      .chn_o_rsci_oswt(chn_o_rsci_oswt),
      .chn_o_rsci_oswt_unreg(chn_o_rsci_oswt_unreg),
      .chn_a_rsci_oswt_unreg_pff(chn_a_rsci_oswt_unreg_iff)
    );
endmodule



